`timescale 1 ps / 1 ps
`define XIL_TIMING

(* dont_touch = "true" *) 
(* NotValidForBitStream *)
module switch_elements
   (enable_i,
    clk_i,
    rst_i,
    info_o);
  input [31:0]enable_i;
  input clk_i;
  input rst_i;
  output [31:0]info_o;

  wire clk_i;
  wire [31:0]enable_i;
  wire [31:0]info_o;
  wire \info_o[28]_INST_0_i_2_n_0 ;
  wire \info_o[29]_INST_0_i_2_n_0 ;
  wire \info_o[29]_INST_0_i_3_n_0 ;
  wire \info_o[30]_INST_0_i_1_n_0 ;
  wire \info_o[31]_INST_0_i_1_n_0 ;
  wire \info_o[31]_INST_0_i_3_n_0 ;
  wire \info_o[3]_INST_0_i_1_n_0 ;
  wire \info_o[3]_INST_0_i_2_n_0 ;
  wire rst_i;
  wire switch_n_32;
  wire switch_n_33;

  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \info_o[28]_INST_0_i_2 
       (.I0(switch_n_33),
        .I1(switch_n_32),
        .I2(enable_i[4]),
        .I3(enable_i[5]),
        .I4(enable_i[1]),
        .I5(enable_i[0]),
        .O(\info_o[28]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000007)) 
    \info_o[29]_INST_0_i_2 
       (.I0(enable_i[3]),
        .I1(enable_i[2]),
        .I2(switch_n_32),
        .I3(enable_i[4]),
        .I4(enable_i[5]),
        .I5(\info_o[29]_INST_0_i_3_n_0 ),
        .O(\info_o[29]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \info_o[29]_INST_0_i_3 
       (.I0(enable_i[1]),
        .I1(enable_i[0]),
        .O(\info_o[29]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \info_o[30]_INST_0_i_1 
       (.I0(enable_i[5]),
        .I1(enable_i[4]),
        .I2(switch_n_32),
        .I3(enable_i[1]),
        .I4(enable_i[0]),
        .I5(enable_i[2]),
        .O(\info_o[30]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \info_o[31]_INST_0_i_1 
       (.I0(\info_o[31]_INST_0_i_3_n_0 ),
        .I1(enable_i[0]),
        .I2(enable_i[1]),
        .O(\info_o[31]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFFFFFFFF)) 
    \info_o[31]_INST_0_i_3 
       (.I0(enable_i[8]),
        .I1(enable_i[9]),
        .I2(enable_i[7]),
        .I3(enable_i[5]),
        .I4(enable_i[4]),
        .I5(enable_i[6]),
        .O(\info_o[31]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFEF)) 
    \info_o[3]_INST_0_i_1 
       (.I0(switch_n_32),
        .I1(enable_i[3]),
        .I2(enable_i[5]),
        .I3(enable_i[4]),
        .I4(enable_i[2]),
        .O(\info_o[3]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \info_o[3]_INST_0_i_2 
       (.I0(\info_o[31]_INST_0_i_3_n_0 ),
        .I1(enable_i[0]),
        .I2(enable_i[1]),
        .O(\info_o[3]_INST_0_i_2_n_0 ));
  switch_elements_aes switch
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .enable_i_3_sp_1(switch_n_33),
        .enable_i_6_sp_1(switch_n_32),
        .info_o(info_o),
        .\info_o[0]_0 (\info_o[31]_INST_0_i_1_n_0 ),
        .info_o_0_sp_1(\info_o[3]_INST_0_i_2_n_0 ),
        .info_o_2_sp_1(\info_o[3]_INST_0_i_1_n_0 ),
        .info_o_4_sp_1(\info_o[28]_INST_0_i_2_n_0 ),
        .info_o_5_sp_1(\info_o[29]_INST_0_i_2_n_0 ),
        .info_o_9_sp_1(\info_o[30]_INST_0_i_1_n_0 ),
        .rst_i(rst_i));
endmodule

(* ORIG_REF_NAME = "aes" *) 
module switch_elements_aes
   (info_o,
    enable_i_6_sp_1,
    enable_i_3_sp_1,
    clk_i,
    rst_i,
    enable_i,
    info_o_0_sp_1,
    \info_o[0]_0 ,
    info_o_2_sp_1,
    info_o_4_sp_1,
    info_o_5_sp_1,
    info_o_9_sp_1);
  output [31:0]info_o;
  output enable_i_6_sp_1;
  output enable_i_3_sp_1;
  input clk_i;
  input rst_i;
  input [31:0]enable_i;
  input info_o_0_sp_1;
  input \info_o[0]_0 ;
  input info_o_2_sp_1;
  input info_o_4_sp_1;
  input info_o_5_sp_1;
  input info_o_9_sp_1;

  wire block_reg;
  wire \block_reg[1][31]_i_1_n_0 ;
  wire \block_reg[2][31]_i_1_n_0 ;
  wire \block_reg[3][31]_i_1_n_0 ;
  wire \block_reg[3][31]_i_2_n_0 ;
  wire clk_i;
  wire config_we4_out;
  wire [127:0]core_block;
  wire [255:0]core_key;
  wire core_ready;
  wire [127:0]core_result;
  wire core_valid;
  wire [31:0]enable_i;
  wire enable_i_3_sn_1;
  wire enable_i_6_sn_1;
  wire [31:0]info_o;
  wire \info_o[0]_0 ;
  wire \info_o[0]_INST_0_i_1_n_0 ;
  wire \info_o[0]_INST_0_i_2_n_0 ;
  wire \info_o[10]_INST_0_i_1_n_0 ;
  wire \info_o[11]_INST_0_i_1_n_0 ;
  wire \info_o[12]_INST_0_i_1_n_0 ;
  wire \info_o[13]_INST_0_i_1_n_0 ;
  wire \info_o[14]_INST_0_i_1_n_0 ;
  wire \info_o[15]_INST_0_i_1_n_0 ;
  wire \info_o[16]_INST_0_i_1_n_0 ;
  wire \info_o[17]_INST_0_i_1_n_0 ;
  wire \info_o[18]_INST_0_i_1_n_0 ;
  wire \info_o[19]_INST_0_i_1_n_0 ;
  wire \info_o[1]_INST_0_i_2_n_0 ;
  wire \info_o[1]_INST_0_i_3_n_0 ;
  wire \info_o[20]_INST_0_i_1_n_0 ;
  wire \info_o[21]_INST_0_i_1_n_0 ;
  wire \info_o[22]_INST_0_i_1_n_0 ;
  wire \info_o[23]_INST_0_i_1_n_0 ;
  wire \info_o[24]_INST_0_i_1_n_0 ;
  wire \info_o[25]_INST_0_i_1_n_0 ;
  wire \info_o[26]_INST_0_i_1_n_0 ;
  wire \info_o[27]_INST_0_i_1_n_0 ;
  wire \info_o[28]_INST_0_i_1_n_0 ;
  wire \info_o[29]_INST_0_i_1_n_0 ;
  wire \info_o[2]_INST_0_i_1_n_0 ;
  wire \info_o[30]_INST_0_i_2_n_0 ;
  wire \info_o[31]_INST_0_i_2_n_0 ;
  wire \info_o[3]_INST_0_i_3_n_0 ;
  wire \info_o[4]_INST_0_i_1_n_0 ;
  wire \info_o[5]_INST_0_i_1_n_0 ;
  wire \info_o[6]_INST_0_i_1_n_0 ;
  wire \info_o[7]_INST_0_i_1_n_0 ;
  wire \info_o[8]_INST_0_i_1_n_0 ;
  wire \info_o[9]_INST_0_i_1_n_0 ;
  wire info_o_0_sn_1;
  wire info_o_2_sn_1;
  wire info_o_4_sn_1;
  wire info_o_5_sn_1;
  wire info_o_9_sn_1;
  wire init_new0_out;
  wire init_reg_i_2_n_0;
  wire init_reg_i_3_n_0;
  wire key_reg;
  wire \key_reg[1][31]_i_1_n_0 ;
  wire \key_reg[2][31]_i_1_n_0 ;
  wire \key_reg[3][31]_i_1_n_0 ;
  wire \key_reg[3][31]_i_2_n_0 ;
  wire \key_reg[4][31]_i_1_n_0 ;
  wire \key_reg[5][31]_i_1_n_0 ;
  wire \key_reg[6][31]_i_1_n_0 ;
  wire \key_reg[7][31]_i_1_n_0 ;
  wire \key_reg[7][31]_i_2_n_0 ;
  wire keylen_reg_reg_rep__0_n_0;
  wire keylen_reg_reg_rep_n_0;
  wire next_new1_out;
  wire [3:0]p_1_in;
  wire ready_reg;
  wire [127:0]result_reg;
  wire rst_i;
  wire valid_reg;

  assign enable_i_3_sp_1 = enable_i_3_sn_1;
  assign enable_i_6_sp_1 = enable_i_6_sn_1;
  assign info_o_0_sn_1 = info_o_0_sp_1;
  assign info_o_2_sn_1 = info_o_2_sp_1;
  assign info_o_4_sn_1 = info_o_4_sp_1;
  assign info_o_5_sn_1 = info_o_5_sp_1;
  assign info_o_9_sn_1 = info_o_9_sp_1;
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \block_reg[0][31]_i_1 
       (.I0(enable_i[1]),
        .I1(enable_i[0]),
        .I2(enable_i[6]),
        .I3(\block_reg[3][31]_i_2_n_0 ),
        .I4(enable_i[3]),
        .I5(enable_i[2]),
        .O(block_reg));
  LUT6 #(
    .INIT(64'h0000000000080000)) 
    \block_reg[1][31]_i_1 
       (.I0(enable_i[1]),
        .I1(enable_i[0]),
        .I2(enable_i[6]),
        .I3(\block_reg[3][31]_i_2_n_0 ),
        .I4(enable_i[2]),
        .I5(enable_i[3]),
        .O(\block_reg[1][31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \block_reg[2][31]_i_1 
       (.I0(enable_i[1]),
        .I1(enable_i[0]),
        .I2(enable_i[6]),
        .I3(\block_reg[3][31]_i_2_n_0 ),
        .I4(enable_i[2]),
        .I5(enable_i[3]),
        .O(\block_reg[2][31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \block_reg[3][31]_i_1 
       (.I0(enable_i[1]),
        .I1(enable_i[0]),
        .I2(enable_i[6]),
        .I3(\block_reg[3][31]_i_2_n_0 ),
        .I4(enable_i[3]),
        .I5(enable_i[2]),
        .O(\block_reg[3][31]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT5 #(
    .INIT(32'hFFFFFFEF)) 
    \block_reg[3][31]_i_2 
       (.I0(enable_i[4]),
        .I1(enable_i[5]),
        .I2(enable_i[7]),
        .I3(enable_i[9]),
        .I4(enable_i[8]),
        .O(\block_reg[3][31]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][0] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(core_block[96]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][10] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(core_block[106]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][11] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(core_block[107]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][12] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(core_block[108]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][13] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(core_block[109]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][14] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(core_block[110]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][15] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(core_block[111]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][16] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(core_block[112]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][17] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(core_block[113]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][18] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(core_block[114]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][19] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(core_block[115]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][1] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(core_block[97]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][20] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(core_block[116]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][21] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(core_block[117]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][22] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(core_block[118]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][23] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(core_block[119]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][24] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(core_block[120]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][25] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(core_block[121]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][26] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(core_block[122]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][27] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(core_block[123]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][28] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(core_block[124]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][29] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(core_block[125]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][2] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(core_block[98]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][30] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(core_block[126]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][31] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(core_block[127]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][3] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(core_block[99]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][4] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(core_block[100]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][5] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(core_block[101]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][6] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(core_block[102]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][7] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(core_block[103]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][8] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(core_block[104]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[0][9] 
       (.C(clk_i),
        .CE(block_reg),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(core_block[105]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][0] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(core_block[64]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][10] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(core_block[74]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][11] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(core_block[75]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][12] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(core_block[76]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][13] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(core_block[77]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][14] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(core_block[78]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][15] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(core_block[79]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][16] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(core_block[80]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][17] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(core_block[81]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][18] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(core_block[82]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][19] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(core_block[83]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][1] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(core_block[65]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][20] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(core_block[84]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][21] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(core_block[85]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][22] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(core_block[86]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][23] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(core_block[87]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][24] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(core_block[88]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][25] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(core_block[89]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][26] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(core_block[90]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][27] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(core_block[91]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][28] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(core_block[92]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][29] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(core_block[93]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][2] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(core_block[66]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][30] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(core_block[94]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][31] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(core_block[95]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][3] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(core_block[67]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][4] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(core_block[68]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][5] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(core_block[69]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][6] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(core_block[70]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][7] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(core_block[71]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][8] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(core_block[72]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[1][9] 
       (.C(clk_i),
        .CE(\block_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(core_block[73]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][0] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(core_block[32]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][10] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(core_block[42]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][11] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(core_block[43]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][12] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(core_block[44]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][13] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(core_block[45]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][14] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(core_block[46]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][15] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(core_block[47]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][16] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(core_block[48]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][17] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(core_block[49]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][18] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(core_block[50]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][19] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(core_block[51]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][1] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(core_block[33]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][20] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(core_block[52]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][21] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(core_block[53]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][22] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(core_block[54]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][23] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(core_block[55]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][24] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(core_block[56]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][25] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(core_block[57]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][26] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(core_block[58]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][27] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(core_block[59]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][28] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(core_block[60]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][29] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(core_block[61]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][2] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(core_block[34]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][30] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(core_block[62]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][31] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(core_block[63]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][3] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(core_block[35]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][4] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(core_block[36]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][5] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(core_block[37]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][6] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(core_block[38]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][7] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(core_block[39]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][8] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(core_block[40]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[2][9] 
       (.C(clk_i),
        .CE(\block_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(core_block[41]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][0] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(core_block[0]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][10] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(core_block[10]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][11] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(core_block[11]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][12] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(core_block[12]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][13] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(core_block[13]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][14] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(core_block[14]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][15] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(core_block[15]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][16] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(core_block[16]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][17] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(core_block[17]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][18] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(core_block[18]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][19] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(core_block[19]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][1] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(core_block[1]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][20] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(core_block[20]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][21] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(core_block[21]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][22] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(core_block[22]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][23] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(core_block[23]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][24] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(core_block[24]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][25] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(core_block[25]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][26] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(core_block[26]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][27] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(core_block[27]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][28] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(core_block[28]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][29] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(core_block[29]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][2] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(core_block[2]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][30] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(core_block[30]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][31] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(core_block[31]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][3] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(core_block[3]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][4] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(core_block[4]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][5] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(core_block[5]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][6] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(core_block[6]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][7] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(core_block[7]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][8] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(core_block[8]));
  FDCE #(
    .INIT(1'b0)) 
    \block_reg_reg[3][9] 
       (.C(clk_i),
        .CE(\block_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(core_block[9]));
  switch_elements_aes_core core
       (.D(core_result),
        .clk_i(clk_i),
        .core_block(core_block),
        .core_key(core_key),
        .core_valid(core_valid),
        .\key_mem_reg[14][127] (keylen_reg_reg_rep__0_n_0),
        .\key_mem_reg[14][36] (keylen_reg_reg_rep_n_0),
        .p_1_in(p_1_in),
        .ready(core_ready),
        .rst_i(rst_i));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    encdec_reg_i_1
       (.I0(enable_i_6_sn_1),
        .I1(enable_i[5]),
        .I2(enable_i[0]),
        .I3(enable_i_3_sn_1),
        .I4(enable_i[4]),
        .I5(enable_i[1]),
        .O(config_we4_out));
  FDCE #(
    .INIT(1'b0)) 
    encdec_reg_reg
       (.C(clk_i),
        .CE(config_we4_out),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(p_1_in[2]));
  LUT5 #(
    .INIT(32'hFF101010)) 
    \info_o[0]_INST_0 
       (.I0(enable_i_6_sn_1),
        .I1(\info_o[0]_INST_0_i_1_n_0 ),
        .I2(info_o_0_sn_1),
        .I3(\info_o[0]_0 ),
        .I4(\info_o[0]_INST_0_i_2_n_0 ),
        .O(info_o[0]));
  LUT6 #(
    .INIT(64'hFBFBFBFFFFFFFBFF)) 
    \info_o[0]_INST_0_i_1 
       (.I0(enable_i[4]),
        .I1(enable_i[5]),
        .I2(enable_i[3]),
        .I3(p_1_in[0]),
        .I4(enable_i[2]),
        .I5(ready_reg),
        .O(\info_o[0]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[0]_INST_0_i_2 
       (.I0(result_reg[0]),
        .I1(result_reg[64]),
        .I2(enable_i[2]),
        .I3(result_reg[32]),
        .I4(enable_i[3]),
        .I5(result_reg[96]),
        .O(\info_o[0]_INST_0_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \info_o[10]_INST_0 
       (.I0(info_o_4_sn_1),
        .I1(\info_o[0]_0 ),
        .I2(\info_o[10]_INST_0_i_1_n_0 ),
        .O(info_o[10]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[10]_INST_0_i_1 
       (.I0(result_reg[10]),
        .I1(result_reg[74]),
        .I2(enable_i[2]),
        .I3(result_reg[42]),
        .I4(enable_i[3]),
        .I5(result_reg[106]),
        .O(\info_o[10]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \info_o[11]_INST_0 
       (.I0(\info_o[0]_0 ),
        .I1(\info_o[11]_INST_0_i_1_n_0 ),
        .O(info_o[11]));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \info_o[11]_INST_0_i_1 
       (.I0(result_reg[43]),
        .I1(result_reg[107]),
        .I2(enable_i[2]),
        .I3(result_reg[11]),
        .I4(enable_i[3]),
        .I5(result_reg[75]),
        .O(\info_o[11]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \info_o[12]_INST_0 
       (.I0(info_o_9_sn_1),
        .I1(\info_o[0]_0 ),
        .I2(\info_o[12]_INST_0_i_1_n_0 ),
        .O(info_o[12]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[12]_INST_0_i_1 
       (.I0(result_reg[12]),
        .I1(result_reg[76]),
        .I2(enable_i[2]),
        .I3(result_reg[44]),
        .I4(enable_i[3]),
        .I5(result_reg[108]),
        .O(\info_o[12]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \info_o[13]_INST_0 
       (.I0(info_o_5_sn_1),
        .I1(\info_o[0]_0 ),
        .I2(\info_o[13]_INST_0_i_1_n_0 ),
        .O(info_o[13]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[13]_INST_0_i_1 
       (.I0(result_reg[13]),
        .I1(result_reg[77]),
        .I2(enable_i[2]),
        .I3(result_reg[45]),
        .I4(enable_i[3]),
        .I5(result_reg[109]),
        .O(\info_o[13]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT4 #(
    .INIT(16'hF222)) 
    \info_o[14]_INST_0 
       (.I0(info_o_9_sn_1),
        .I1(enable_i[3]),
        .I2(\info_o[0]_0 ),
        .I3(\info_o[14]_INST_0_i_1_n_0 ),
        .O(info_o[14]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[14]_INST_0_i_1 
       (.I0(result_reg[14]),
        .I1(result_reg[78]),
        .I2(enable_i[2]),
        .I3(result_reg[46]),
        .I4(enable_i[3]),
        .I5(result_reg[110]),
        .O(\info_o[14]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \info_o[15]_INST_0 
       (.I0(\info_o[0]_0 ),
        .I1(\info_o[15]_INST_0_i_1_n_0 ),
        .O(info_o[15]));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \info_o[15]_INST_0_i_1 
       (.I0(result_reg[47]),
        .I1(result_reg[111]),
        .I2(enable_i[2]),
        .I3(result_reg[15]),
        .I4(enable_i[3]),
        .I5(result_reg[79]),
        .O(\info_o[15]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT4 #(
    .INIT(16'hF222)) 
    \info_o[16]_INST_0 
       (.I0(info_o_9_sn_1),
        .I1(enable_i[3]),
        .I2(\info_o[0]_0 ),
        .I3(\info_o[16]_INST_0_i_1_n_0 ),
        .O(info_o[16]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[16]_INST_0_i_1 
       (.I0(result_reg[16]),
        .I1(result_reg[80]),
        .I2(enable_i[2]),
        .I3(result_reg[48]),
        .I4(enable_i[3]),
        .I5(result_reg[112]),
        .O(\info_o[16]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \info_o[17]_INST_0 
       (.I0(info_o_4_sn_1),
        .I1(\info_o[0]_0 ),
        .I2(\info_o[17]_INST_0_i_1_n_0 ),
        .O(info_o[17]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[17]_INST_0_i_1 
       (.I0(result_reg[17]),
        .I1(result_reg[81]),
        .I2(enable_i[2]),
        .I3(result_reg[49]),
        .I4(enable_i[3]),
        .I5(result_reg[113]),
        .O(\info_o[17]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \info_o[18]_INST_0 
       (.I0(info_o_9_sn_1),
        .I1(\info_o[0]_0 ),
        .I2(\info_o[18]_INST_0_i_1_n_0 ),
        .O(info_o[18]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[18]_INST_0_i_1 
       (.I0(result_reg[18]),
        .I1(result_reg[82]),
        .I2(enable_i[2]),
        .I3(result_reg[50]),
        .I4(enable_i[3]),
        .I5(result_reg[114]),
        .O(\info_o[18]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \info_o[19]_INST_0 
       (.I0(info_o_4_sn_1),
        .I1(\info_o[0]_0 ),
        .I2(\info_o[19]_INST_0_i_1_n_0 ),
        .O(info_o[19]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[19]_INST_0_i_1 
       (.I0(result_reg[19]),
        .I1(result_reg[83]),
        .I2(enable_i[2]),
        .I3(result_reg[51]),
        .I4(enable_i[3]),
        .I5(result_reg[115]),
        .O(\info_o[19]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFF101010)) 
    \info_o[1]_INST_0 
       (.I0(enable_i_6_sn_1),
        .I1(\info_o[1]_INST_0_i_2_n_0 ),
        .I2(info_o_0_sn_1),
        .I3(\info_o[0]_0 ),
        .I4(\info_o[1]_INST_0_i_3_n_0 ),
        .O(info_o[1]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \info_o[1]_INST_0_i_1 
       (.I0(enable_i[6]),
        .I1(enable_i[9]),
        .I2(enable_i[8]),
        .I3(enable_i[7]),
        .O(enable_i_6_sn_1));
  LUT6 #(
    .INIT(64'hFBFBFBFFFFFFFBFF)) 
    \info_o[1]_INST_0_i_2 
       (.I0(enable_i[4]),
        .I1(enable_i[5]),
        .I2(enable_i[3]),
        .I3(p_1_in[1]),
        .I4(enable_i[2]),
        .I5(valid_reg),
        .O(\info_o[1]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[1]_INST_0_i_3 
       (.I0(result_reg[1]),
        .I1(result_reg[65]),
        .I2(enable_i[2]),
        .I3(result_reg[33]),
        .I4(enable_i[3]),
        .I5(result_reg[97]),
        .O(\info_o[1]_INST_0_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \info_o[20]_INST_0 
       (.I0(\info_o[20]_INST_0_i_1_n_0 ),
        .I1(\info_o[0]_0 ),
        .O(info_o[20]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[20]_INST_0_i_1 
       (.I0(result_reg[20]),
        .I1(result_reg[84]),
        .I2(enable_i[2]),
        .I3(result_reg[52]),
        .I4(enable_i[3]),
        .I5(result_reg[116]),
        .O(\info_o[20]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \info_o[21]_INST_0 
       (.I0(info_o_5_sn_1),
        .I1(\info_o[0]_0 ),
        .I2(\info_o[21]_INST_0_i_1_n_0 ),
        .O(info_o[21]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[21]_INST_0_i_1 
       (.I0(result_reg[21]),
        .I1(result_reg[85]),
        .I2(enable_i[2]),
        .I3(result_reg[53]),
        .I4(enable_i[3]),
        .I5(result_reg[117]),
        .O(\info_o[21]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT4 #(
    .INIT(16'hF222)) 
    \info_o[22]_INST_0 
       (.I0(info_o_9_sn_1),
        .I1(enable_i[3]),
        .I2(\info_o[0]_0 ),
        .I3(\info_o[22]_INST_0_i_1_n_0 ),
        .O(info_o[22]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[22]_INST_0_i_1 
       (.I0(result_reg[22]),
        .I1(result_reg[86]),
        .I2(enable_i[2]),
        .I3(result_reg[54]),
        .I4(enable_i[3]),
        .I5(result_reg[118]),
        .O(\info_o[22]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \info_o[23]_INST_0 
       (.I0(\info_o[23]_INST_0_i_1_n_0 ),
        .I1(\info_o[0]_0 ),
        .O(info_o[23]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[23]_INST_0_i_1 
       (.I0(result_reg[23]),
        .I1(result_reg[87]),
        .I2(enable_i[2]),
        .I3(result_reg[55]),
        .I4(enable_i[3]),
        .I5(result_reg[119]),
        .O(\info_o[23]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT4 #(
    .INIT(16'hF222)) 
    \info_o[24]_INST_0 
       (.I0(info_o_9_sn_1),
        .I1(enable_i[3]),
        .I2(\info_o[0]_0 ),
        .I3(\info_o[24]_INST_0_i_1_n_0 ),
        .O(info_o[24]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[24]_INST_0_i_1 
       (.I0(result_reg[24]),
        .I1(result_reg[88]),
        .I2(enable_i[2]),
        .I3(result_reg[56]),
        .I4(enable_i[3]),
        .I5(result_reg[120]),
        .O(\info_o[24]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \info_o[25]_INST_0 
       (.I0(\info_o[0]_0 ),
        .I1(\info_o[25]_INST_0_i_1_n_0 ),
        .O(info_o[25]));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \info_o[25]_INST_0_i_1 
       (.I0(result_reg[57]),
        .I1(result_reg[121]),
        .I2(enable_i[2]),
        .I3(result_reg[25]),
        .I4(enable_i[3]),
        .I5(result_reg[89]),
        .O(\info_o[25]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \info_o[26]_INST_0 
       (.I0(\info_o[0]_0 ),
        .I1(\info_o[26]_INST_0_i_1_n_0 ),
        .O(info_o[26]));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \info_o[26]_INST_0_i_1 
       (.I0(result_reg[58]),
        .I1(result_reg[122]),
        .I2(enable_i[2]),
        .I3(result_reg[26]),
        .I4(enable_i[3]),
        .I5(result_reg[90]),
        .O(\info_o[26]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \info_o[27]_INST_0 
       (.I0(\info_o[0]_0 ),
        .I1(\info_o[27]_INST_0_i_1_n_0 ),
        .O(info_o[27]));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \info_o[27]_INST_0_i_1 
       (.I0(result_reg[59]),
        .I1(result_reg[123]),
        .I2(enable_i[2]),
        .I3(result_reg[27]),
        .I4(enable_i[3]),
        .I5(result_reg[91]),
        .O(\info_o[27]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    \info_o[28]_INST_0 
       (.I0(\info_o[0]_0 ),
        .I1(\info_o[28]_INST_0_i_1_n_0 ),
        .I2(info_o_4_sn_1),
        .O(info_o[28]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[28]_INST_0_i_1 
       (.I0(result_reg[28]),
        .I1(result_reg[92]),
        .I2(enable_i[2]),
        .I3(result_reg[60]),
        .I4(enable_i[3]),
        .I5(result_reg[124]),
        .O(\info_o[28]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \info_o[28]_INST_0_i_3 
       (.I0(enable_i[3]),
        .I1(enable_i[2]),
        .O(enable_i_3_sn_1));
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    \info_o[29]_INST_0 
       (.I0(\info_o[0]_0 ),
        .I1(\info_o[29]_INST_0_i_1_n_0 ),
        .I2(info_o_5_sn_1),
        .O(info_o[29]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[29]_INST_0_i_1 
       (.I0(result_reg[29]),
        .I1(result_reg[93]),
        .I2(enable_i[2]),
        .I3(result_reg[61]),
        .I4(enable_i[3]),
        .I5(result_reg[125]),
        .O(\info_o[29]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \info_o[2]_INST_0 
       (.I0(info_o_2_sn_1),
        .I1(p_1_in[2]),
        .I2(info_o_0_sn_1),
        .I3(\info_o[0]_0 ),
        .I4(\info_o[2]_INST_0_i_1_n_0 ),
        .O(info_o[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[2]_INST_0_i_1 
       (.I0(result_reg[2]),
        .I1(result_reg[66]),
        .I2(enable_i[2]),
        .I3(result_reg[34]),
        .I4(enable_i[3]),
        .I5(result_reg[98]),
        .O(\info_o[2]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT4 #(
    .INIT(16'hF222)) 
    \info_o[30]_INST_0 
       (.I0(info_o_9_sn_1),
        .I1(enable_i[3]),
        .I2(\info_o[0]_0 ),
        .I3(\info_o[30]_INST_0_i_2_n_0 ),
        .O(info_o[30]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[30]_INST_0_i_2 
       (.I0(result_reg[30]),
        .I1(result_reg[94]),
        .I2(enable_i[2]),
        .I3(result_reg[62]),
        .I4(enable_i[3]),
        .I5(result_reg[126]),
        .O(\info_o[30]_INST_0_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \info_o[31]_INST_0 
       (.I0(\info_o[0]_0 ),
        .I1(\info_o[31]_INST_0_i_2_n_0 ),
        .O(info_o[31]));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \info_o[31]_INST_0_i_2 
       (.I0(result_reg[63]),
        .I1(result_reg[127]),
        .I2(enable_i[2]),
        .I3(result_reg[31]),
        .I4(enable_i[3]),
        .I5(result_reg[95]),
        .O(\info_o[31]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \info_o[3]_INST_0 
       (.I0(info_o_2_sn_1),
        .I1(p_1_in[3]),
        .I2(info_o_0_sn_1),
        .I3(\info_o[0]_0 ),
        .I4(\info_o[3]_INST_0_i_3_n_0 ),
        .O(info_o[3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[3]_INST_0_i_3 
       (.I0(result_reg[3]),
        .I1(result_reg[67]),
        .I2(enable_i[2]),
        .I3(result_reg[35]),
        .I4(enable_i[3]),
        .I5(result_reg[99]),
        .O(\info_o[3]_INST_0_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \info_o[4]_INST_0 
       (.I0(info_o_4_sn_1),
        .I1(\info_o[0]_0 ),
        .I2(\info_o[4]_INST_0_i_1_n_0 ),
        .O(info_o[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[4]_INST_0_i_1 
       (.I0(result_reg[4]),
        .I1(result_reg[68]),
        .I2(enable_i[2]),
        .I3(result_reg[36]),
        .I4(enable_i[3]),
        .I5(result_reg[100]),
        .O(\info_o[4]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \info_o[5]_INST_0 
       (.I0(info_o_5_sn_1),
        .I1(\info_o[0]_0 ),
        .I2(\info_o[5]_INST_0_i_1_n_0 ),
        .O(info_o[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[5]_INST_0_i_1 
       (.I0(result_reg[5]),
        .I1(result_reg[69]),
        .I2(enable_i[2]),
        .I3(result_reg[37]),
        .I4(enable_i[3]),
        .I5(result_reg[101]),
        .O(\info_o[5]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \info_o[6]_INST_0 
       (.I0(\info_o[6]_INST_0_i_1_n_0 ),
        .I1(\info_o[0]_0 ),
        .O(info_o[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[6]_INST_0_i_1 
       (.I0(result_reg[6]),
        .I1(result_reg[70]),
        .I2(enable_i[2]),
        .I3(result_reg[38]),
        .I4(enable_i[3]),
        .I5(result_reg[102]),
        .O(\info_o[6]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \info_o[7]_INST_0 
       (.I0(\info_o[7]_INST_0_i_1_n_0 ),
        .I1(\info_o[0]_0 ),
        .O(info_o[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[7]_INST_0_i_1 
       (.I0(result_reg[7]),
        .I1(result_reg[71]),
        .I2(enable_i[2]),
        .I3(result_reg[39]),
        .I4(enable_i[3]),
        .I5(result_reg[103]),
        .O(\info_o[7]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT4 #(
    .INIT(16'hF222)) 
    \info_o[8]_INST_0 
       (.I0(info_o_9_sn_1),
        .I1(enable_i[3]),
        .I2(\info_o[0]_0 ),
        .I3(\info_o[8]_INST_0_i_1_n_0 ),
        .O(info_o[8]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[8]_INST_0_i_1 
       (.I0(result_reg[8]),
        .I1(result_reg[72]),
        .I2(enable_i[2]),
        .I3(result_reg[40]),
        .I4(enable_i[3]),
        .I5(result_reg[104]),
        .O(\info_o[8]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \info_o[9]_INST_0 
       (.I0(info_o_9_sn_1),
        .I1(\info_o[0]_0 ),
        .I2(\info_o[9]_INST_0_i_1_n_0 ),
        .O(info_o[9]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \info_o[9]_INST_0_i_1 
       (.I0(result_reg[9]),
        .I1(result_reg[73]),
        .I2(enable_i[2]),
        .I3(result_reg[41]),
        .I4(enable_i[3]),
        .I5(result_reg[105]),
        .O(\info_o[9]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    init_reg_i_1
       (.I0(enable_i[0]),
        .I1(enable_i[4]),
        .I2(init_reg_i_2_n_0),
        .I3(init_reg_i_3_n_0),
        .I4(enable_i[3]),
        .O(init_new0_out));
  LUT5 #(
    .INIT(32'h00000800)) 
    init_reg_i_2
       (.I0(enable_i[1]),
        .I1(enable_i[0]),
        .I2(enable_i[6]),
        .I3(enable_i[5]),
        .I4(enable_i[2]),
        .O(init_reg_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    init_reg_i_3
       (.I0(enable_i[7]),
        .I1(enable_i[8]),
        .I2(enable_i[9]),
        .O(init_reg_i_3_n_0));
  FDCE #(
    .INIT(1'b0)) 
    init_reg_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(init_new0_out),
        .Q(p_1_in[0]));
  LUT3 #(
    .INIT(8'h01)) 
    \key_reg[0][31]_i_1 
       (.I0(enable_i[3]),
        .I1(enable_i[2]),
        .I2(\key_reg[3][31]_i_2_n_0 ),
        .O(key_reg));
  LUT3 #(
    .INIT(8'h02)) 
    \key_reg[1][31]_i_1 
       (.I0(enable_i[2]),
        .I1(enable_i[3]),
        .I2(\key_reg[3][31]_i_2_n_0 ),
        .O(\key_reg[1][31]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \key_reg[2][31]_i_1 
       (.I0(enable_i[2]),
        .I1(enable_i[3]),
        .I2(\key_reg[3][31]_i_2_n_0 ),
        .O(\key_reg[2][31]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \key_reg[3][31]_i_1 
       (.I0(enable_i[3]),
        .I1(enable_i[2]),
        .I2(\key_reg[3][31]_i_2_n_0 ),
        .O(\key_reg[3][31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFBFFF)) 
    \key_reg[3][31]_i_2 
       (.I0(enable_i[4]),
        .I1(enable_i[0]),
        .I2(enable_i[1]),
        .I3(enable_i[6]),
        .I4(enable_i[5]),
        .I5(init_reg_i_3_n_0),
        .O(\key_reg[3][31]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \key_reg[4][31]_i_1 
       (.I0(\key_reg[7][31]_i_2_n_0 ),
        .I1(enable_i[3]),
        .I2(enable_i[2]),
        .O(\key_reg[4][31]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \key_reg[5][31]_i_1 
       (.I0(\key_reg[7][31]_i_2_n_0 ),
        .I1(enable_i[2]),
        .I2(enable_i[3]),
        .O(\key_reg[5][31]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \key_reg[6][31]_i_1 
       (.I0(enable_i[2]),
        .I1(enable_i[3]),
        .I2(\key_reg[7][31]_i_2_n_0 ),
        .O(\key_reg[6][31]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \key_reg[7][31]_i_1 
       (.I0(\key_reg[7][31]_i_2_n_0 ),
        .I1(enable_i[3]),
        .I2(enable_i[2]),
        .O(\key_reg[7][31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \key_reg[7][31]_i_2 
       (.I0(enable_i[4]),
        .I1(enable_i[0]),
        .I2(enable_i[1]),
        .I3(enable_i[6]),
        .I4(enable_i[5]),
        .I5(init_reg_i_3_n_0),
        .O(\key_reg[7][31]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][0] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(core_key[224]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][10] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(core_key[234]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][11] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(core_key[235]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][12] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(core_key[236]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][13] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(core_key[237]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][14] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(core_key[238]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][15] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(core_key[239]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][16] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(core_key[240]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][17] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(core_key[241]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][18] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(core_key[242]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][19] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(core_key[243]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][1] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(core_key[225]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][20] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(core_key[244]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][21] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(core_key[245]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][22] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(core_key[246]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][23] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(core_key[247]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][24] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(core_key[248]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][25] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(core_key[249]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][26] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(core_key[250]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][27] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(core_key[251]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][28] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(core_key[252]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][29] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(core_key[253]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][2] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(core_key[226]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][30] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(core_key[254]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][31] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(core_key[255]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][3] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(core_key[227]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][4] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(core_key[228]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][5] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(core_key[229]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][6] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(core_key[230]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][7] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(core_key[231]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][8] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(core_key[232]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[0][9] 
       (.C(clk_i),
        .CE(key_reg),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(core_key[233]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][0] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(core_key[192]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][10] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(core_key[202]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][11] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(core_key[203]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][12] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(core_key[204]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][13] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(core_key[205]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][14] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(core_key[206]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][15] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(core_key[207]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][16] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(core_key[208]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][17] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(core_key[209]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][18] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(core_key[210]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][19] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(core_key[211]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][1] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(core_key[193]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][20] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(core_key[212]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][21] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(core_key[213]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][22] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(core_key[214]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][23] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(core_key[215]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][24] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(core_key[216]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][25] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(core_key[217]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][26] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(core_key[218]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][27] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(core_key[219]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][28] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(core_key[220]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][29] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(core_key[221]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][2] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(core_key[194]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][30] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(core_key[222]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][31] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(core_key[223]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][3] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(core_key[195]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][4] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(core_key[196]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][5] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(core_key[197]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][6] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(core_key[198]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][7] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(core_key[199]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][8] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(core_key[200]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[1][9] 
       (.C(clk_i),
        .CE(\key_reg[1][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(core_key[201]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][0] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(core_key[160]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][10] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(core_key[170]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][11] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(core_key[171]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][12] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(core_key[172]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][13] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(core_key[173]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][14] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(core_key[174]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][15] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(core_key[175]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][16] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(core_key[176]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][17] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(core_key[177]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][18] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(core_key[178]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][19] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(core_key[179]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][1] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(core_key[161]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][20] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(core_key[180]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][21] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(core_key[181]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][22] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(core_key[182]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][23] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(core_key[183]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][24] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(core_key[184]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][25] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(core_key[185]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][26] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(core_key[186]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][27] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(core_key[187]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][28] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(core_key[188]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][29] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(core_key[189]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][2] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(core_key[162]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][30] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(core_key[190]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][31] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(core_key[191]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][3] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(core_key[163]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][4] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(core_key[164]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][5] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(core_key[165]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][6] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(core_key[166]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][7] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(core_key[167]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][8] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(core_key[168]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[2][9] 
       (.C(clk_i),
        .CE(\key_reg[2][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(core_key[169]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][0] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(core_key[128]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][10] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(core_key[138]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][11] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(core_key[139]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][12] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(core_key[140]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][13] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(core_key[141]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][14] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(core_key[142]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][15] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(core_key[143]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][16] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(core_key[144]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][17] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(core_key[145]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][18] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(core_key[146]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][19] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(core_key[147]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][1] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(core_key[129]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][20] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(core_key[148]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][21] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(core_key[149]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][22] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(core_key[150]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][23] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(core_key[151]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][24] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(core_key[152]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][25] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(core_key[153]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][26] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(core_key[154]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][27] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(core_key[155]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][28] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(core_key[156]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][29] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(core_key[157]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][2] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(core_key[130]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][30] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(core_key[158]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][31] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(core_key[159]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][3] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(core_key[131]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][4] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(core_key[132]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][5] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(core_key[133]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][6] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(core_key[134]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][7] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(core_key[135]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][8] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(core_key[136]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[3][9] 
       (.C(clk_i),
        .CE(\key_reg[3][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(core_key[137]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][0] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(core_key[96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][10] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(core_key[106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][11] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(core_key[107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][12] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(core_key[108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][13] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(core_key[109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][14] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(core_key[110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][15] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(core_key[111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][16] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(core_key[112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][17] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(core_key[113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][18] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(core_key[114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][19] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(core_key[115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][1] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(core_key[97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][20] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(core_key[116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][21] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(core_key[117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][22] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(core_key[118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][23] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(core_key[119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][24] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(core_key[120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][25] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(core_key[121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][26] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(core_key[122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][27] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(core_key[123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][28] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(core_key[124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][29] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(core_key[125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][2] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(core_key[98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][30] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(core_key[126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][31] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(core_key[127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][3] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(core_key[99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][4] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(core_key[100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][5] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(core_key[101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][6] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(core_key[102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][7] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(core_key[103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][8] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(core_key[104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[4][9] 
       (.C(clk_i),
        .CE(\key_reg[4][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(core_key[105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][0] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(core_key[64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][10] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(core_key[74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][11] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(core_key[75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][12] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(core_key[76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][13] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(core_key[77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][14] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(core_key[78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][15] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(core_key[79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][16] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(core_key[80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][17] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(core_key[81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][18] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(core_key[82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][19] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(core_key[83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][1] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(core_key[65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][20] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(core_key[84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][21] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(core_key[85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][22] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(core_key[86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][23] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(core_key[87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][24] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(core_key[88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][25] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(core_key[89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][26] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(core_key[90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][27] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(core_key[91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][28] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(core_key[92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][29] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(core_key[93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][2] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(core_key[66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][30] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(core_key[94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][31] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(core_key[95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][3] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(core_key[67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][4] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(core_key[68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][5] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(core_key[69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][6] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(core_key[70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][7] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(core_key[71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][8] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(core_key[72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[5][9] 
       (.C(clk_i),
        .CE(\key_reg[5][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(core_key[73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][0] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(core_key[32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][10] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(core_key[42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][11] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(core_key[43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][12] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(core_key[44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][13] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(core_key[45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][14] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(core_key[46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][15] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(core_key[47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][16] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(core_key[48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][17] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(core_key[49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][18] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(core_key[50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][19] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(core_key[51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][1] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(core_key[33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][20] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(core_key[52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][21] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(core_key[53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][22] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(core_key[54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][23] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(core_key[55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][24] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(core_key[56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][25] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(core_key[57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][26] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(core_key[58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][27] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(core_key[59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][28] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(core_key[60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][29] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(core_key[61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][2] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(core_key[34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][30] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(core_key[62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][31] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(core_key[63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][3] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(core_key[35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][4] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(core_key[36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][5] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(core_key[37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][6] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(core_key[38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][7] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(core_key[39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][8] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(core_key[40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[6][9] 
       (.C(clk_i),
        .CE(\key_reg[6][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(core_key[41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][0] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(core_key[0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][10] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(core_key[10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][11] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(core_key[11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][12] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(core_key[12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][13] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(core_key[13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][14] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(core_key[14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][15] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(core_key[15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][16] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(core_key[16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][17] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(core_key[17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][18] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(core_key[18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][19] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(core_key[19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][1] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(core_key[1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][20] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(core_key[20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][21] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(core_key[21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][22] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(core_key[22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][23] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(core_key[23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][24] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(core_key[24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][25] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(core_key[25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][26] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(core_key[26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][27] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(core_key[27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][28] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(core_key[28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][29] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(core_key[29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][2] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(core_key[2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][30] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(core_key[30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][31] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(core_key[31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][3] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(core_key[3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][4] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(core_key[4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][5] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(core_key[5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][6] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(core_key[6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][7] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(core_key[7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][8] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(core_key[8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_reg_reg[7][9] 
       (.C(clk_i),
        .CE(\key_reg[7][31]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(core_key[9]));
  (* ORIG_CELL_NAME = "keylen_reg_reg" *) 
  FDCE #(
    .INIT(1'b0)) 
    keylen_reg_reg
       (.C(clk_i),
        .CE(config_we4_out),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(p_1_in[3]));
  (* ORIG_CELL_NAME = "keylen_reg_reg" *) 
  FDCE #(
    .INIT(1'b0)) 
    keylen_reg_reg_rep
       (.C(clk_i),
        .CE(config_we4_out),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(keylen_reg_reg_rep_n_0));
  (* ORIG_CELL_NAME = "keylen_reg_reg" *) 
  FDCE #(
    .INIT(1'b0)) 
    keylen_reg_reg_rep__0
       (.C(clk_i),
        .CE(config_we4_out),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(keylen_reg_reg_rep__0_n_0));
  LUT5 #(
    .INIT(32'h00000020)) 
    next_reg_i_1
       (.I0(init_reg_i_2_n_0),
        .I1(enable_i[4]),
        .I2(enable_i[1]),
        .I3(enable_i[3]),
        .I4(init_reg_i_3_n_0),
        .O(next_new1_out));
  FDCE #(
    .INIT(1'b0)) 
    next_reg_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(next_new1_out),
        .Q(p_1_in[1]));
  FDCE #(
    .INIT(1'b0)) 
    ready_reg_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_ready),
        .Q(ready_reg));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[0]),
        .Q(result_reg[0]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[100] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[100]),
        .Q(result_reg[100]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[101] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[101]),
        .Q(result_reg[101]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[102] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[102]),
        .Q(result_reg[102]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[103] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[103]),
        .Q(result_reg[103]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[104] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[104]),
        .Q(result_reg[104]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[105] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[105]),
        .Q(result_reg[105]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[106] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[106]),
        .Q(result_reg[106]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[107] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[107]),
        .Q(result_reg[107]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[108] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[108]),
        .Q(result_reg[108]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[109] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[109]),
        .Q(result_reg[109]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[10]),
        .Q(result_reg[10]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[110] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[110]),
        .Q(result_reg[110]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[111] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[111]),
        .Q(result_reg[111]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[112] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[112]),
        .Q(result_reg[112]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[113] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[113]),
        .Q(result_reg[113]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[114] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[114]),
        .Q(result_reg[114]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[115] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[115]),
        .Q(result_reg[115]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[116] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[116]),
        .Q(result_reg[116]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[117] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[117]),
        .Q(result_reg[117]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[118] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[118]),
        .Q(result_reg[118]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[119] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[119]),
        .Q(result_reg[119]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[11]),
        .Q(result_reg[11]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[120] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[120]),
        .Q(result_reg[120]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[121] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[121]),
        .Q(result_reg[121]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[122] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[122]),
        .Q(result_reg[122]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[123] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[123]),
        .Q(result_reg[123]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[124] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[124]),
        .Q(result_reg[124]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[125] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[125]),
        .Q(result_reg[125]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[126] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[126]),
        .Q(result_reg[126]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[127] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[127]),
        .Q(result_reg[127]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[12]),
        .Q(result_reg[12]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[13]),
        .Q(result_reg[13]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[14]),
        .Q(result_reg[14]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[15]),
        .Q(result_reg[15]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[16]),
        .Q(result_reg[16]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[17]),
        .Q(result_reg[17]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[18]),
        .Q(result_reg[18]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[19]),
        .Q(result_reg[19]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[1]),
        .Q(result_reg[1]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[20]),
        .Q(result_reg[20]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[21]),
        .Q(result_reg[21]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[22]),
        .Q(result_reg[22]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[23]),
        .Q(result_reg[23]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[24]),
        .Q(result_reg[24]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[25]),
        .Q(result_reg[25]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[26]),
        .Q(result_reg[26]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[27]),
        .Q(result_reg[27]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[28]),
        .Q(result_reg[28]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[29]),
        .Q(result_reg[29]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[2]),
        .Q(result_reg[2]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[30]),
        .Q(result_reg[30]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[31]),
        .Q(result_reg[31]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[32] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[32]),
        .Q(result_reg[32]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[33] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[33]),
        .Q(result_reg[33]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[34] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[34]),
        .Q(result_reg[34]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[35] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[35]),
        .Q(result_reg[35]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[36] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[36]),
        .Q(result_reg[36]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[37] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[37]),
        .Q(result_reg[37]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[38] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[38]),
        .Q(result_reg[38]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[39] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[39]),
        .Q(result_reg[39]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[3]),
        .Q(result_reg[3]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[40] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[40]),
        .Q(result_reg[40]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[41] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[41]),
        .Q(result_reg[41]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[42] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[42]),
        .Q(result_reg[42]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[43] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[43]),
        .Q(result_reg[43]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[44] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[44]),
        .Q(result_reg[44]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[45] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[45]),
        .Q(result_reg[45]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[46] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[46]),
        .Q(result_reg[46]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[47] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[47]),
        .Q(result_reg[47]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[48] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[48]),
        .Q(result_reg[48]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[49] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[49]),
        .Q(result_reg[49]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[4]),
        .Q(result_reg[4]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[50] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[50]),
        .Q(result_reg[50]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[51] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[51]),
        .Q(result_reg[51]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[52] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[52]),
        .Q(result_reg[52]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[53] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[53]),
        .Q(result_reg[53]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[54] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[54]),
        .Q(result_reg[54]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[55] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[55]),
        .Q(result_reg[55]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[56] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[56]),
        .Q(result_reg[56]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[57] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[57]),
        .Q(result_reg[57]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[58] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[58]),
        .Q(result_reg[58]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[59] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[59]),
        .Q(result_reg[59]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[5]),
        .Q(result_reg[5]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[60] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[60]),
        .Q(result_reg[60]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[61] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[61]),
        .Q(result_reg[61]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[62] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[62]),
        .Q(result_reg[62]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[63] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[63]),
        .Q(result_reg[63]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[64] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[64]),
        .Q(result_reg[64]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[65] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[65]),
        .Q(result_reg[65]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[66] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[66]),
        .Q(result_reg[66]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[67] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[67]),
        .Q(result_reg[67]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[68] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[68]),
        .Q(result_reg[68]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[69] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[69]),
        .Q(result_reg[69]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[6]),
        .Q(result_reg[6]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[70] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[70]),
        .Q(result_reg[70]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[71] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[71]),
        .Q(result_reg[71]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[72] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[72]),
        .Q(result_reg[72]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[73] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[73]),
        .Q(result_reg[73]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[74] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[74]),
        .Q(result_reg[74]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[75] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[75]),
        .Q(result_reg[75]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[76] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[76]),
        .Q(result_reg[76]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[77] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[77]),
        .Q(result_reg[77]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[78] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[78]),
        .Q(result_reg[78]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[79] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[79]),
        .Q(result_reg[79]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[7]),
        .Q(result_reg[7]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[80] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[80]),
        .Q(result_reg[80]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[81] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[81]),
        .Q(result_reg[81]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[82] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[82]),
        .Q(result_reg[82]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[83] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[83]),
        .Q(result_reg[83]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[84] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[84]),
        .Q(result_reg[84]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[85] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[85]),
        .Q(result_reg[85]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[86] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[86]),
        .Q(result_reg[86]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[87] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[87]),
        .Q(result_reg[87]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[88] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[88]),
        .Q(result_reg[88]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[89] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[89]),
        .Q(result_reg[89]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[8]),
        .Q(result_reg[8]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[90] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[90]),
        .Q(result_reg[90]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[91] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[91]),
        .Q(result_reg[91]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[92] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[92]),
        .Q(result_reg[92]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[93] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[93]),
        .Q(result_reg[93]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[94] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[94]),
        .Q(result_reg[94]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[95] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[95]),
        .Q(result_reg[95]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[96] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[96]),
        .Q(result_reg[96]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[97] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[97]),
        .Q(result_reg[97]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[98] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[98]),
        .Q(result_reg[98]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[99] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[99]),
        .Q(result_reg[99]));
  FDCE #(
    .INIT(1'b0)) 
    \result_reg_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_result[9]),
        .Q(result_reg[9]));
  FDCE #(
    .INIT(1'b0)) 
    valid_reg_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(core_valid),
        .Q(valid_reg));
endmodule

(* ORIG_REF_NAME = "aes_core" *) 
module switch_elements_aes_core
   (ready,
    core_valid,
    D,
    p_1_in,
    core_block,
    core_key,
    clk_i,
    rst_i,
    \key_mem_reg[14][36] ,
    \key_mem_reg[14][127] );
  output ready;
  output core_valid;
  output [127:0]D;
  input [3:0]p_1_in;
  input [127:0]core_block;
  input [255:0]core_key;
  input clk_i;
  input rst_i;
  input \key_mem_reg[14][36] ;
  input \key_mem_reg[14][127] ;

  wire [127:0]D;
  wire [87:1]addroundkey_return;
  wire [1:0]aes_core_ctrl_new;
  wire [1:0]aes_core_ctrl_reg;
  wire clk_i;
  wire [127:0]core_block;
  wire [255:0]core_key;
  wire core_valid;
  wire dec_block_n_128;
  wire [127:0]dec_new_block;
  wire dec_ready;
  wire [3:0]dec_round_nr;
  wire enc_block_n_0;
  wire enc_block_n_1;
  wire enc_block_n_100;
  wire enc_block_n_101;
  wire enc_block_n_102;
  wire enc_block_n_103;
  wire enc_block_n_104;
  wire enc_block_n_105;
  wire enc_block_n_106;
  wire enc_block_n_107;
  wire enc_block_n_108;
  wire enc_block_n_109;
  wire enc_block_n_110;
  wire enc_block_n_111;
  wire enc_block_n_112;
  wire enc_block_n_113;
  wire enc_block_n_114;
  wire enc_block_n_115;
  wire enc_block_n_116;
  wire enc_block_n_117;
  wire enc_block_n_118;
  wire enc_block_n_119;
  wire enc_block_n_120;
  wire enc_block_n_121;
  wire enc_block_n_122;
  wire enc_block_n_123;
  wire enc_block_n_124;
  wire enc_block_n_125;
  wire enc_block_n_126;
  wire enc_block_n_127;
  wire enc_block_n_128;
  wire enc_block_n_129;
  wire enc_block_n_130;
  wire enc_block_n_131;
  wire enc_block_n_132;
  wire enc_block_n_133;
  wire enc_block_n_134;
  wire enc_block_n_135;
  wire enc_block_n_136;
  wire enc_block_n_137;
  wire enc_block_n_138;
  wire enc_block_n_139;
  wire enc_block_n_140;
  wire enc_block_n_141;
  wire enc_block_n_142;
  wire enc_block_n_143;
  wire enc_block_n_144;
  wire enc_block_n_145;
  wire enc_block_n_146;
  wire enc_block_n_147;
  wire enc_block_n_148;
  wire enc_block_n_149;
  wire enc_block_n_150;
  wire enc_block_n_22;
  wire enc_block_n_23;
  wire enc_block_n_24;
  wire enc_block_n_25;
  wire enc_block_n_26;
  wire enc_block_n_27;
  wire enc_block_n_28;
  wire enc_block_n_281;
  wire enc_block_n_282;
  wire enc_block_n_283;
  wire enc_block_n_284;
  wire enc_block_n_285;
  wire enc_block_n_286;
  wire enc_block_n_287;
  wire enc_block_n_288;
  wire enc_block_n_289;
  wire enc_block_n_29;
  wire enc_block_n_30;
  wire enc_block_n_31;
  wire enc_block_n_32;
  wire enc_block_n_33;
  wire enc_block_n_34;
  wire enc_block_n_35;
  wire enc_block_n_36;
  wire enc_block_n_37;
  wire enc_block_n_38;
  wire enc_block_n_39;
  wire enc_block_n_40;
  wire enc_block_n_41;
  wire enc_block_n_42;
  wire enc_block_n_43;
  wire enc_block_n_44;
  wire enc_block_n_45;
  wire enc_block_n_46;
  wire enc_block_n_47;
  wire enc_block_n_48;
  wire enc_block_n_49;
  wire enc_block_n_50;
  wire enc_block_n_51;
  wire enc_block_n_52;
  wire enc_block_n_53;
  wire enc_block_n_54;
  wire enc_block_n_55;
  wire enc_block_n_56;
  wire enc_block_n_57;
  wire enc_block_n_58;
  wire enc_block_n_59;
  wire enc_block_n_60;
  wire enc_block_n_61;
  wire enc_block_n_62;
  wire enc_block_n_63;
  wire enc_block_n_64;
  wire enc_block_n_65;
  wire enc_block_n_66;
  wire enc_block_n_67;
  wire enc_block_n_68;
  wire enc_block_n_69;
  wire enc_block_n_70;
  wire enc_block_n_71;
  wire enc_block_n_72;
  wire enc_block_n_73;
  wire enc_block_n_74;
  wire enc_block_n_75;
  wire enc_block_n_76;
  wire enc_block_n_77;
  wire enc_block_n_78;
  wire enc_block_n_79;
  wire enc_block_n_80;
  wire enc_block_n_81;
  wire enc_block_n_82;
  wire enc_block_n_83;
  wire enc_block_n_84;
  wire enc_block_n_85;
  wire enc_block_n_86;
  wire enc_block_n_87;
  wire enc_block_n_88;
  wire enc_block_n_89;
  wire enc_block_n_90;
  wire enc_block_n_91;
  wire enc_block_n_92;
  wire enc_block_n_93;
  wire enc_block_n_94;
  wire enc_block_n_95;
  wire enc_block_n_96;
  wire enc_block_n_97;
  wire enc_block_n_98;
  wire enc_block_n_99;
  wire enc_ready;
  wire init_state;
  wire [7:0]inv_mixcolumns_return0110_out__47;
  wire [7:1]inv_mixcolumns_return0117_out__50;
  wire [7:0]inv_mixcolumns_return0124_out__47;
  wire [7:1]inv_mixcolumns_return0134_out__63;
  wire [7:0]inv_mixcolumns_return0142_out__55;
  wire [7:1]inv_mixcolumns_return0149_out__55;
  wire [7:0]inv_mixcolumns_return0156_out__63;
  wire [7:1]inv_mixcolumns_return0166_out__55;
  wire [7:0]inv_mixcolumns_return0174_out__63;
  wire [7:1]inv_mixcolumns_return0181_out__58;
  wire [7:0]inv_mixcolumns_return0188_out__55;
  wire [7:1]inv_mixcolumns_return0198_out__63;
  wire [7:0]inv_mixcolumns_return0206_out__55;
  wire [7:1]inv_mixcolumns_return0213_out__55;
  wire [7:0]inv_mixcolumns_return0220_out__63;
  wire [7:1]inv_mixcolumns_return0__55;
  wire \key_mem_reg[14][127] ;
  wire \key_mem_reg[14][36] ;
  wire key_ready;
  wire keymem_n_0;
  wire keymem_n_1;
  wire keymem_n_10;
  wire keymem_n_100;
  wire keymem_n_101;
  wire keymem_n_102;
  wire keymem_n_103;
  wire keymem_n_104;
  wire keymem_n_105;
  wire keymem_n_107;
  wire keymem_n_108;
  wire keymem_n_109;
  wire keymem_n_11;
  wire keymem_n_110;
  wire keymem_n_111;
  wire keymem_n_112;
  wire keymem_n_12;
  wire keymem_n_13;
  wire keymem_n_14;
  wire keymem_n_15;
  wire keymem_n_16;
  wire keymem_n_17;
  wire keymem_n_18;
  wire keymem_n_19;
  wire keymem_n_2;
  wire keymem_n_20;
  wire keymem_n_21;
  wire keymem_n_23;
  wire keymem_n_24;
  wire keymem_n_241;
  wire keymem_n_242;
  wire keymem_n_243;
  wire keymem_n_244;
  wire keymem_n_245;
  wire keymem_n_246;
  wire keymem_n_247;
  wire keymem_n_25;
  wire keymem_n_26;
  wire keymem_n_27;
  wire keymem_n_28;
  wire keymem_n_288;
  wire keymem_n_289;
  wire keymem_n_29;
  wire keymem_n_290;
  wire keymem_n_291;
  wire keymem_n_292;
  wire keymem_n_293;
  wire keymem_n_294;
  wire keymem_n_295;
  wire keymem_n_296;
  wire keymem_n_297;
  wire keymem_n_3;
  wire keymem_n_30;
  wire keymem_n_31;
  wire keymem_n_32;
  wire keymem_n_33;
  wire keymem_n_34;
  wire keymem_n_36;
  wire keymem_n_37;
  wire keymem_n_38;
  wire keymem_n_39;
  wire keymem_n_4;
  wire keymem_n_40;
  wire keymem_n_41;
  wire keymem_n_43;
  wire keymem_n_44;
  wire keymem_n_45;
  wire keymem_n_46;
  wire keymem_n_47;
  wire keymem_n_48;
  wire keymem_n_49;
  wire keymem_n_5;
  wire keymem_n_51;
  wire keymem_n_52;
  wire keymem_n_53;
  wire keymem_n_54;
  wire keymem_n_55;
  wire keymem_n_56;
  wire keymem_n_57;
  wire keymem_n_58;
  wire keymem_n_59;
  wire keymem_n_6;
  wire keymem_n_60;
  wire keymem_n_61;
  wire keymem_n_62;
  wire keymem_n_64;
  wire keymem_n_65;
  wire keymem_n_66;
  wire keymem_n_67;
  wire keymem_n_68;
  wire keymem_n_69;
  wire keymem_n_71;
  wire keymem_n_72;
  wire keymem_n_73;
  wire keymem_n_74;
  wire keymem_n_75;
  wire keymem_n_76;
  wire keymem_n_77;
  wire keymem_n_79;
  wire keymem_n_8;
  wire keymem_n_80;
  wire keymem_n_81;
  wire keymem_n_82;
  wire keymem_n_83;
  wire keymem_n_84;
  wire keymem_n_85;
  wire keymem_n_86;
  wire keymem_n_87;
  wire keymem_n_88;
  wire keymem_n_89;
  wire keymem_n_9;
  wire keymem_n_90;
  wire keymem_n_92;
  wire keymem_n_93;
  wire keymem_n_94;
  wire keymem_n_95;
  wire keymem_n_96;
  wire keymem_n_97;
  wire keymem_n_98;
  wire keymem_n_99;
  wire [31:0]keymem_sboxw;
  wire [3:0]muxed_round_nr;
  wire [31:6]muxed_sboxw;
  wire [31:0]new_sboxw;
  wire [16:0]new_sboxw_0;
  wire [1:1]op126_in;
  wire [0:0]op127_in;
  wire [1:1]op158_in;
  wire [0:0]op159_in;
  wire [0:0]op191_in;
  wire [0:0]op96_in;
  wire [1:1]p_0_in31_in;
  wire [1:1]p_0_in38_in;
  wire [1:1]p_0_in46_in;
  wire [1:1]p_0_in54_in;
  wire [127:24]p_0_out;
  wire [31:24]p_19_in;
  wire [3:0]p_1_in;
  wire [31:24]rconw;
  wire ready;
  wire ready_new;
  wire ready_we;
  wire [127:0]round_key;
  wire rst_i;
  wire [0:0]update_type__0;

  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \FSM_sequential_aes_core_ctrl_reg[0]_i_1 
       (.I0(p_1_in[0]),
        .I1(aes_core_ctrl_reg[0]),
        .I2(aes_core_ctrl_reg[1]),
        .O(aes_core_ctrl_new[0]));
  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \FSM_sequential_aes_core_ctrl_reg[1]_i_2 
       (.I0(p_1_in[0]),
        .I1(p_1_in[1]),
        .I2(aes_core_ctrl_reg[0]),
        .I3(aes_core_ctrl_reg[1]),
        .O(aes_core_ctrl_new[1]));
  (* FSM_ENCODED_STATES = "CTRL_INIT:01,CTRL_IDLE:00,CTRL_NEXT:10" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_aes_core_ctrl_reg_reg[0] 
       (.C(clk_i),
        .CE(ready_we),
        .CLR(rst_i),
        .D(aes_core_ctrl_new[0]),
        .Q(aes_core_ctrl_reg[0]));
  (* FSM_ENCODED_STATES = "CTRL_INIT:01,CTRL_IDLE:00,CTRL_NEXT:10" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_aes_core_ctrl_reg_reg[1] 
       (.C(clk_i),
        .CE(ready_we),
        .CLR(rst_i),
        .D(aes_core_ctrl_new[1]),
        .Q(aes_core_ctrl_reg[1]));
  switch_elements_aes_decipher_block dec_block
       (.\FSM_sequential_dec_ctrl_reg_reg[0]_0 (update_type__0),
        .\FSM_sequential_dec_ctrl_reg_reg[1]_0 (dec_block_n_128),
        .Q(dec_round_nr),
        .addroundkey_return({addroundkey_return[87:81],addroundkey_return[71:65],addroundkey_return[47:40],addroundkey_return[23:17],addroundkey_return[15:1]}),
        .\block_w0_reg_reg[0]_0 (keymem_n_244),
        .\block_w0_reg_reg[0]_1 (keymem_n_288),
        .\block_w0_reg_reg[10]_0 (keymem_n_17),
        .\block_w0_reg_reg[12]_0 (keymem_n_16),
        .\block_w0_reg_reg[13]_0 (keymem_n_15),
        .\block_w0_reg_reg[14]_0 (keymem_n_14),
        .\block_w0_reg_reg[15]_0 (keymem_n_13),
        .\block_w0_reg_reg[16]_0 (keymem_n_247),
        .\block_w0_reg_reg[16]_1 (keymem_n_294),
        .\block_w0_reg_reg[17]_0 (keymem_n_12),
        .\block_w0_reg_reg[19]_0 (keymem_n_11),
        .\block_w0_reg_reg[1]_0 (keymem_n_27),
        .\block_w0_reg_reg[20]_0 (keymem_n_10),
        .\block_w0_reg_reg[21]_0 (keymem_n_9),
        .\block_w0_reg_reg[22]_0 (keymem_n_8),
        .\block_w0_reg_reg[23]_0 (keymem_n_6),
        .\block_w0_reg_reg[24]_0 (keymem_n_5),
        .\block_w0_reg_reg[25]_0 (keymem_n_4),
        .\block_w0_reg_reg[28]_0 (keymem_n_3),
        .\block_w0_reg_reg[29]_0 (keymem_n_2),
        .\block_w0_reg_reg[2]_0 (keymem_n_26),
        .\block_w0_reg_reg[30]_0 (keymem_n_1),
        .\block_w0_reg_reg[31]_0 (keymem_n_0),
        .\block_w0_reg_reg[3]_0 (keymem_n_25),
        .\block_w0_reg_reg[4]_0 (keymem_n_24),
        .\block_w0_reg_reg[5]_0 (keymem_n_23),
        .\block_w0_reg_reg[6]_0 (keymem_n_21),
        .\block_w0_reg_reg[7]_0 (keymem_n_20),
        .\block_w0_reg_reg[8]_0 (keymem_n_19),
        .\block_w0_reg_reg[9]_0 (keymem_n_18),
        .\block_w1_reg_reg[0]_0 (keymem_n_246),
        .\block_w1_reg_reg[0]_1 (keymem_n_289),
        .\block_w1_reg_reg[10]_0 (keymem_n_46),
        .\block_w1_reg_reg[12]_0 (keymem_n_45),
        .\block_w1_reg_reg[13]_0 (keymem_n_44),
        .\block_w1_reg_reg[14]_0 (keymem_n_43),
        .\block_w1_reg_reg[15]_0 (keymem_n_41),
        .\block_w1_reg_reg[16]_0 (keymem_n_241),
        .\block_w1_reg_reg[16]_1 (keymem_n_295),
        .\block_w1_reg_reg[17]_0 (keymem_n_40),
        .\block_w1_reg_reg[19]_0 (keymem_n_39),
        .\block_w1_reg_reg[1]_0 (keymem_n_55),
        .\block_w1_reg_reg[20]_0 (keymem_n_38),
        .\block_w1_reg_reg[21]_0 (keymem_n_37),
        .\block_w1_reg_reg[22]_0 (keymem_n_36),
        .\block_w1_reg_reg[23]_0 (keymem_n_34),
        .\block_w1_reg_reg[24]_0 (keymem_n_33),
        .\block_w1_reg_reg[25]_0 (keymem_n_32),
        .\block_w1_reg_reg[28]_0 (keymem_n_31),
        .\block_w1_reg_reg[29]_0 (keymem_n_30),
        .\block_w1_reg_reg[2]_0 (keymem_n_54),
        .\block_w1_reg_reg[30]_0 (keymem_n_29),
        .\block_w1_reg_reg[31]_0 (keymem_n_28),
        .\block_w1_reg_reg[3]_0 (keymem_n_53),
        .\block_w1_reg_reg[4]_0 (keymem_n_52),
        .\block_w1_reg_reg[5]_0 (keymem_n_51),
        .\block_w1_reg_reg[6]_0 (keymem_n_49),
        .\block_w1_reg_reg[7]_0 (keymem_n_48),
        .\block_w1_reg_reg[8]_0 (keymem_n_47),
        .\block_w1_reg_reg[9]_0 (keymem_n_292),
        .\block_w2_reg_reg[0]_0 (keymem_n_112),
        .\block_w2_reg_reg[0]_1 (keymem_n_290),
        .\block_w2_reg_reg[10]_0 (keymem_n_74),
        .\block_w2_reg_reg[12]_0 (keymem_n_73),
        .\block_w2_reg_reg[13]_0 (keymem_n_72),
        .\block_w2_reg_reg[14]_0 (keymem_n_71),
        .\block_w2_reg_reg[15]_0 (keymem_n_69),
        .\block_w2_reg_reg[16]_0 (keymem_n_243),
        .\block_w2_reg_reg[16]_1 (keymem_n_296),
        .\block_w2_reg_reg[17]_0 (keymem_n_68),
        .\block_w2_reg_reg[19]_0 (keymem_n_67),
        .\block_w2_reg_reg[1]_0 (keymem_n_83),
        .\block_w2_reg_reg[20]_0 (keymem_n_66),
        .\block_w2_reg_reg[21]_0 (keymem_n_65),
        .\block_w2_reg_reg[22]_0 (keymem_n_64),
        .\block_w2_reg_reg[23]_0 (keymem_n_62),
        .\block_w2_reg_reg[24]_0 (keymem_n_61),
        .\block_w2_reg_reg[25]_0 (keymem_n_60),
        .\block_w2_reg_reg[28]_0 (keymem_n_59),
        .\block_w2_reg_reg[29]_0 (keymem_n_58),
        .\block_w2_reg_reg[2]_0 (keymem_n_82),
        .\block_w2_reg_reg[30]_0 (keymem_n_57),
        .\block_w2_reg_reg[31]_0 (keymem_n_56),
        .\block_w2_reg_reg[3]_0 (keymem_n_81),
        .\block_w2_reg_reg[4]_0 (keymem_n_80),
        .\block_w2_reg_reg[5]_0 (keymem_n_79),
        .\block_w2_reg_reg[6]_0 (keymem_n_77),
        .\block_w2_reg_reg[7]_0 (keymem_n_76),
        .\block_w2_reg_reg[8]_0 (keymem_n_75),
        .\block_w2_reg_reg[9]_0 (keymem_n_293),
        .\block_w3_reg_reg[0]_0 (keymem_n_242),
        .\block_w3_reg_reg[0]_1 (keymem_n_291),
        .\block_w3_reg_reg[10]_0 (keymem_n_101),
        .\block_w3_reg_reg[12]_0 (keymem_n_100),
        .\block_w3_reg_reg[13]_0 (keymem_n_99),
        .\block_w3_reg_reg[14]_0 (keymem_n_98),
        .\block_w3_reg_reg[15]_0 (keymem_n_97),
        .\block_w3_reg_reg[16]_0 (keymem_n_245),
        .\block_w3_reg_reg[16]_1 (keymem_n_297),
        .\block_w3_reg_reg[17]_0 (keymem_n_96),
        .\block_w3_reg_reg[19]_0 (keymem_n_95),
        .\block_w3_reg_reg[1]_0 (keymem_n_111),
        .\block_w3_reg_reg[20]_0 (keymem_n_94),
        .\block_w3_reg_reg[21]_0 (keymem_n_93),
        .\block_w3_reg_reg[22]_0 (keymem_n_92),
        .\block_w3_reg_reg[23]_0 (keymem_n_90),
        .\block_w3_reg_reg[24]_0 (keymem_n_89),
        .\block_w3_reg_reg[25]_0 (keymem_n_88),
        .\block_w3_reg_reg[28]_0 (keymem_n_87),
        .\block_w3_reg_reg[29]_0 (keymem_n_86),
        .\block_w3_reg_reg[2]_0 (keymem_n_110),
        .\block_w3_reg_reg[30]_0 (keymem_n_85),
        .\block_w3_reg_reg[31]_0 (keymem_n_84),
        .\block_w3_reg_reg[3]_0 (keymem_n_109),
        .\block_w3_reg_reg[4]_0 (keymem_n_108),
        .\block_w3_reg_reg[5]_0 (keymem_n_107),
        .\block_w3_reg_reg[6]_0 (keymem_n_105),
        .\block_w3_reg_reg[7]_0 (keymem_n_104),
        .\block_w3_reg_reg[8]_0 (keymem_n_103),
        .\block_w3_reg_reg[9]_0 (keymem_n_102),
        .clk_i(clk_i),
        .dec_new_block(dec_new_block),
        .dec_ready(dec_ready),
        .inv_mixcolumns_return0110_out__47({inv_mixcolumns_return0110_out__47[7:2],inv_mixcolumns_return0110_out__47[0]}),
        .inv_mixcolumns_return0117_out__50(inv_mixcolumns_return0117_out__50),
        .inv_mixcolumns_return0124_out__47(inv_mixcolumns_return0124_out__47),
        .inv_mixcolumns_return0134_out__63(inv_mixcolumns_return0134_out__63),
        .inv_mixcolumns_return0142_out__55(inv_mixcolumns_return0142_out__55),
        .inv_mixcolumns_return0149_out__55(inv_mixcolumns_return0149_out__55),
        .inv_mixcolumns_return0156_out__63(inv_mixcolumns_return0156_out__63),
        .inv_mixcolumns_return0166_out__55(inv_mixcolumns_return0166_out__55),
        .inv_mixcolumns_return0174_out__63(inv_mixcolumns_return0174_out__63),
        .inv_mixcolumns_return0181_out__58(inv_mixcolumns_return0181_out__58),
        .inv_mixcolumns_return0188_out__55(inv_mixcolumns_return0188_out__55),
        .inv_mixcolumns_return0198_out__63(inv_mixcolumns_return0198_out__63),
        .inv_mixcolumns_return0206_out__55({inv_mixcolumns_return0206_out__55[7:2],inv_mixcolumns_return0206_out__55[0]}),
        .inv_mixcolumns_return0213_out__55(inv_mixcolumns_return0213_out__55),
        .inv_mixcolumns_return0220_out__63(inv_mixcolumns_return0220_out__63),
        .inv_mixcolumns_return0__55(inv_mixcolumns_return0__55),
        .\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11 ({new_sboxw_0[16],new_sboxw_0[9],new_sboxw_0[0]}),
        .op126_in(op126_in),
        .op127_in(op127_in),
        .op158_in(op158_in),
        .op159_in(op159_in),
        .op191_in(op191_in),
        .op96_in(op96_in),
        .p_0_in31_in(p_0_in31_in),
        .p_0_in38_in(p_0_in38_in),
        .p_0_in46_in(p_0_in46_in),
        .p_0_in54_in(p_0_in54_in),
        .p_0_out({p_0_out[127:113],p_0_out[111:97],p_0_out[95:88],p_0_out[79:72],p_0_out[63:49],p_0_out[39:33],p_0_out[31:24]}),
        .p_1_in(p_1_in[3:1]),
        .round_key({round_key[123:122],round_key[114],round_key[107],round_key[91:90],round_key[82],round_key[75],round_key[59:58],round_key[50],round_key[43],round_key[27:26],round_key[18],round_key[11]}),
        .rst_i(rst_i));
  switch_elements_aes_encipher_block enc_block
       (.D(D),
        .E(ready_we),
        .Q(keymem_sboxw),
        .addroundkey_return({addroundkey_return[84:83],addroundkey_return[81],addroundkey_return[68:67],addroundkey_return[65],addroundkey_return[44:43],addroundkey_return[41],addroundkey_return[20:19],addroundkey_return[17],addroundkey_return[12:11],addroundkey_return[9],addroundkey_return[4:3],addroundkey_return[1]}),
        .\block_w2_reg[28]_i_3 (dec_round_nr),
        .clk_i(clk_i),
        .core_block({core_block[127:125],core_block[122],core_block[120:117],core_block[114],core_block[112:109],core_block[106],core_block[104:101],core_block[98],core_block[96:93],core_block[90],core_block[88:85],core_block[82],core_block[80:77],core_block[74],core_block[72:69],core_block[66],core_block[64:61],core_block[58],core_block[56:53],core_block[50],core_block[48:45],core_block[42],core_block[40:37],core_block[34],core_block[32:29],core_block[26],core_block[24:21],core_block[18],core_block[16:13],core_block[10],core_block[8:5],core_block[2],core_block[0]}),
        .core_valid(core_valid),
        .dec_new_block(dec_new_block),
        .dec_ready(dec_ready),
        .enc_ready(enc_ready),
        .init_state(init_state),
        .key_ready(key_ready),
        .muxed_round_nr(muxed_round_nr),
        .new_sboxw(new_sboxw),
        .next_reg_reg(enc_block_n_150),
        .p_0_out({p_0_out[124:123],p_0_out[121],p_0_out[116:115],p_0_out[113],p_0_out[108:107],p_0_out[105],p_0_out[100:99],p_0_out[97],p_0_out[92:91],p_0_out[89],p_0_out[76:75],p_0_out[73],p_0_out[60:59],p_0_out[57],p_0_out[52:51],p_0_out[49],p_0_out[36:35],p_0_out[33],p_0_out[28:27],p_0_out[25]}),
        .p_19_in(p_19_in),
        .p_1_in(p_1_in),
        .\prev_key1_reg[127]_i_5 (rconw),
        .\prev_key1_reg_reg[0] (enc_block_n_22),
        .\prev_key1_reg_reg[0]_0 (enc_block_n_23),
        .\prev_key1_reg_reg[0]_1 (enc_block_n_24),
        .\prev_key1_reg_reg[0]_10 (enc_block_n_33),
        .\prev_key1_reg_reg[0]_11 (enc_block_n_34),
        .\prev_key1_reg_reg[0]_12 (enc_block_n_35),
        .\prev_key1_reg_reg[0]_13 (enc_block_n_36),
        .\prev_key1_reg_reg[0]_14 (enc_block_n_37),
        .\prev_key1_reg_reg[0]_15 (enc_block_n_38),
        .\prev_key1_reg_reg[0]_16 (enc_block_n_39),
        .\prev_key1_reg_reg[0]_17 (enc_block_n_40),
        .\prev_key1_reg_reg[0]_18 (enc_block_n_41),
        .\prev_key1_reg_reg[0]_19 (enc_block_n_42),
        .\prev_key1_reg_reg[0]_2 (enc_block_n_25),
        .\prev_key1_reg_reg[0]_20 (enc_block_n_43),
        .\prev_key1_reg_reg[0]_21 (enc_block_n_44),
        .\prev_key1_reg_reg[0]_22 (enc_block_n_45),
        .\prev_key1_reg_reg[0]_23 (enc_block_n_46),
        .\prev_key1_reg_reg[0]_24 (enc_block_n_47),
        .\prev_key1_reg_reg[0]_25 (enc_block_n_48),
        .\prev_key1_reg_reg[0]_26 (enc_block_n_49),
        .\prev_key1_reg_reg[0]_27 (enc_block_n_50),
        .\prev_key1_reg_reg[0]_28 (enc_block_n_51),
        .\prev_key1_reg_reg[0]_29 (enc_block_n_52),
        .\prev_key1_reg_reg[0]_3 (enc_block_n_26),
        .\prev_key1_reg_reg[0]_30 (enc_block_n_53),
        .\prev_key1_reg_reg[0]_4 (enc_block_n_27),
        .\prev_key1_reg_reg[0]_5 (enc_block_n_28),
        .\prev_key1_reg_reg[0]_6 (enc_block_n_29),
        .\prev_key1_reg_reg[0]_7 (enc_block_n_30),
        .\prev_key1_reg_reg[0]_8 (enc_block_n_31),
        .\prev_key1_reg_reg[0]_9 (enc_block_n_32),
        .\prev_key1_reg_reg[16] (enc_block_n_86),
        .\prev_key1_reg_reg[16]_0 (enc_block_n_87),
        .\prev_key1_reg_reg[16]_1 (enc_block_n_88),
        .\prev_key1_reg_reg[16]_10 (enc_block_n_97),
        .\prev_key1_reg_reg[16]_11 (enc_block_n_98),
        .\prev_key1_reg_reg[16]_12 (enc_block_n_99),
        .\prev_key1_reg_reg[16]_13 (enc_block_n_100),
        .\prev_key1_reg_reg[16]_14 (enc_block_n_101),
        .\prev_key1_reg_reg[16]_15 (enc_block_n_102),
        .\prev_key1_reg_reg[16]_16 (enc_block_n_103),
        .\prev_key1_reg_reg[16]_17 (enc_block_n_104),
        .\prev_key1_reg_reg[16]_18 (enc_block_n_105),
        .\prev_key1_reg_reg[16]_19 (enc_block_n_106),
        .\prev_key1_reg_reg[16]_2 (enc_block_n_89),
        .\prev_key1_reg_reg[16]_20 (enc_block_n_107),
        .\prev_key1_reg_reg[16]_21 (enc_block_n_108),
        .\prev_key1_reg_reg[16]_22 (enc_block_n_109),
        .\prev_key1_reg_reg[16]_23 (enc_block_n_110),
        .\prev_key1_reg_reg[16]_24 (enc_block_n_111),
        .\prev_key1_reg_reg[16]_25 (enc_block_n_112),
        .\prev_key1_reg_reg[16]_26 (enc_block_n_113),
        .\prev_key1_reg_reg[16]_27 (enc_block_n_114),
        .\prev_key1_reg_reg[16]_28 (enc_block_n_115),
        .\prev_key1_reg_reg[16]_29 (enc_block_n_116),
        .\prev_key1_reg_reg[16]_3 (enc_block_n_90),
        .\prev_key1_reg_reg[16]_30 (enc_block_n_117),
        .\prev_key1_reg_reg[16]_4 (enc_block_n_91),
        .\prev_key1_reg_reg[16]_5 (enc_block_n_92),
        .\prev_key1_reg_reg[16]_6 (enc_block_n_93),
        .\prev_key1_reg_reg[16]_7 (enc_block_n_94),
        .\prev_key1_reg_reg[16]_8 (enc_block_n_95),
        .\prev_key1_reg_reg[16]_9 (enc_block_n_96),
        .\prev_key1_reg_reg[24] (enc_block_n_118),
        .\prev_key1_reg_reg[24]_0 (enc_block_n_119),
        .\prev_key1_reg_reg[24]_1 (enc_block_n_120),
        .\prev_key1_reg_reg[24]_10 (enc_block_n_129),
        .\prev_key1_reg_reg[24]_11 (enc_block_n_130),
        .\prev_key1_reg_reg[24]_12 (enc_block_n_131),
        .\prev_key1_reg_reg[24]_13 (enc_block_n_132),
        .\prev_key1_reg_reg[24]_14 (enc_block_n_133),
        .\prev_key1_reg_reg[24]_15 (enc_block_n_134),
        .\prev_key1_reg_reg[24]_16 (enc_block_n_135),
        .\prev_key1_reg_reg[24]_17 (enc_block_n_136),
        .\prev_key1_reg_reg[24]_18 (enc_block_n_137),
        .\prev_key1_reg_reg[24]_19 (enc_block_n_138),
        .\prev_key1_reg_reg[24]_2 (enc_block_n_121),
        .\prev_key1_reg_reg[24]_20 (enc_block_n_139),
        .\prev_key1_reg_reg[24]_21 (enc_block_n_140),
        .\prev_key1_reg_reg[24]_22 (enc_block_n_141),
        .\prev_key1_reg_reg[24]_23 (enc_block_n_142),
        .\prev_key1_reg_reg[24]_24 (enc_block_n_143),
        .\prev_key1_reg_reg[24]_25 (enc_block_n_144),
        .\prev_key1_reg_reg[24]_26 (enc_block_n_145),
        .\prev_key1_reg_reg[24]_27 (enc_block_n_146),
        .\prev_key1_reg_reg[24]_28 (enc_block_n_147),
        .\prev_key1_reg_reg[24]_29 (enc_block_n_148),
        .\prev_key1_reg_reg[24]_3 (enc_block_n_122),
        .\prev_key1_reg_reg[24]_30 (enc_block_n_149),
        .\prev_key1_reg_reg[24]_4 (enc_block_n_123),
        .\prev_key1_reg_reg[24]_5 (enc_block_n_124),
        .\prev_key1_reg_reg[24]_6 (enc_block_n_125),
        .\prev_key1_reg_reg[24]_7 (enc_block_n_126),
        .\prev_key1_reg_reg[24]_8 (enc_block_n_127),
        .\prev_key1_reg_reg[24]_9 (enc_block_n_128),
        .\prev_key1_reg_reg[31] ({muxed_sboxw[31:30],muxed_sboxw[23:22],muxed_sboxw[15:14],muxed_sboxw[7:6]}),
        .\prev_key1_reg_reg[8] (enc_block_n_54),
        .\prev_key1_reg_reg[8]_0 (enc_block_n_55),
        .\prev_key1_reg_reg[8]_1 (enc_block_n_56),
        .\prev_key1_reg_reg[8]_10 (enc_block_n_65),
        .\prev_key1_reg_reg[8]_11 (enc_block_n_66),
        .\prev_key1_reg_reg[8]_12 (enc_block_n_67),
        .\prev_key1_reg_reg[8]_13 (enc_block_n_68),
        .\prev_key1_reg_reg[8]_14 (enc_block_n_69),
        .\prev_key1_reg_reg[8]_15 (enc_block_n_70),
        .\prev_key1_reg_reg[8]_16 (enc_block_n_71),
        .\prev_key1_reg_reg[8]_17 (enc_block_n_72),
        .\prev_key1_reg_reg[8]_18 (enc_block_n_73),
        .\prev_key1_reg_reg[8]_19 (enc_block_n_74),
        .\prev_key1_reg_reg[8]_2 (enc_block_n_57),
        .\prev_key1_reg_reg[8]_20 (enc_block_n_75),
        .\prev_key1_reg_reg[8]_21 (enc_block_n_76),
        .\prev_key1_reg_reg[8]_22 (enc_block_n_77),
        .\prev_key1_reg_reg[8]_23 (enc_block_n_78),
        .\prev_key1_reg_reg[8]_24 (enc_block_n_79),
        .\prev_key1_reg_reg[8]_25 (enc_block_n_80),
        .\prev_key1_reg_reg[8]_26 (enc_block_n_81),
        .\prev_key1_reg_reg[8]_27 (enc_block_n_82),
        .\prev_key1_reg_reg[8]_28 (enc_block_n_83),
        .\prev_key1_reg_reg[8]_29 (enc_block_n_84),
        .\prev_key1_reg_reg[8]_3 (enc_block_n_58),
        .\prev_key1_reg_reg[8]_30 (enc_block_n_85),
        .\prev_key1_reg_reg[8]_4 (enc_block_n_59),
        .\prev_key1_reg_reg[8]_5 (enc_block_n_60),
        .\prev_key1_reg_reg[8]_6 (enc_block_n_61),
        .\prev_key1_reg_reg[8]_7 (enc_block_n_62),
        .\prev_key1_reg_reg[8]_8 (enc_block_n_63),
        .\prev_key1_reg_reg[8]_9 (enc_block_n_64),
        .result_valid_reg_reg(aes_core_ctrl_reg),
        .\round_ctr_reg_reg[0]_0 (enc_block_n_286),
        .\round_ctr_reg_reg[0]_1 (enc_block_n_287),
        .\round_ctr_reg_reg[0]_2 (enc_block_n_288),
        .\round_ctr_reg_reg[0]_3 (enc_block_n_289),
        .\round_ctr_reg_reg[1]_0 (enc_block_n_0),
        .\round_ctr_reg_reg[1]_1 (enc_block_n_1),
        .\round_ctr_reg_reg[1]_2 (enc_block_n_283),
        .\round_ctr_reg_reg[1]_3 (enc_block_n_284),
        .\round_ctr_reg_reg[1]_4 (enc_block_n_285),
        .\round_ctr_reg_reg[3]_0 (enc_block_n_281),
        .\round_ctr_reg_reg[3]_1 (enc_block_n_282),
        .round_key(round_key),
        .rst_i(rst_i));
  switch_elements_aes_key_mem keymem
       (.Q(keymem_sboxw),
        .addroundkey_return({addroundkey_return[87:81],addroundkey_return[71:65],addroundkey_return[47:40],addroundkey_return[23:17],addroundkey_return[15:1]}),
        .\block_reg_reg[0][0] (keymem_n_242),
        .\block_reg_reg[0][16] (keymem_n_241),
        .\block_reg_reg[1][0] (keymem_n_244),
        .\block_reg_reg[1][16] (keymem_n_243),
        .\block_reg_reg[2][0] (keymem_n_246),
        .\block_reg_reg[2][16] (keymem_n_245),
        .\block_reg_reg[3][0] (keymem_n_112),
        .\block_reg_reg[3][16] (keymem_n_247),
        .\block_w0_reg[31]_i_6__0_0 (enc_block_n_1),
        .\block_w0_reg[31]_i_6__0_1 (enc_block_n_288),
        .\block_w0_reg_reg[0] (p_0_in54_in),
        .\block_w0_reg_reg[0]_0 (keymem_n_295),
        .\block_w0_reg_reg[0]_1 (update_type__0),
        .\block_w0_reg_reg[10] (keymem_n_17),
        .\block_w0_reg_reg[12] (keymem_n_16),
        .\block_w0_reg_reg[13] (keymem_n_15),
        .\block_w0_reg_reg[14] (keymem_n_14),
        .\block_w0_reg_reg[15] (keymem_n_13),
        .\block_w0_reg_reg[16] (op191_in),
        .\block_w0_reg_reg[16]_0 ({new_sboxw_0[16],new_sboxw_0[9],new_sboxw_0[0]}),
        .\block_w0_reg_reg[17] (keymem_n_12),
        .\block_w0_reg_reg[19] (keymem_n_11),
        .\block_w0_reg_reg[1] (keymem_n_27),
        .\block_w0_reg_reg[20] (keymem_n_10),
        .\block_w0_reg_reg[21] (keymem_n_9),
        .\block_w0_reg_reg[22] (keymem_n_8),
        .\block_w0_reg_reg[23] (keymem_n_6),
        .\block_w0_reg_reg[24] (keymem_n_5),
        .\block_w0_reg_reg[25] (keymem_n_4),
        .\block_w0_reg_reg[28] (keymem_n_3),
        .\block_w0_reg_reg[29] (keymem_n_2),
        .\block_w0_reg_reg[2] (keymem_n_26),
        .\block_w0_reg_reg[30] (keymem_n_1),
        .\block_w0_reg_reg[31] (keymem_n_0),
        .\block_w0_reg_reg[31]_0 (keymem_n_291),
        .\block_w0_reg_reg[31]_1 (dec_block_n_128),
        .\block_w0_reg_reg[31]_2 (enc_block_n_281),
        .\block_w0_reg_reg[3] (keymem_n_25),
        .\block_w0_reg_reg[4] (keymem_n_24),
        .\block_w0_reg_reg[5] (keymem_n_23),
        .\block_w0_reg_reg[6] (keymem_n_21),
        .\block_w0_reg_reg[7] (keymem_n_20),
        .\block_w0_reg_reg[8] (keymem_n_19),
        .\block_w0_reg_reg[8]_0 (keymem_n_293),
        .\block_w0_reg_reg[9] (keymem_n_18),
        .\block_w1_reg[29]_i_4_0 (enc_block_n_283),
        .\block_w1_reg[29]_i_4_1 (enc_block_n_286),
        .\block_w1_reg_reg[0] (p_0_in46_in),
        .\block_w1_reg_reg[0]_0 (keymem_n_296),
        .\block_w1_reg_reg[10] (keymem_n_46),
        .\block_w1_reg_reg[12] (keymem_n_45),
        .\block_w1_reg_reg[13] (keymem_n_44),
        .\block_w1_reg_reg[14] (keymem_n_43),
        .\block_w1_reg_reg[15] (keymem_n_41),
        .\block_w1_reg_reg[16] (op159_in),
        .\block_w1_reg_reg[17] (keymem_n_40),
        .\block_w1_reg_reg[19] (keymem_n_39),
        .\block_w1_reg_reg[1] (keymem_n_55),
        .\block_w1_reg_reg[20] (keymem_n_38),
        .\block_w1_reg_reg[21] (keymem_n_37),
        .\block_w1_reg_reg[22] (keymem_n_36),
        .\block_w1_reg_reg[23] (keymem_n_34),
        .\block_w1_reg_reg[24] (keymem_n_33),
        .\block_w1_reg_reg[25] (keymem_n_32),
        .\block_w1_reg_reg[28] (keymem_n_31),
        .\block_w1_reg_reg[29] (keymem_n_30),
        .\block_w1_reg_reg[2] (keymem_n_54),
        .\block_w1_reg_reg[30] (keymem_n_29),
        .\block_w1_reg_reg[31] (keymem_n_28),
        .\block_w1_reg_reg[31]_0 (keymem_n_288),
        .\block_w1_reg_reg[3] (keymem_n_53),
        .\block_w1_reg_reg[4] (keymem_n_52),
        .\block_w1_reg_reg[5] (keymem_n_51),
        .\block_w1_reg_reg[6] (keymem_n_49),
        .\block_w1_reg_reg[7] (keymem_n_48),
        .\block_w1_reg_reg[8] (keymem_n_47),
        .\block_w1_reg_reg[9] (op158_in),
        .\block_w2_reg[29]_i_4_0 (enc_block_n_284),
        .\block_w2_reg[29]_i_4_1 (enc_block_n_287),
        .\block_w2_reg_reg[0] (p_0_in38_in),
        .\block_w2_reg_reg[0]_0 (keymem_n_297),
        .\block_w2_reg_reg[10] (keymem_n_74),
        .\block_w2_reg_reg[12] (keymem_n_73),
        .\block_w2_reg_reg[13] (keymem_n_72),
        .\block_w2_reg_reg[14] (keymem_n_71),
        .\block_w2_reg_reg[15] (keymem_n_69),
        .\block_w2_reg_reg[16] (op127_in),
        .\block_w2_reg_reg[17] (keymem_n_68),
        .\block_w2_reg_reg[19] (keymem_n_67),
        .\block_w2_reg_reg[1] (keymem_n_83),
        .\block_w2_reg_reg[20] (keymem_n_66),
        .\block_w2_reg_reg[21] (keymem_n_65),
        .\block_w2_reg_reg[22] (keymem_n_64),
        .\block_w2_reg_reg[23] (keymem_n_62),
        .\block_w2_reg_reg[24] (keymem_n_61),
        .\block_w2_reg_reg[25] (keymem_n_60),
        .\block_w2_reg_reg[28] (keymem_n_59),
        .\block_w2_reg_reg[29] (keymem_n_58),
        .\block_w2_reg_reg[2] (keymem_n_82),
        .\block_w2_reg_reg[30] (keymem_n_57),
        .\block_w2_reg_reg[31] (keymem_n_56),
        .\block_w2_reg_reg[31]_0 (keymem_n_289),
        .\block_w2_reg_reg[3] (keymem_n_81),
        .\block_w2_reg_reg[4] (keymem_n_80),
        .\block_w2_reg_reg[5] (keymem_n_79),
        .\block_w2_reg_reg[6] (keymem_n_77),
        .\block_w2_reg_reg[7] (keymem_n_76),
        .\block_w2_reg_reg[8] (keymem_n_75),
        .\block_w2_reg_reg[9] (op126_in),
        .\block_w3_reg[1]_i_4__0_0 (enc_block_n_0),
        .\block_w3_reg[30]_i_4_0 (enc_block_n_285),
        .\block_w3_reg[30]_i_4_1 (enc_block_n_289),
        .\block_w3_reg_reg[0] (p_0_in31_in),
        .\block_w3_reg_reg[0]_0 (keymem_n_294),
        .\block_w3_reg_reg[10] (keymem_n_101),
        .\block_w3_reg_reg[12] (keymem_n_100),
        .\block_w3_reg_reg[13] (keymem_n_99),
        .\block_w3_reg_reg[14] (keymem_n_98),
        .\block_w3_reg_reg[15] (keymem_n_97),
        .\block_w3_reg_reg[16] (op96_in),
        .\block_w3_reg_reg[17] (keymem_n_96),
        .\block_w3_reg_reg[19] (keymem_n_95),
        .\block_w3_reg_reg[1] (keymem_n_111),
        .\block_w3_reg_reg[20] (keymem_n_94),
        .\block_w3_reg_reg[21] (keymem_n_93),
        .\block_w3_reg_reg[22] (keymem_n_92),
        .\block_w3_reg_reg[23] (keymem_n_90),
        .\block_w3_reg_reg[24] (keymem_n_89),
        .\block_w3_reg_reg[25] (keymem_n_88),
        .\block_w3_reg_reg[26] (enc_block_n_282),
        .\block_w3_reg_reg[28] (keymem_n_87),
        .\block_w3_reg_reg[29] (keymem_n_86),
        .\block_w3_reg_reg[2] (keymem_n_110),
        .\block_w3_reg_reg[30] (keymem_n_85),
        .\block_w3_reg_reg[31] (keymem_n_84),
        .\block_w3_reg_reg[31]_0 (keymem_n_290),
        .\block_w3_reg_reg[3] (keymem_n_109),
        .\block_w3_reg_reg[4] (keymem_n_108),
        .\block_w3_reg_reg[5] (keymem_n_107),
        .\block_w3_reg_reg[6] (keymem_n_105),
        .\block_w3_reg_reg[7] (keymem_n_104),
        .\block_w3_reg_reg[8] (keymem_n_103),
        .\block_w3_reg_reg[8]_0 (keymem_n_292),
        .\block_w3_reg_reg[9] (keymem_n_102),
        .clk_i(clk_i),
        .core_block(core_block),
        .core_key(core_key),
        .dec_new_block(dec_new_block),
        .dec_ready(dec_ready),
        .enc_ready(enc_ready),
        .init_state(init_state),
        .inv_mixcolumns_return0110_out__47({inv_mixcolumns_return0110_out__47[7:2],inv_mixcolumns_return0110_out__47[0]}),
        .inv_mixcolumns_return0117_out__50(inv_mixcolumns_return0117_out__50),
        .inv_mixcolumns_return0124_out__47(inv_mixcolumns_return0124_out__47),
        .inv_mixcolumns_return0134_out__63(inv_mixcolumns_return0134_out__63),
        .inv_mixcolumns_return0142_out__55(inv_mixcolumns_return0142_out__55),
        .inv_mixcolumns_return0149_out__55(inv_mixcolumns_return0149_out__55),
        .inv_mixcolumns_return0156_out__63(inv_mixcolumns_return0156_out__63),
        .inv_mixcolumns_return0166_out__55(inv_mixcolumns_return0166_out__55),
        .inv_mixcolumns_return0174_out__63(inv_mixcolumns_return0174_out__63),
        .inv_mixcolumns_return0181_out__58(inv_mixcolumns_return0181_out__58),
        .inv_mixcolumns_return0188_out__55(inv_mixcolumns_return0188_out__55),
        .inv_mixcolumns_return0198_out__63(inv_mixcolumns_return0198_out__63),
        .inv_mixcolumns_return0206_out__55({inv_mixcolumns_return0206_out__55[7:2],inv_mixcolumns_return0206_out__55[0]}),
        .inv_mixcolumns_return0213_out__55(inv_mixcolumns_return0213_out__55),
        .inv_mixcolumns_return0220_out__63(inv_mixcolumns_return0220_out__63),
        .inv_mixcolumns_return0__55(inv_mixcolumns_return0__55),
        .\key_mem_reg[14][127]_0 (\key_mem_reg[14][127] ),
        .\key_mem_reg[14][36]_0 (\key_mem_reg[14][36] ),
        .key_ready(key_ready),
        .muxed_round_nr(muxed_round_nr),
        .new_sboxw(new_sboxw),
        .p_0_out({p_0_out[127:113],p_0_out[111:97],p_0_out[95:88],p_0_out[79:72],p_0_out[63:49],p_0_out[39:33],p_0_out[31:24]}),
        .p_19_in(p_19_in),
        .p_1_in({p_1_in[3:2],p_1_in[0]}),
        .\rcon_reg_reg[7]_0 (rconw),
        .ready_new(ready_new),
        .ready_reg_reg_0(aes_core_ctrl_reg),
        .round_key(round_key),
        .rst_i(rst_i));
  FDPE #(
    .INIT(1'b1)) 
    ready_reg_reg
       (.C(clk_i),
        .CE(ready_we),
        .D(ready_new),
        .PRE(rst_i),
        .Q(ready));
  FDCE #(
    .INIT(1'b0)) 
    result_valid_reg_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(enc_block_n_150),
        .Q(core_valid));
  switch_elements_aes_sbox sbox_inst
       (.\block_w2_reg_reg[0]_i_5_0 (enc_block_n_22),
        .\block_w2_reg_reg[0]_i_5_1 (enc_block_n_30),
        .\block_w2_reg_reg[0]_i_5_2 (enc_block_n_38),
        .\block_w2_reg_reg[0]_i_5_3 (enc_block_n_46),
        .\block_w2_reg_reg[1]_i_5_0 (enc_block_n_23),
        .\block_w2_reg_reg[1]_i_5_1 (enc_block_n_31),
        .\block_w2_reg_reg[1]_i_5_2 (enc_block_n_39),
        .\block_w2_reg_reg[1]_i_5_3 (enc_block_n_47),
        .\block_w2_reg_reg[2]_i_5_0 (enc_block_n_24),
        .\block_w2_reg_reg[2]_i_5_1 (enc_block_n_32),
        .\block_w2_reg_reg[2]_i_5_2 (enc_block_n_40),
        .\block_w2_reg_reg[2]_i_5_3 (enc_block_n_48),
        .\block_w2_reg_reg[3]_i_5_0 (enc_block_n_25),
        .\block_w2_reg_reg[3]_i_5_1 (enc_block_n_33),
        .\block_w2_reg_reg[3]_i_5_2 (enc_block_n_41),
        .\block_w2_reg_reg[3]_i_5_3 (enc_block_n_49),
        .\block_w2_reg_reg[4]_i_6_0 (enc_block_n_26),
        .\block_w2_reg_reg[4]_i_6_1 (enc_block_n_34),
        .\block_w2_reg_reg[4]_i_6_2 (enc_block_n_42),
        .\block_w2_reg_reg[4]_i_6_3 (enc_block_n_50),
        .\block_w2_reg_reg[5]_i_5_0 (enc_block_n_27),
        .\block_w2_reg_reg[5]_i_5_1 (enc_block_n_35),
        .\block_w2_reg_reg[5]_i_5_2 (enc_block_n_43),
        .\block_w2_reg_reg[5]_i_5_3 (enc_block_n_51),
        .\block_w2_reg_reg[6]_i_5_0 (enc_block_n_28),
        .\block_w2_reg_reg[6]_i_5_1 (enc_block_n_36),
        .\block_w2_reg_reg[6]_i_5_2 (enc_block_n_44),
        .\block_w2_reg_reg[6]_i_5_3 (enc_block_n_52),
        .\block_w2_reg_reg[7]_i_5_0 (enc_block_n_29),
        .\block_w2_reg_reg[7]_i_5_1 (enc_block_n_37),
        .\block_w2_reg_reg[7]_i_5_2 (enc_block_n_45),
        .\block_w2_reg_reg[7]_i_5_3 (enc_block_n_53),
        .\block_w3_reg[31]_i_3 ({muxed_sboxw[31:30],muxed_sboxw[23:22],muxed_sboxw[15:14],muxed_sboxw[7:6]}),
        .new_sboxw(new_sboxw),
        .\sbox_inferred__0/block_w2_reg_reg[10]_i_5_0 (enc_block_n_56),
        .\sbox_inferred__0/block_w2_reg_reg[10]_i_5_1 (enc_block_n_64),
        .\sbox_inferred__0/block_w2_reg_reg[10]_i_5_2 (enc_block_n_72),
        .\sbox_inferred__0/block_w2_reg_reg[10]_i_5_3 (enc_block_n_80),
        .\sbox_inferred__0/block_w2_reg_reg[11]_i_5_0 (enc_block_n_57),
        .\sbox_inferred__0/block_w2_reg_reg[11]_i_5_1 (enc_block_n_65),
        .\sbox_inferred__0/block_w2_reg_reg[11]_i_5_2 (enc_block_n_73),
        .\sbox_inferred__0/block_w2_reg_reg[11]_i_5_3 (enc_block_n_81),
        .\sbox_inferred__0/block_w2_reg_reg[12]_i_5_0 (enc_block_n_58),
        .\sbox_inferred__0/block_w2_reg_reg[12]_i_5_1 (enc_block_n_66),
        .\sbox_inferred__0/block_w2_reg_reg[12]_i_5_2 (enc_block_n_74),
        .\sbox_inferred__0/block_w2_reg_reg[12]_i_5_3 (enc_block_n_82),
        .\sbox_inferred__0/block_w2_reg_reg[13]_i_5_0 (enc_block_n_59),
        .\sbox_inferred__0/block_w2_reg_reg[13]_i_5_1 (enc_block_n_67),
        .\sbox_inferred__0/block_w2_reg_reg[13]_i_5_2 (enc_block_n_75),
        .\sbox_inferred__0/block_w2_reg_reg[13]_i_5_3 (enc_block_n_83),
        .\sbox_inferred__0/block_w2_reg_reg[14]_i_5_0 (enc_block_n_60),
        .\sbox_inferred__0/block_w2_reg_reg[14]_i_5_1 (enc_block_n_68),
        .\sbox_inferred__0/block_w2_reg_reg[14]_i_5_2 (enc_block_n_76),
        .\sbox_inferred__0/block_w2_reg_reg[14]_i_5_3 (enc_block_n_84),
        .\sbox_inferred__0/block_w2_reg_reg[15]_i_5_0 (enc_block_n_61),
        .\sbox_inferred__0/block_w2_reg_reg[15]_i_5_1 (enc_block_n_69),
        .\sbox_inferred__0/block_w2_reg_reg[15]_i_5_2 (enc_block_n_77),
        .\sbox_inferred__0/block_w2_reg_reg[15]_i_5_3 (enc_block_n_85),
        .\sbox_inferred__0/block_w2_reg_reg[8]_i_5_0 (enc_block_n_54),
        .\sbox_inferred__0/block_w2_reg_reg[8]_i_5_1 (enc_block_n_62),
        .\sbox_inferred__0/block_w2_reg_reg[8]_i_5_2 (enc_block_n_70),
        .\sbox_inferred__0/block_w2_reg_reg[8]_i_5_3 (enc_block_n_78),
        .\sbox_inferred__0/block_w2_reg_reg[9]_i_6_0 (enc_block_n_55),
        .\sbox_inferred__0/block_w2_reg_reg[9]_i_6_1 (enc_block_n_63),
        .\sbox_inferred__0/block_w2_reg_reg[9]_i_6_2 (enc_block_n_71),
        .\sbox_inferred__0/block_w2_reg_reg[9]_i_6_3 (enc_block_n_79),
        .\sbox_inferred__1/block_w2_reg_reg[16]_i_5_0 (enc_block_n_86),
        .\sbox_inferred__1/block_w2_reg_reg[16]_i_5_1 (enc_block_n_94),
        .\sbox_inferred__1/block_w2_reg_reg[16]_i_5_2 (enc_block_n_102),
        .\sbox_inferred__1/block_w2_reg_reg[16]_i_5_3 (enc_block_n_110),
        .\sbox_inferred__1/block_w2_reg_reg[17]_i_5_0 (enc_block_n_87),
        .\sbox_inferred__1/block_w2_reg_reg[17]_i_5_1 (enc_block_n_95),
        .\sbox_inferred__1/block_w2_reg_reg[17]_i_5_2 (enc_block_n_103),
        .\sbox_inferred__1/block_w2_reg_reg[17]_i_5_3 (enc_block_n_111),
        .\sbox_inferred__1/block_w2_reg_reg[18]_i_5_0 (enc_block_n_88),
        .\sbox_inferred__1/block_w2_reg_reg[18]_i_5_1 (enc_block_n_96),
        .\sbox_inferred__1/block_w2_reg_reg[18]_i_5_2 (enc_block_n_104),
        .\sbox_inferred__1/block_w2_reg_reg[18]_i_5_3 (enc_block_n_112),
        .\sbox_inferred__1/block_w2_reg_reg[19]_i_5_0 (enc_block_n_89),
        .\sbox_inferred__1/block_w2_reg_reg[19]_i_5_1 (enc_block_n_97),
        .\sbox_inferred__1/block_w2_reg_reg[19]_i_5_2 (enc_block_n_105),
        .\sbox_inferred__1/block_w2_reg_reg[19]_i_5_3 (enc_block_n_113),
        .\sbox_inferred__1/block_w2_reg_reg[20]_i_6_0 (enc_block_n_90),
        .\sbox_inferred__1/block_w2_reg_reg[20]_i_6_1 (enc_block_n_98),
        .\sbox_inferred__1/block_w2_reg_reg[20]_i_6_2 (enc_block_n_106),
        .\sbox_inferred__1/block_w2_reg_reg[20]_i_6_3 (enc_block_n_114),
        .\sbox_inferred__1/block_w2_reg_reg[21]_i_5_0 (enc_block_n_91),
        .\sbox_inferred__1/block_w2_reg_reg[21]_i_5_1 (enc_block_n_99),
        .\sbox_inferred__1/block_w2_reg_reg[21]_i_5_2 (enc_block_n_107),
        .\sbox_inferred__1/block_w2_reg_reg[21]_i_5_3 (enc_block_n_115),
        .\sbox_inferred__1/block_w2_reg_reg[22]_i_5_0 (enc_block_n_92),
        .\sbox_inferred__1/block_w2_reg_reg[22]_i_5_1 (enc_block_n_100),
        .\sbox_inferred__1/block_w2_reg_reg[22]_i_5_2 (enc_block_n_108),
        .\sbox_inferred__1/block_w2_reg_reg[22]_i_5_3 (enc_block_n_116),
        .\sbox_inferred__1/block_w2_reg_reg[23]_i_5_0 (enc_block_n_93),
        .\sbox_inferred__1/block_w2_reg_reg[23]_i_5_1 (enc_block_n_101),
        .\sbox_inferred__1/block_w2_reg_reg[23]_i_5_2 (enc_block_n_109),
        .\sbox_inferred__1/block_w2_reg_reg[23]_i_5_3 (enc_block_n_117),
        .\sbox_inferred__2/block_w2_reg_reg[24]_i_5_0 (enc_block_n_118),
        .\sbox_inferred__2/block_w2_reg_reg[24]_i_5_1 (enc_block_n_126),
        .\sbox_inferred__2/block_w2_reg_reg[24]_i_5_2 (enc_block_n_134),
        .\sbox_inferred__2/block_w2_reg_reg[24]_i_5_3 (enc_block_n_142),
        .\sbox_inferred__2/block_w2_reg_reg[25]_i_6_0 (enc_block_n_119),
        .\sbox_inferred__2/block_w2_reg_reg[25]_i_6_1 (enc_block_n_127),
        .\sbox_inferred__2/block_w2_reg_reg[25]_i_6_2 (enc_block_n_135),
        .\sbox_inferred__2/block_w2_reg_reg[25]_i_6_3 (enc_block_n_143),
        .\sbox_inferred__2/block_w2_reg_reg[26]_i_5_0 (enc_block_n_120),
        .\sbox_inferred__2/block_w2_reg_reg[26]_i_5_1 (enc_block_n_128),
        .\sbox_inferred__2/block_w2_reg_reg[26]_i_5_2 (enc_block_n_136),
        .\sbox_inferred__2/block_w2_reg_reg[26]_i_5_3 (enc_block_n_144),
        .\sbox_inferred__2/block_w2_reg_reg[27]_i_5_0 (enc_block_n_121),
        .\sbox_inferred__2/block_w2_reg_reg[27]_i_5_1 (enc_block_n_129),
        .\sbox_inferred__2/block_w2_reg_reg[27]_i_5_2 (enc_block_n_137),
        .\sbox_inferred__2/block_w2_reg_reg[27]_i_5_3 (enc_block_n_145),
        .\sbox_inferred__2/block_w2_reg_reg[28]_i_5_0 (enc_block_n_122),
        .\sbox_inferred__2/block_w2_reg_reg[28]_i_5_1 (enc_block_n_130),
        .\sbox_inferred__2/block_w2_reg_reg[28]_i_5_2 (enc_block_n_138),
        .\sbox_inferred__2/block_w2_reg_reg[28]_i_5_3 (enc_block_n_146),
        .\sbox_inferred__2/block_w2_reg_reg[29]_i_5_0 (enc_block_n_123),
        .\sbox_inferred__2/block_w2_reg_reg[29]_i_5_1 (enc_block_n_131),
        .\sbox_inferred__2/block_w2_reg_reg[29]_i_5_2 (enc_block_n_139),
        .\sbox_inferred__2/block_w2_reg_reg[29]_i_5_3 (enc_block_n_147),
        .\sbox_inferred__2/block_w2_reg_reg[30]_i_5_0 (enc_block_n_124),
        .\sbox_inferred__2/block_w2_reg_reg[30]_i_5_1 (enc_block_n_132),
        .\sbox_inferred__2/block_w2_reg_reg[30]_i_5_2 (enc_block_n_140),
        .\sbox_inferred__2/block_w2_reg_reg[30]_i_5_3 (enc_block_n_148),
        .\sbox_inferred__2/block_w2_reg_reg[31]_i_10_0 (enc_block_n_125),
        .\sbox_inferred__2/block_w2_reg_reg[31]_i_10_1 (enc_block_n_133),
        .\sbox_inferred__2/block_w2_reg_reg[31]_i_10_2 (enc_block_n_141),
        .\sbox_inferred__2/block_w2_reg_reg[31]_i_10_3 (enc_block_n_149));
endmodule

(* ORIG_REF_NAME = "aes_decipher_block" *) 
module switch_elements_aes_decipher_block
   (dec_new_block,
    \FSM_sequential_dec_ctrl_reg_reg[1]_0 ,
    Q,
    \FSM_sequential_dec_ctrl_reg_reg[0]_0 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11 ,
    dec_ready,
    round_key,
    \block_w3_reg_reg[16]_0 ,
    \block_w3_reg_reg[16]_1 ,
    op96_in,
    \block_w2_reg_reg[16]_0 ,
    \block_w2_reg_reg[16]_1 ,
    op127_in,
    \block_w1_reg_reg[16]_0 ,
    \block_w1_reg_reg[16]_1 ,
    op159_in,
    \block_w0_reg_reg[16]_0 ,
    \block_w0_reg_reg[16]_1 ,
    op191_in,
    \block_w2_reg_reg[9]_0 ,
    op126_in,
    \block_w1_reg_reg[9]_0 ,
    op158_in,
    \block_w3_reg_reg[0]_0 ,
    \block_w3_reg_reg[0]_1 ,
    p_0_in31_in,
    \block_w2_reg_reg[0]_0 ,
    \block_w2_reg_reg[0]_1 ,
    p_0_in38_in,
    \block_w1_reg_reg[0]_0 ,
    \block_w1_reg_reg[0]_1 ,
    p_0_in46_in,
    \block_w0_reg_reg[0]_0 ,
    \block_w0_reg_reg[0]_1 ,
    p_0_in54_in,
    \block_w0_reg_reg[1]_0 ,
    addroundkey_return,
    inv_mixcolumns_return0166_out__55,
    \block_w1_reg_reg[1]_0 ,
    p_0_out,
    inv_mixcolumns_return0134_out__63,
    \block_w2_reg_reg[1]_0 ,
    inv_mixcolumns_return0__55,
    \block_w3_reg_reg[1]_0 ,
    inv_mixcolumns_return0198_out__63,
    \block_w0_reg_reg[2]_0 ,
    \block_w1_reg_reg[2]_0 ,
    \block_w2_reg_reg[2]_0 ,
    \block_w3_reg_reg[2]_0 ,
    \block_w0_reg_reg[3]_0 ,
    \block_w1_reg_reg[3]_0 ,
    \block_w2_reg_reg[3]_0 ,
    \block_w3_reg_reg[3]_0 ,
    \block_w0_reg_reg[4]_0 ,
    \block_w1_reg_reg[4]_0 ,
    \block_w2_reg_reg[4]_0 ,
    \block_w3_reg_reg[4]_0 ,
    \block_w0_reg_reg[5]_0 ,
    \block_w1_reg_reg[5]_0 ,
    \block_w2_reg_reg[5]_0 ,
    \block_w3_reg_reg[5]_0 ,
    \block_w0_reg_reg[6]_0 ,
    \block_w1_reg_reg[6]_0 ,
    \block_w2_reg_reg[6]_0 ,
    \block_w3_reg_reg[6]_0 ,
    \block_w0_reg_reg[7]_0 ,
    \block_w1_reg_reg[7]_0 ,
    \block_w2_reg_reg[7]_0 ,
    \block_w3_reg_reg[7]_0 ,
    \block_w0_reg_reg[8]_0 ,
    inv_mixcolumns_return0142_out__55,
    \block_w1_reg_reg[8]_0 ,
    inv_mixcolumns_return0110_out__47,
    \block_w2_reg_reg[8]_0 ,
    inv_mixcolumns_return0206_out__55,
    \block_w3_reg_reg[8]_0 ,
    inv_mixcolumns_return0174_out__63,
    \block_w0_reg_reg[9]_0 ,
    \block_w3_reg_reg[9]_0 ,
    \block_w0_reg_reg[10]_0 ,
    \block_w1_reg_reg[10]_0 ,
    \block_w2_reg_reg[10]_0 ,
    \block_w3_reg_reg[10]_0 ,
    \block_w0_reg_reg[12]_0 ,
    \block_w1_reg_reg[12]_0 ,
    \block_w2_reg_reg[12]_0 ,
    \block_w3_reg_reg[12]_0 ,
    \block_w0_reg_reg[13]_0 ,
    \block_w1_reg_reg[13]_0 ,
    \block_w2_reg_reg[13]_0 ,
    \block_w3_reg_reg[13]_0 ,
    \block_w0_reg_reg[14]_0 ,
    \block_w1_reg_reg[14]_0 ,
    \block_w2_reg_reg[14]_0 ,
    \block_w3_reg_reg[14]_0 ,
    \block_w0_reg_reg[15]_0 ,
    \block_w1_reg_reg[15]_0 ,
    \block_w2_reg_reg[15]_0 ,
    \block_w3_reg_reg[15]_0 ,
    \block_w0_reg_reg[17]_0 ,
    inv_mixcolumns_return0117_out__50,
    \block_w1_reg_reg[17]_0 ,
    inv_mixcolumns_return0213_out__55,
    \block_w2_reg_reg[17]_0 ,
    inv_mixcolumns_return0181_out__58,
    \block_w3_reg_reg[17]_0 ,
    inv_mixcolumns_return0149_out__55,
    \block_w0_reg_reg[19]_0 ,
    \block_w1_reg_reg[19]_0 ,
    \block_w2_reg_reg[19]_0 ,
    \block_w3_reg_reg[19]_0 ,
    \block_w0_reg_reg[20]_0 ,
    \block_w1_reg_reg[20]_0 ,
    \block_w2_reg_reg[20]_0 ,
    \block_w3_reg_reg[20]_0 ,
    \block_w0_reg_reg[21]_0 ,
    \block_w1_reg_reg[21]_0 ,
    \block_w2_reg_reg[21]_0 ,
    \block_w3_reg_reg[21]_0 ,
    \block_w0_reg_reg[22]_0 ,
    \block_w1_reg_reg[22]_0 ,
    \block_w2_reg_reg[22]_0 ,
    \block_w3_reg_reg[22]_0 ,
    \block_w0_reg_reg[23]_0 ,
    \block_w1_reg_reg[23]_0 ,
    \block_w2_reg_reg[23]_0 ,
    \block_w3_reg_reg[23]_0 ,
    \block_w0_reg_reg[24]_0 ,
    inv_mixcolumns_return0220_out__63,
    \block_w1_reg_reg[24]_0 ,
    inv_mixcolumns_return0188_out__55,
    \block_w2_reg_reg[24]_0 ,
    inv_mixcolumns_return0156_out__63,
    \block_w3_reg_reg[24]_0 ,
    inv_mixcolumns_return0124_out__47,
    \block_w0_reg_reg[25]_0 ,
    \block_w1_reg_reg[25]_0 ,
    \block_w2_reg_reg[25]_0 ,
    \block_w3_reg_reg[25]_0 ,
    \block_w0_reg_reg[28]_0 ,
    \block_w1_reg_reg[28]_0 ,
    \block_w2_reg_reg[28]_0 ,
    \block_w3_reg_reg[28]_0 ,
    \block_w0_reg_reg[29]_0 ,
    \block_w1_reg_reg[29]_0 ,
    \block_w2_reg_reg[29]_0 ,
    \block_w3_reg_reg[29]_0 ,
    \block_w0_reg_reg[30]_0 ,
    \block_w1_reg_reg[30]_0 ,
    \block_w2_reg_reg[30]_0 ,
    \block_w3_reg_reg[30]_0 ,
    \block_w0_reg_reg[31]_0 ,
    \block_w1_reg_reg[31]_0 ,
    \block_w2_reg_reg[31]_0 ,
    \block_w3_reg_reg[31]_0 ,
    p_1_in,
    clk_i,
    rst_i);
  output [127:0]dec_new_block;
  output \FSM_sequential_dec_ctrl_reg_reg[1]_0 ;
  output [3:0]Q;
  output [0:0]\FSM_sequential_dec_ctrl_reg_reg[0]_0 ;
  output [2:0]\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11 ;
  output dec_ready;
  input [15:0]round_key;
  input \block_w3_reg_reg[16]_0 ;
  input \block_w3_reg_reg[16]_1 ;
  input [0:0]op96_in;
  input \block_w2_reg_reg[16]_0 ;
  input \block_w2_reg_reg[16]_1 ;
  input [0:0]op127_in;
  input \block_w1_reg_reg[16]_0 ;
  input \block_w1_reg_reg[16]_1 ;
  input [0:0]op159_in;
  input \block_w0_reg_reg[16]_0 ;
  input \block_w0_reg_reg[16]_1 ;
  input [0:0]op191_in;
  input \block_w2_reg_reg[9]_0 ;
  input [0:0]op126_in;
  input \block_w1_reg_reg[9]_0 ;
  input [0:0]op158_in;
  input \block_w3_reg_reg[0]_0 ;
  input \block_w3_reg_reg[0]_1 ;
  input [0:0]p_0_in31_in;
  input \block_w2_reg_reg[0]_0 ;
  input \block_w2_reg_reg[0]_1 ;
  input [0:0]p_0_in38_in;
  input \block_w1_reg_reg[0]_0 ;
  input \block_w1_reg_reg[0]_1 ;
  input [0:0]p_0_in46_in;
  input \block_w0_reg_reg[0]_0 ;
  input \block_w0_reg_reg[0]_1 ;
  input [0:0]p_0_in54_in;
  input \block_w0_reg_reg[1]_0 ;
  input [43:0]addroundkey_return;
  input [6:0]inv_mixcolumns_return0166_out__55;
  input \block_w1_reg_reg[1]_0 ;
  input [75:0]p_0_out;
  input [6:0]inv_mixcolumns_return0134_out__63;
  input \block_w2_reg_reg[1]_0 ;
  input [6:0]inv_mixcolumns_return0__55;
  input \block_w3_reg_reg[1]_0 ;
  input [6:0]inv_mixcolumns_return0198_out__63;
  input \block_w0_reg_reg[2]_0 ;
  input \block_w1_reg_reg[2]_0 ;
  input \block_w2_reg_reg[2]_0 ;
  input \block_w3_reg_reg[2]_0 ;
  input \block_w0_reg_reg[3]_0 ;
  input \block_w1_reg_reg[3]_0 ;
  input \block_w2_reg_reg[3]_0 ;
  input \block_w3_reg_reg[3]_0 ;
  input \block_w0_reg_reg[4]_0 ;
  input \block_w1_reg_reg[4]_0 ;
  input \block_w2_reg_reg[4]_0 ;
  input \block_w3_reg_reg[4]_0 ;
  input \block_w0_reg_reg[5]_0 ;
  input \block_w1_reg_reg[5]_0 ;
  input \block_w2_reg_reg[5]_0 ;
  input \block_w3_reg_reg[5]_0 ;
  input \block_w0_reg_reg[6]_0 ;
  input \block_w1_reg_reg[6]_0 ;
  input \block_w2_reg_reg[6]_0 ;
  input \block_w3_reg_reg[6]_0 ;
  input \block_w0_reg_reg[7]_0 ;
  input \block_w1_reg_reg[7]_0 ;
  input \block_w2_reg_reg[7]_0 ;
  input \block_w3_reg_reg[7]_0 ;
  input \block_w0_reg_reg[8]_0 ;
  input [7:0]inv_mixcolumns_return0142_out__55;
  input \block_w1_reg_reg[8]_0 ;
  input [6:0]inv_mixcolumns_return0110_out__47;
  input \block_w2_reg_reg[8]_0 ;
  input [6:0]inv_mixcolumns_return0206_out__55;
  input \block_w3_reg_reg[8]_0 ;
  input [7:0]inv_mixcolumns_return0174_out__63;
  input \block_w0_reg_reg[9]_0 ;
  input \block_w3_reg_reg[9]_0 ;
  input \block_w0_reg_reg[10]_0 ;
  input \block_w1_reg_reg[10]_0 ;
  input \block_w2_reg_reg[10]_0 ;
  input \block_w3_reg_reg[10]_0 ;
  input \block_w0_reg_reg[12]_0 ;
  input \block_w1_reg_reg[12]_0 ;
  input \block_w2_reg_reg[12]_0 ;
  input \block_w3_reg_reg[12]_0 ;
  input \block_w0_reg_reg[13]_0 ;
  input \block_w1_reg_reg[13]_0 ;
  input \block_w2_reg_reg[13]_0 ;
  input \block_w3_reg_reg[13]_0 ;
  input \block_w0_reg_reg[14]_0 ;
  input \block_w1_reg_reg[14]_0 ;
  input \block_w2_reg_reg[14]_0 ;
  input \block_w3_reg_reg[14]_0 ;
  input \block_w0_reg_reg[15]_0 ;
  input \block_w1_reg_reg[15]_0 ;
  input \block_w2_reg_reg[15]_0 ;
  input \block_w3_reg_reg[15]_0 ;
  input \block_w0_reg_reg[17]_0 ;
  input [6:0]inv_mixcolumns_return0117_out__50;
  input \block_w1_reg_reg[17]_0 ;
  input [6:0]inv_mixcolumns_return0213_out__55;
  input \block_w2_reg_reg[17]_0 ;
  input [6:0]inv_mixcolumns_return0181_out__58;
  input \block_w3_reg_reg[17]_0 ;
  input [6:0]inv_mixcolumns_return0149_out__55;
  input \block_w0_reg_reg[19]_0 ;
  input \block_w1_reg_reg[19]_0 ;
  input \block_w2_reg_reg[19]_0 ;
  input \block_w3_reg_reg[19]_0 ;
  input \block_w0_reg_reg[20]_0 ;
  input \block_w1_reg_reg[20]_0 ;
  input \block_w2_reg_reg[20]_0 ;
  input \block_w3_reg_reg[20]_0 ;
  input \block_w0_reg_reg[21]_0 ;
  input \block_w1_reg_reg[21]_0 ;
  input \block_w2_reg_reg[21]_0 ;
  input \block_w3_reg_reg[21]_0 ;
  input \block_w0_reg_reg[22]_0 ;
  input \block_w1_reg_reg[22]_0 ;
  input \block_w2_reg_reg[22]_0 ;
  input \block_w3_reg_reg[22]_0 ;
  input \block_w0_reg_reg[23]_0 ;
  input \block_w1_reg_reg[23]_0 ;
  input \block_w2_reg_reg[23]_0 ;
  input \block_w3_reg_reg[23]_0 ;
  input \block_w0_reg_reg[24]_0 ;
  input [7:0]inv_mixcolumns_return0220_out__63;
  input \block_w1_reg_reg[24]_0 ;
  input [7:0]inv_mixcolumns_return0188_out__55;
  input \block_w2_reg_reg[24]_0 ;
  input [7:0]inv_mixcolumns_return0156_out__63;
  input \block_w3_reg_reg[24]_0 ;
  input [7:0]inv_mixcolumns_return0124_out__47;
  input \block_w0_reg_reg[25]_0 ;
  input \block_w1_reg_reg[25]_0 ;
  input \block_w2_reg_reg[25]_0 ;
  input \block_w3_reg_reg[25]_0 ;
  input \block_w0_reg_reg[28]_0 ;
  input \block_w1_reg_reg[28]_0 ;
  input \block_w2_reg_reg[28]_0 ;
  input \block_w3_reg_reg[28]_0 ;
  input \block_w0_reg_reg[29]_0 ;
  input \block_w1_reg_reg[29]_0 ;
  input \block_w2_reg_reg[29]_0 ;
  input \block_w3_reg_reg[29]_0 ;
  input \block_w0_reg_reg[30]_0 ;
  input \block_w1_reg_reg[30]_0 ;
  input \block_w2_reg_reg[30]_0 ;
  input \block_w3_reg_reg[30]_0 ;
  input \block_w0_reg_reg[31]_0 ;
  input \block_w1_reg_reg[31]_0 ;
  input \block_w2_reg_reg[31]_0 ;
  input \block_w3_reg_reg[31]_0 ;
  input [2:0]p_1_in;
  input clk_i;
  input rst_i;

  wire \FSM_sequential_dec_ctrl_reg[1]_i_1_n_0 ;
  wire \FSM_sequential_dec_ctrl_reg[1]_i_3_n_0 ;
  wire [0:0]\FSM_sequential_dec_ctrl_reg_reg[0]_0 ;
  wire \FSM_sequential_dec_ctrl_reg_reg[1]_0 ;
  wire [3:0]Q;
  wire [43:0]addroundkey_return;
  wire \block_w0_reg[0]_i_1_n_0 ;
  wire \block_w0_reg[10]_i_3_n_0 ;
  wire \block_w0_reg[11]_i_2__0_n_0 ;
  wire \block_w0_reg[11]_i_3_n_0 ;
  wire \block_w0_reg[12]_i_3_n_0 ;
  wire \block_w0_reg[13]_i_3_n_0 ;
  wire \block_w0_reg[14]_i_3_n_0 ;
  wire \block_w0_reg[15]_i_3_n_0 ;
  wire \block_w0_reg[16]_i_1_n_0 ;
  wire \block_w0_reg[17]_i_3_n_0 ;
  wire \block_w0_reg[18]_i_2__0_n_0 ;
  wire \block_w0_reg[18]_i_3_n_0 ;
  wire \block_w0_reg[19]_i_3_n_0 ;
  wire \block_w0_reg[1]_i_3_n_0 ;
  wire \block_w0_reg[20]_i_3_n_0 ;
  wire \block_w0_reg[21]_i_3_n_0 ;
  wire \block_w0_reg[22]_i_3_n_0 ;
  wire \block_w0_reg[23]_i_3_n_0 ;
  wire \block_w0_reg[24]_i_3_n_0 ;
  wire \block_w0_reg[25]_i_3_n_0 ;
  wire \block_w0_reg[26]_i_2__0_n_0 ;
  wire \block_w0_reg[26]_i_3_n_0 ;
  wire \block_w0_reg[27]_i_2__0_n_0 ;
  wire \block_w0_reg[27]_i_3_n_0 ;
  wire \block_w0_reg[28]_i_3_n_0 ;
  wire \block_w0_reg[29]_i_3_n_0 ;
  wire \block_w0_reg[2]_i_3_n_0 ;
  wire \block_w0_reg[30]_i_3_n_0 ;
  wire \block_w0_reg[31]_i_4_n_0 ;
  wire \block_w0_reg[3]_i_3_n_0 ;
  wire \block_w0_reg[4]_i_3_n_0 ;
  wire \block_w0_reg[5]_i_3_n_0 ;
  wire \block_w0_reg[6]_i_3_n_0 ;
  wire \block_w0_reg[7]_i_3_n_0 ;
  wire \block_w0_reg[8]_i_3_n_0 ;
  wire \block_w0_reg[9]_i_3_n_0 ;
  wire \block_w0_reg_reg[0]_0 ;
  wire \block_w0_reg_reg[0]_1 ;
  wire \block_w0_reg_reg[10]_0 ;
  wire \block_w0_reg_reg[10]_i_1_n_0 ;
  wire \block_w0_reg_reg[11]_i_1_n_0 ;
  wire \block_w0_reg_reg[12]_0 ;
  wire \block_w0_reg_reg[12]_i_1_n_0 ;
  wire \block_w0_reg_reg[13]_0 ;
  wire \block_w0_reg_reg[13]_i_1_n_0 ;
  wire \block_w0_reg_reg[14]_0 ;
  wire \block_w0_reg_reg[14]_i_1_n_0 ;
  wire \block_w0_reg_reg[15]_0 ;
  wire \block_w0_reg_reg[15]_i_1_n_0 ;
  wire \block_w0_reg_reg[16]_0 ;
  wire \block_w0_reg_reg[16]_1 ;
  wire \block_w0_reg_reg[17]_0 ;
  wire \block_w0_reg_reg[17]_i_1_n_0 ;
  wire \block_w0_reg_reg[18]_i_1_n_0 ;
  wire \block_w0_reg_reg[19]_0 ;
  wire \block_w0_reg_reg[19]_i_1_n_0 ;
  wire \block_w0_reg_reg[1]_0 ;
  wire \block_w0_reg_reg[1]_i_1_n_0 ;
  wire \block_w0_reg_reg[20]_0 ;
  wire \block_w0_reg_reg[20]_i_1_n_0 ;
  wire \block_w0_reg_reg[21]_0 ;
  wire \block_w0_reg_reg[21]_i_1_n_0 ;
  wire \block_w0_reg_reg[22]_0 ;
  wire \block_w0_reg_reg[22]_i_1_n_0 ;
  wire \block_w0_reg_reg[23]_0 ;
  wire \block_w0_reg_reg[23]_i_1_n_0 ;
  wire \block_w0_reg_reg[24]_0 ;
  wire \block_w0_reg_reg[24]_i_1_n_0 ;
  wire \block_w0_reg_reg[25]_0 ;
  wire \block_w0_reg_reg[25]_i_1_n_0 ;
  wire \block_w0_reg_reg[26]_i_1_n_0 ;
  wire \block_w0_reg_reg[27]_i_1_n_0 ;
  wire \block_w0_reg_reg[28]_0 ;
  wire \block_w0_reg_reg[28]_i_1_n_0 ;
  wire \block_w0_reg_reg[29]_0 ;
  wire \block_w0_reg_reg[29]_i_1_n_0 ;
  wire \block_w0_reg_reg[2]_0 ;
  wire \block_w0_reg_reg[2]_i_1_n_0 ;
  wire \block_w0_reg_reg[30]_0 ;
  wire \block_w0_reg_reg[30]_i_1_n_0 ;
  wire \block_w0_reg_reg[31]_0 ;
  wire \block_w0_reg_reg[31]_i_2_n_0 ;
  wire \block_w0_reg_reg[3]_0 ;
  wire \block_w0_reg_reg[3]_i_1_n_0 ;
  wire \block_w0_reg_reg[4]_0 ;
  wire \block_w0_reg_reg[4]_i_1_n_0 ;
  wire \block_w0_reg_reg[5]_0 ;
  wire \block_w0_reg_reg[5]_i_1_n_0 ;
  wire \block_w0_reg_reg[6]_0 ;
  wire \block_w0_reg_reg[6]_i_1_n_0 ;
  wire \block_w0_reg_reg[7]_0 ;
  wire \block_w0_reg_reg[7]_i_1_n_0 ;
  wire \block_w0_reg_reg[8]_0 ;
  wire \block_w0_reg_reg[8]_i_1_n_0 ;
  wire \block_w0_reg_reg[9]_0 ;
  wire \block_w0_reg_reg[9]_i_1_n_0 ;
  wire block_w0_we;
  wire \block_w1_reg[0]_i_1_n_0 ;
  wire \block_w1_reg[10]_i_3_n_0 ;
  wire \block_w1_reg[11]_i_2__0_n_0 ;
  wire \block_w1_reg[11]_i_3_n_0 ;
  wire \block_w1_reg[12]_i_3_n_0 ;
  wire \block_w1_reg[13]_i_3_n_0 ;
  wire \block_w1_reg[14]_i_3_n_0 ;
  wire \block_w1_reg[15]_i_3_n_0 ;
  wire \block_w1_reg[16]_i_1_n_0 ;
  wire \block_w1_reg[17]_i_3_n_0 ;
  wire \block_w1_reg[18]_i_2__0_n_0 ;
  wire \block_w1_reg[18]_i_3_n_0 ;
  wire \block_w1_reg[19]_i_3_n_0 ;
  wire \block_w1_reg[1]_i_3_n_0 ;
  wire \block_w1_reg[20]_i_3_n_0 ;
  wire \block_w1_reg[21]_i_3_n_0 ;
  wire \block_w1_reg[22]_i_3_n_0 ;
  wire \block_w1_reg[23]_i_3_n_0 ;
  wire \block_w1_reg[24]_i_3_n_0 ;
  wire \block_w1_reg[25]_i_3_n_0 ;
  wire \block_w1_reg[26]_i_2__0_n_0 ;
  wire \block_w1_reg[26]_i_3_n_0 ;
  wire \block_w1_reg[27]_i_2__0_n_0 ;
  wire \block_w1_reg[27]_i_3_n_0 ;
  wire \block_w1_reg[28]_i_3_n_0 ;
  wire \block_w1_reg[29]_i_3_n_0 ;
  wire \block_w1_reg[2]_i_3_n_0 ;
  wire \block_w1_reg[30]_i_3_n_0 ;
  wire \block_w1_reg[31]_i_4_n_0 ;
  wire \block_w1_reg[3]_i_3_n_0 ;
  wire \block_w1_reg[4]_i_3_n_0 ;
  wire \block_w1_reg[5]_i_3_n_0 ;
  wire \block_w1_reg[6]_i_3_n_0 ;
  wire \block_w1_reg[7]_i_3_n_0 ;
  wire \block_w1_reg[8]_i_3_n_0 ;
  wire \block_w1_reg[9]_i_1_n_0 ;
  wire \block_w1_reg[9]_i_2__0_n_0 ;
  wire \block_w1_reg_reg[0]_0 ;
  wire \block_w1_reg_reg[0]_1 ;
  wire \block_w1_reg_reg[10]_0 ;
  wire \block_w1_reg_reg[10]_i_1_n_0 ;
  wire \block_w1_reg_reg[11]_i_1_n_0 ;
  wire \block_w1_reg_reg[12]_0 ;
  wire \block_w1_reg_reg[12]_i_1_n_0 ;
  wire \block_w1_reg_reg[13]_0 ;
  wire \block_w1_reg_reg[13]_i_1_n_0 ;
  wire \block_w1_reg_reg[14]_0 ;
  wire \block_w1_reg_reg[14]_i_1_n_0 ;
  wire \block_w1_reg_reg[15]_0 ;
  wire \block_w1_reg_reg[15]_i_1_n_0 ;
  wire \block_w1_reg_reg[16]_0 ;
  wire \block_w1_reg_reg[16]_1 ;
  wire \block_w1_reg_reg[17]_0 ;
  wire \block_w1_reg_reg[17]_i_1_n_0 ;
  wire \block_w1_reg_reg[18]_i_1_n_0 ;
  wire \block_w1_reg_reg[19]_0 ;
  wire \block_w1_reg_reg[19]_i_1_n_0 ;
  wire \block_w1_reg_reg[1]_0 ;
  wire \block_w1_reg_reg[1]_i_1_n_0 ;
  wire \block_w1_reg_reg[20]_0 ;
  wire \block_w1_reg_reg[20]_i_1_n_0 ;
  wire \block_w1_reg_reg[21]_0 ;
  wire \block_w1_reg_reg[21]_i_1_n_0 ;
  wire \block_w1_reg_reg[22]_0 ;
  wire \block_w1_reg_reg[22]_i_1_n_0 ;
  wire \block_w1_reg_reg[23]_0 ;
  wire \block_w1_reg_reg[23]_i_1_n_0 ;
  wire \block_w1_reg_reg[24]_0 ;
  wire \block_w1_reg_reg[24]_i_1_n_0 ;
  wire \block_w1_reg_reg[25]_0 ;
  wire \block_w1_reg_reg[25]_i_1_n_0 ;
  wire \block_w1_reg_reg[26]_i_1_n_0 ;
  wire \block_w1_reg_reg[27]_i_1_n_0 ;
  wire \block_w1_reg_reg[28]_0 ;
  wire \block_w1_reg_reg[28]_i_1_n_0 ;
  wire \block_w1_reg_reg[29]_0 ;
  wire \block_w1_reg_reg[29]_i_1_n_0 ;
  wire \block_w1_reg_reg[2]_0 ;
  wire \block_w1_reg_reg[2]_i_1_n_0 ;
  wire \block_w1_reg_reg[30]_0 ;
  wire \block_w1_reg_reg[30]_i_1_n_0 ;
  wire \block_w1_reg_reg[31]_0 ;
  wire \block_w1_reg_reg[31]_i_2_n_0 ;
  wire \block_w1_reg_reg[3]_0 ;
  wire \block_w1_reg_reg[3]_i_1_n_0 ;
  wire \block_w1_reg_reg[4]_0 ;
  wire \block_w1_reg_reg[4]_i_1_n_0 ;
  wire \block_w1_reg_reg[5]_0 ;
  wire \block_w1_reg_reg[5]_i_1_n_0 ;
  wire \block_w1_reg_reg[6]_0 ;
  wire \block_w1_reg_reg[6]_i_1_n_0 ;
  wire \block_w1_reg_reg[7]_0 ;
  wire \block_w1_reg_reg[7]_i_1_n_0 ;
  wire \block_w1_reg_reg[8]_0 ;
  wire \block_w1_reg_reg[8]_i_1_n_0 ;
  wire \block_w1_reg_reg[9]_0 ;
  wire block_w1_we;
  wire \block_w2_reg[10]_i_3_n_0 ;
  wire \block_w2_reg[11]_i_2__0_n_0 ;
  wire \block_w2_reg[11]_i_3_n_0 ;
  wire \block_w2_reg[12]_i_3_n_0 ;
  wire \block_w2_reg[13]_i_3_n_0 ;
  wire \block_w2_reg[14]_i_3_n_0 ;
  wire \block_w2_reg[15]_i_3_n_0 ;
  wire \block_w2_reg[17]_i_3_n_0 ;
  wire \block_w2_reg[18]_i_2__0_n_0 ;
  wire \block_w2_reg[18]_i_3_n_0 ;
  wire \block_w2_reg[19]_i_3_n_0 ;
  wire \block_w2_reg[1]_i_3_n_0 ;
  wire \block_w2_reg[20]_i_3_n_0 ;
  wire \block_w2_reg[21]_i_3_n_0 ;
  wire \block_w2_reg[22]_i_3_n_0 ;
  wire \block_w2_reg[23]_i_3_n_0 ;
  wire \block_w2_reg[24]_i_3_n_0 ;
  wire \block_w2_reg[25]_i_3_n_0 ;
  wire \block_w2_reg[26]_i_2__0_n_0 ;
  wire \block_w2_reg[26]_i_3_n_0 ;
  wire \block_w2_reg[27]_i_2__0_n_0 ;
  wire \block_w2_reg[27]_i_3_n_0 ;
  wire \block_w2_reg[28]_i_3_n_0 ;
  wire \block_w2_reg[29]_i_3_n_0 ;
  wire \block_w2_reg[2]_i_3_n_0 ;
  wire \block_w2_reg[30]_i_3_n_0 ;
  wire \block_w2_reg[31]_i_4_n_0 ;
  wire \block_w2_reg[3]_i_3_n_0 ;
  wire \block_w2_reg[4]_i_3_n_0 ;
  wire \block_w2_reg[5]_i_3_n_0 ;
  wire \block_w2_reg[6]_i_3_n_0 ;
  wire \block_w2_reg[7]_i_3_n_0 ;
  wire \block_w2_reg[8]_i_3_n_0 ;
  wire \block_w2_reg[9]_i_2_n_0 ;
  wire \block_w2_reg_reg[0]_0 ;
  wire \block_w2_reg_reg[0]_1 ;
  wire \block_w2_reg_reg[10]_0 ;
  wire \block_w2_reg_reg[12]_0 ;
  wire \block_w2_reg_reg[13]_0 ;
  wire \block_w2_reg_reg[14]_0 ;
  wire \block_w2_reg_reg[15]_0 ;
  wire \block_w2_reg_reg[16]_0 ;
  wire \block_w2_reg_reg[16]_1 ;
  wire \block_w2_reg_reg[17]_0 ;
  wire \block_w2_reg_reg[19]_0 ;
  wire \block_w2_reg_reg[1]_0 ;
  wire \block_w2_reg_reg[20]_0 ;
  wire \block_w2_reg_reg[21]_0 ;
  wire \block_w2_reg_reg[22]_0 ;
  wire \block_w2_reg_reg[23]_0 ;
  wire \block_w2_reg_reg[24]_0 ;
  wire \block_w2_reg_reg[25]_0 ;
  wire \block_w2_reg_reg[28]_0 ;
  wire \block_w2_reg_reg[29]_0 ;
  wire \block_w2_reg_reg[2]_0 ;
  wire \block_w2_reg_reg[30]_0 ;
  wire \block_w2_reg_reg[31]_0 ;
  wire \block_w2_reg_reg[3]_0 ;
  wire \block_w2_reg_reg[4]_0 ;
  wire \block_w2_reg_reg[5]_0 ;
  wire \block_w2_reg_reg[6]_0 ;
  wire \block_w2_reg_reg[7]_0 ;
  wire \block_w2_reg_reg[8]_0 ;
  wire \block_w2_reg_reg[9]_0 ;
  wire block_w2_we;
  wire \block_w3_reg[0]_i_1_n_0 ;
  wire \block_w3_reg[10]_i_3_n_0 ;
  wire \block_w3_reg[11]_i_2__0_n_0 ;
  wire \block_w3_reg[11]_i_3_n_0 ;
  wire \block_w3_reg[12]_i_3_n_0 ;
  wire \block_w3_reg[13]_i_3_n_0 ;
  wire \block_w3_reg[14]_i_3_n_0 ;
  wire \block_w3_reg[15]_i_3_n_0 ;
  wire \block_w3_reg[16]_i_1_n_0 ;
  wire \block_w3_reg[17]_i_3_n_0 ;
  wire \block_w3_reg[18]_i_2__0_n_0 ;
  wire \block_w3_reg[18]_i_3_n_0 ;
  wire \block_w3_reg[19]_i_3_n_0 ;
  wire \block_w3_reg[1]_i_3_n_0 ;
  wire \block_w3_reg[20]_i_3_n_0 ;
  wire \block_w3_reg[21]_i_3_n_0 ;
  wire \block_w3_reg[22]_i_3_n_0 ;
  wire \block_w3_reg[23]_i_3_n_0 ;
  wire \block_w3_reg[24]_i_3_n_0 ;
  wire \block_w3_reg[25]_i_3_n_0 ;
  wire \block_w3_reg[26]_i_2__0_n_0 ;
  wire \block_w3_reg[26]_i_3_n_0 ;
  wire \block_w3_reg[27]_i_2__0_n_0 ;
  wire \block_w3_reg[27]_i_3_n_0 ;
  wire \block_w3_reg[28]_i_3_n_0 ;
  wire \block_w3_reg[29]_i_3_n_0 ;
  wire \block_w3_reg[2]_i_3_n_0 ;
  wire \block_w3_reg[30]_i_3_n_0 ;
  wire \block_w3_reg[31]_i_3__0_n_0 ;
  wire \block_w3_reg[31]_i_5_n_0 ;
  wire \block_w3_reg[3]_i_3_n_0 ;
  wire \block_w3_reg[4]_i_3_n_0 ;
  wire \block_w3_reg[5]_i_3_n_0 ;
  wire \block_w3_reg[6]_i_3_n_0 ;
  wire \block_w3_reg[7]_i_3_n_0 ;
  wire \block_w3_reg[8]_i_3_n_0 ;
  wire \block_w3_reg[9]_i_3_n_0 ;
  wire \block_w3_reg_reg[0]_0 ;
  wire \block_w3_reg_reg[0]_1 ;
  wire \block_w3_reg_reg[10]_0 ;
  wire \block_w3_reg_reg[10]_i_1_n_0 ;
  wire \block_w3_reg_reg[11]_i_1_n_0 ;
  wire \block_w3_reg_reg[12]_0 ;
  wire \block_w3_reg_reg[12]_i_1_n_0 ;
  wire \block_w3_reg_reg[13]_0 ;
  wire \block_w3_reg_reg[13]_i_1_n_0 ;
  wire \block_w3_reg_reg[14]_0 ;
  wire \block_w3_reg_reg[14]_i_1_n_0 ;
  wire \block_w3_reg_reg[15]_0 ;
  wire \block_w3_reg_reg[15]_i_1_n_0 ;
  wire \block_w3_reg_reg[16]_0 ;
  wire \block_w3_reg_reg[16]_1 ;
  wire \block_w3_reg_reg[17]_0 ;
  wire \block_w3_reg_reg[17]_i_1_n_0 ;
  wire \block_w3_reg_reg[18]_i_1_n_0 ;
  wire \block_w3_reg_reg[19]_0 ;
  wire \block_w3_reg_reg[19]_i_1_n_0 ;
  wire \block_w3_reg_reg[1]_0 ;
  wire \block_w3_reg_reg[1]_i_1_n_0 ;
  wire \block_w3_reg_reg[20]_0 ;
  wire \block_w3_reg_reg[20]_i_1_n_0 ;
  wire \block_w3_reg_reg[21]_0 ;
  wire \block_w3_reg_reg[21]_i_1_n_0 ;
  wire \block_w3_reg_reg[22]_0 ;
  wire \block_w3_reg_reg[22]_i_1_n_0 ;
  wire \block_w3_reg_reg[23]_0 ;
  wire \block_w3_reg_reg[23]_i_1_n_0 ;
  wire \block_w3_reg_reg[24]_0 ;
  wire \block_w3_reg_reg[24]_i_1_n_0 ;
  wire \block_w3_reg_reg[25]_0 ;
  wire \block_w3_reg_reg[25]_i_1_n_0 ;
  wire \block_w3_reg_reg[26]_i_1_n_0 ;
  wire \block_w3_reg_reg[27]_i_1_n_0 ;
  wire \block_w3_reg_reg[28]_0 ;
  wire \block_w3_reg_reg[28]_i_1_n_0 ;
  wire \block_w3_reg_reg[29]_0 ;
  wire \block_w3_reg_reg[29]_i_1_n_0 ;
  wire \block_w3_reg_reg[2]_0 ;
  wire \block_w3_reg_reg[2]_i_1_n_0 ;
  wire \block_w3_reg_reg[30]_0 ;
  wire \block_w3_reg_reg[30]_i_1_n_0 ;
  wire \block_w3_reg_reg[31]_0 ;
  wire \block_w3_reg_reg[31]_i_2_n_0 ;
  wire \block_w3_reg_reg[3]_0 ;
  wire \block_w3_reg_reg[3]_i_1_n_0 ;
  wire \block_w3_reg_reg[4]_0 ;
  wire \block_w3_reg_reg[4]_i_1_n_0 ;
  wire \block_w3_reg_reg[5]_0 ;
  wire \block_w3_reg_reg[5]_i_1_n_0 ;
  wire \block_w3_reg_reg[6]_0 ;
  wire \block_w3_reg_reg[6]_i_1_n_0 ;
  wire \block_w3_reg_reg[7]_0 ;
  wire \block_w3_reg_reg[7]_i_1_n_0 ;
  wire \block_w3_reg_reg[8]_0 ;
  wire \block_w3_reg_reg[8]_i_1_n_0 ;
  wire \block_w3_reg_reg[9]_0 ;
  wire \block_w3_reg_reg[9]_i_1_n_0 ;
  wire block_w3_we;
  wire clk_i;
  wire [1:0]dec_ctrl_new;
  wire [1:1]dec_ctrl_reg;
  wire [127:0]dec_new_block;
  wire dec_ready;
  wire g0_b0__0_n_0;
  wire g0_b0__1_n_0;
  wire g0_b0__2_n_0;
  wire g0_b0_n_0;
  wire g0_b1__0_n_0;
  wire g0_b1__1_n_0;
  wire g0_b1__2_n_0;
  wire g0_b1_n_0;
  wire g0_b2__0_n_0;
  wire g0_b2__1_n_0;
  wire g0_b2__2_n_0;
  wire g0_b2_n_0;
  wire g0_b3__0_n_0;
  wire g0_b3__1_n_0;
  wire g0_b3__2_n_0;
  wire g0_b3_n_0;
  wire g0_b4__0_n_0;
  wire g0_b4__1_n_0;
  wire g0_b4__2_n_0;
  wire g0_b4_n_0;
  wire g0_b5__0_n_0;
  wire g0_b5__1_n_0;
  wire g0_b5__2_n_0;
  wire g0_b5_n_0;
  wire g0_b6__0_n_0;
  wire g0_b6__1_n_0;
  wire g0_b6__2_n_0;
  wire g0_b6_n_0;
  wire g0_b7__0_n_0;
  wire g0_b7__1_n_0;
  wire g0_b7__2_n_0;
  wire g0_b7_n_0;
  wire g1_b0__0_n_0;
  wire g1_b0__1_n_0;
  wire g1_b0__2_n_0;
  wire g1_b0_n_0;
  wire g1_b1__0_n_0;
  wire g1_b1__1_n_0;
  wire g1_b1__2_n_0;
  wire g1_b1_n_0;
  wire g1_b2__0_n_0;
  wire g1_b2__1_n_0;
  wire g1_b2__2_n_0;
  wire g1_b2_n_0;
  wire g1_b3__0_n_0;
  wire g1_b3__1_n_0;
  wire g1_b3__2_n_0;
  wire g1_b3_n_0;
  wire g1_b4__0_n_0;
  wire g1_b4__1_n_0;
  wire g1_b4__2_n_0;
  wire g1_b4_n_0;
  wire g1_b5__0_n_0;
  wire g1_b5__1_n_0;
  wire g1_b5__2_n_0;
  wire g1_b5_n_0;
  wire g1_b6__0_n_0;
  wire g1_b6__1_n_0;
  wire g1_b6__2_n_0;
  wire g1_b6_n_0;
  wire g1_b7__0_n_0;
  wire g1_b7__1_n_0;
  wire g1_b7__2_n_0;
  wire g1_b7_n_0;
  wire g2_b0__0_n_0;
  wire g2_b0__1_n_0;
  wire g2_b0__2_n_0;
  wire g2_b0_n_0;
  wire g2_b1__0_n_0;
  wire g2_b1__1_n_0;
  wire g2_b1__2_n_0;
  wire g2_b1_n_0;
  wire g2_b2__0_n_0;
  wire g2_b2__1_n_0;
  wire g2_b2__2_n_0;
  wire g2_b2_n_0;
  wire g2_b3__0_n_0;
  wire g2_b3__1_n_0;
  wire g2_b3__2_n_0;
  wire g2_b3_n_0;
  wire g2_b4__0_n_0;
  wire g2_b4__1_n_0;
  wire g2_b4__2_n_0;
  wire g2_b4_n_0;
  wire g2_b5__0_n_0;
  wire g2_b5__1_n_0;
  wire g2_b5__2_n_0;
  wire g2_b5_n_0;
  wire g2_b6__0_n_0;
  wire g2_b6__1_n_0;
  wire g2_b6__2_n_0;
  wire g2_b6_n_0;
  wire g2_b7__0_n_0;
  wire g2_b7__1_n_0;
  wire g2_b7__2_n_0;
  wire g2_b7_n_0;
  wire g3_b0__0_n_0;
  wire g3_b0__1_n_0;
  wire g3_b0__2_n_0;
  wire g3_b0_n_0;
  wire g3_b1__0_n_0;
  wire g3_b1__1_n_0;
  wire g3_b1__2_n_0;
  wire g3_b1_n_0;
  wire g3_b2__0_n_0;
  wire g3_b2__1_n_0;
  wire g3_b2__2_n_0;
  wire g3_b2_n_0;
  wire g3_b3__0_n_0;
  wire g3_b3__1_n_0;
  wire g3_b3__2_n_0;
  wire g3_b3_n_0;
  wire g3_b4__0_n_0;
  wire g3_b4__1_n_0;
  wire g3_b4__2_n_0;
  wire g3_b4_n_0;
  wire g3_b5__0_n_0;
  wire g3_b5__1_n_0;
  wire g3_b5__2_n_0;
  wire g3_b5_n_0;
  wire g3_b6__0_n_0;
  wire g3_b6__1_n_0;
  wire g3_b6__2_n_0;
  wire g3_b6_n_0;
  wire g3_b7__0_n_0;
  wire g3_b7__1_n_0;
  wire g3_b7__2_n_0;
  wire g3_b7_n_0;
  wire [6:0]inv_mixcolumns_return0110_out__47;
  wire [6:0]inv_mixcolumns_return0117_out__50;
  wire [7:0]inv_mixcolumns_return0124_out__47;
  wire [6:0]inv_mixcolumns_return0134_out__63;
  wire [7:0]inv_mixcolumns_return0142_out__55;
  wire [6:0]inv_mixcolumns_return0149_out__55;
  wire [7:0]inv_mixcolumns_return0156_out__63;
  wire [6:0]inv_mixcolumns_return0166_out__55;
  wire [7:0]inv_mixcolumns_return0174_out__63;
  wire [6:0]inv_mixcolumns_return0181_out__58;
  wire [7:0]inv_mixcolumns_return0188_out__55;
  wire [6:0]inv_mixcolumns_return0198_out__63;
  wire [6:0]inv_mixcolumns_return0206_out__55;
  wire [6:0]inv_mixcolumns_return0213_out__55;
  wire [7:0]inv_mixcolumns_return0220_out__63;
  wire [6:0]inv_mixcolumns_return0__55;
  wire [2:0]\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11 ;
  wire [31:1]new_sboxw;
  wire [0:0]op126_in;
  wire [0:0]op127_in;
  wire [0:0]op158_in;
  wire [0:0]op159_in;
  wire [0:0]op191_in;
  wire [0:0]op96_in;
  wire [1:0]p_0_in;
  wire [0:0]p_0_in31_in;
  wire [0:0]p_0_in38_in;
  wire [0:0]p_0_in46_in;
  wire [0:0]p_0_in54_in;
  wire [31:0]p_0_in__0;
  wire [75:0]p_0_out;
  wire [2:0]p_1_in;
  wire ready_new;
  wire ready_reg_i_1__0_n_0;
  wire ready_reg_i_2_n_0;
  wire round_ctr_dec__1;
  wire [3:0]round_ctr_new;
  wire round_ctr_set__1;
  wire round_ctr_we;
  wire [15:0]round_key;
  wire rst_i;
  wire [1:0]sword_ctr_new;
  wire sword_ctr_rst;
  wire sword_ctr_we;
  wire [31:0]tmp_sboxw;
  wire [31:0]tmp_sboxw_0;
  wire [1:1]update_type__0;

  LUT6 #(
    .INIT(64'h00000000F4040404)) 
    \FSM_sequential_dec_ctrl_reg[0]_i_1 
       (.I0(p_1_in[1]),
        .I1(p_1_in[0]),
        .I2(dec_ctrl_reg),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(sword_ctr_rst),
        .O(dec_ctrl_new[0]));
  LUT6 #(
    .INIT(64'hFFBAAABAAABAAABA)) 
    \FSM_sequential_dec_ctrl_reg[1]_i_1 
       (.I0(sword_ctr_rst),
        .I1(p_1_in[1]),
        .I2(p_1_in[0]),
        .I3(dec_ctrl_reg),
        .I4(p_0_in[1]),
        .I5(p_0_in[0]),
        .O(\FSM_sequential_dec_ctrl_reg[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT5 #(
    .INIT(32'hB8888888)) 
    \FSM_sequential_dec_ctrl_reg[1]_i_2 
       (.I0(\FSM_sequential_dec_ctrl_reg[1]_i_3_n_0 ),
        .I1(sword_ctr_rst),
        .I2(p_0_in[1]),
        .I3(p_0_in[0]),
        .I4(dec_ctrl_reg),
        .O(dec_ctrl_new[1]));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    \FSM_sequential_dec_ctrl_reg[1]_i_3 
       (.I0(Q[3]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(dec_ctrl_reg),
        .O(\FSM_sequential_dec_ctrl_reg[1]_i_3_n_0 ));
  (* FSM_ENCODED_STATES = "CTRL_INIT:01,CTRL_MAIN:11,CTRL_IDLE:00,CTRL_SBOX:10" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_dec_ctrl_reg_reg[0] 
       (.C(clk_i),
        .CE(\FSM_sequential_dec_ctrl_reg[1]_i_1_n_0 ),
        .CLR(rst_i),
        .D(dec_ctrl_new[0]),
        .Q(sword_ctr_rst));
  (* FSM_ENCODED_STATES = "CTRL_INIT:01,CTRL_MAIN:11,CTRL_IDLE:00,CTRL_SBOX:10" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_dec_ctrl_reg_reg[1] 
       (.C(clk_i),
        .CE(\FSM_sequential_dec_ctrl_reg[1]_i_1_n_0 ),
        .CLR(rst_i),
        .D(dec_ctrl_new[1]),
        .Q(dec_ctrl_reg));
  LUT6 #(
    .INIT(64'hBA10BA1044440000)) 
    \block_w0_reg[0]_i_1 
       (.I0(update_type__0),
        .I1(ready_new),
        .I2(\block_w0_reg_reg[0]_0 ),
        .I3(\block_w0_reg_reg[0]_1 ),
        .I4(p_0_in54_in),
        .I5(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w0_reg[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[10]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[24]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[10]),
        .I5(inv_mixcolumns_return0142_out__55[2]),
        .O(\block_w0_reg[10]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w0_reg[11]_i_2__0 
       (.I0(round_key[12]),
        .I1(dec_new_block[107]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w0_reg[11]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[11]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[25]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[11]),
        .I5(inv_mixcolumns_return0142_out__55[3]),
        .O(\block_w0_reg[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[12]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[26]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[12]),
        .I5(inv_mixcolumns_return0142_out__55[4]),
        .O(\block_w0_reg[12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[13]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[27]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[13]),
        .I5(inv_mixcolumns_return0142_out__55[5]),
        .O(\block_w0_reg[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[14]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[28]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[14]),
        .I5(inv_mixcolumns_return0142_out__55[6]),
        .O(\block_w0_reg[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[15]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[29]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[15]),
        .I5(inv_mixcolumns_return0142_out__55[7]),
        .O(\block_w0_reg[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBA10BA1044440000)) 
    \block_w0_reg[16]_i_1 
       (.I0(update_type__0),
        .I1(ready_new),
        .I2(\block_w0_reg_reg[16]_0 ),
        .I3(\block_w0_reg_reg[16]_1 ),
        .I4(op191_in),
        .I5(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w0_reg[16]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[17]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[15]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[17]),
        .I5(inv_mixcolumns_return0117_out__50[0]),
        .O(\block_w0_reg[17]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w0_reg[18]_i_2__0 
       (.I0(dec_new_block[114]),
        .I1(round_key[13]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w0_reg[18]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[18]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[16]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[18]),
        .I5(inv_mixcolumns_return0117_out__50[1]),
        .O(\block_w0_reg[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[19]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[17]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[19]),
        .I5(inv_mixcolumns_return0117_out__50[2]),
        .O(\block_w0_reg[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[1]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[30]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[1]),
        .I5(inv_mixcolumns_return0166_out__55[0]),
        .O(\block_w0_reg[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[20]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[18]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[20]),
        .I5(inv_mixcolumns_return0117_out__50[3]),
        .O(\block_w0_reg[20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[21]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[19]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[21]),
        .I5(inv_mixcolumns_return0117_out__50[4]),
        .O(\block_w0_reg[21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[22]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[20]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[22]),
        .I5(inv_mixcolumns_return0117_out__50[5]),
        .O(\block_w0_reg[22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[23]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[21]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[23]),
        .I5(inv_mixcolumns_return0117_out__50[6]),
        .O(\block_w0_reg[23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[24]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[68]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[24]),
        .I5(inv_mixcolumns_return0220_out__63[0]),
        .O(\block_w0_reg[24]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[25]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[69]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[25]),
        .I5(inv_mixcolumns_return0220_out__63[1]),
        .O(\block_w0_reg[25]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w0_reg[26]_i_2__0 
       (.I0(dec_new_block[122]),
        .I1(round_key[14]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w0_reg[26]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[26]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[70]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[26]),
        .I5(inv_mixcolumns_return0220_out__63[2]),
        .O(\block_w0_reg[26]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w0_reg[27]_i_2__0 
       (.I0(dec_new_block[123]),
        .I1(round_key[15]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w0_reg[27]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[27]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[71]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[27]),
        .I5(inv_mixcolumns_return0220_out__63[3]),
        .O(\block_w0_reg[27]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[28]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[72]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[28]),
        .I5(inv_mixcolumns_return0220_out__63[4]),
        .O(\block_w0_reg[28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[29]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[73]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[29]),
        .I5(inv_mixcolumns_return0220_out__63[5]),
        .O(\block_w0_reg[29]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[2]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[31]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[2]),
        .I5(inv_mixcolumns_return0166_out__55[1]),
        .O(\block_w0_reg[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[30]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[74]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[30]),
        .I5(inv_mixcolumns_return0220_out__63[6]),
        .O(\block_w0_reg[30]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h46464656)) 
    \block_w0_reg[31]_i_1 
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(p_0_in[0]),
        .I4(p_0_in[1]),
        .O(block_w0_we));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[31]_i_4 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[75]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[31]),
        .I5(inv_mixcolumns_return0220_out__63[7]),
        .O(\block_w0_reg[31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[3]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[32]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[3]),
        .I5(inv_mixcolumns_return0166_out__55[2]),
        .O(\block_w0_reg[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[4]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[33]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[4]),
        .I5(inv_mixcolumns_return0166_out__55[3]),
        .O(\block_w0_reg[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[5]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[34]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[5]),
        .I5(inv_mixcolumns_return0166_out__55[4]),
        .O(\block_w0_reg[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[6]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[35]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[6]),
        .I5(inv_mixcolumns_return0166_out__55[5]),
        .O(\block_w0_reg[6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[7]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[36]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[7]),
        .I5(inv_mixcolumns_return0166_out__55[6]),
        .O(\block_w0_reg[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[8]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[22]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[8]),
        .I5(inv_mixcolumns_return0142_out__55[0]),
        .O(\block_w0_reg[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w0_reg[9]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[23]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11 [1]),
        .I5(inv_mixcolumns_return0142_out__55[1]),
        .O(\block_w0_reg[9]_i_3_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[0] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[0]_i_1_n_0 ),
        .Q(dec_new_block[96]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[10] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[10]_i_1_n_0 ),
        .Q(dec_new_block[106]));
  MUXF7 \block_w0_reg_reg[10]_i_1 
       (.I0(\block_w0_reg_reg[10]_0 ),
        .I1(\block_w0_reg[10]_i_3_n_0 ),
        .O(\block_w0_reg_reg[10]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[11] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[11]_i_1_n_0 ),
        .Q(dec_new_block[107]));
  MUXF7 \block_w0_reg_reg[11]_i_1 
       (.I0(\block_w0_reg[11]_i_2__0_n_0 ),
        .I1(\block_w0_reg[11]_i_3_n_0 ),
        .O(\block_w0_reg_reg[11]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[12] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[12]_i_1_n_0 ),
        .Q(dec_new_block[108]));
  MUXF7 \block_w0_reg_reg[12]_i_1 
       (.I0(\block_w0_reg_reg[12]_0 ),
        .I1(\block_w0_reg[12]_i_3_n_0 ),
        .O(\block_w0_reg_reg[12]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[13] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[13]_i_1_n_0 ),
        .Q(dec_new_block[109]));
  MUXF7 \block_w0_reg_reg[13]_i_1 
       (.I0(\block_w0_reg_reg[13]_0 ),
        .I1(\block_w0_reg[13]_i_3_n_0 ),
        .O(\block_w0_reg_reg[13]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[14] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[14]_i_1_n_0 ),
        .Q(dec_new_block[110]));
  MUXF7 \block_w0_reg_reg[14]_i_1 
       (.I0(\block_w0_reg_reg[14]_0 ),
        .I1(\block_w0_reg[14]_i_3_n_0 ),
        .O(\block_w0_reg_reg[14]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[15] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[15]_i_1_n_0 ),
        .Q(dec_new_block[111]));
  MUXF7 \block_w0_reg_reg[15]_i_1 
       (.I0(\block_w0_reg_reg[15]_0 ),
        .I1(\block_w0_reg[15]_i_3_n_0 ),
        .O(\block_w0_reg_reg[15]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[16] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[16]_i_1_n_0 ),
        .Q(dec_new_block[112]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[17] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[17]_i_1_n_0 ),
        .Q(dec_new_block[113]));
  MUXF7 \block_w0_reg_reg[17]_i_1 
       (.I0(\block_w0_reg_reg[17]_0 ),
        .I1(\block_w0_reg[17]_i_3_n_0 ),
        .O(\block_w0_reg_reg[17]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[18] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[18]_i_1_n_0 ),
        .Q(dec_new_block[114]));
  MUXF7 \block_w0_reg_reg[18]_i_1 
       (.I0(\block_w0_reg[18]_i_2__0_n_0 ),
        .I1(\block_w0_reg[18]_i_3_n_0 ),
        .O(\block_w0_reg_reg[18]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[19] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[19]_i_1_n_0 ),
        .Q(dec_new_block[115]));
  MUXF7 \block_w0_reg_reg[19]_i_1 
       (.I0(\block_w0_reg_reg[19]_0 ),
        .I1(\block_w0_reg[19]_i_3_n_0 ),
        .O(\block_w0_reg_reg[19]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[1] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[1]_i_1_n_0 ),
        .Q(dec_new_block[97]));
  MUXF7 \block_w0_reg_reg[1]_i_1 
       (.I0(\block_w0_reg_reg[1]_0 ),
        .I1(\block_w0_reg[1]_i_3_n_0 ),
        .O(\block_w0_reg_reg[1]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[20] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[20]_i_1_n_0 ),
        .Q(dec_new_block[116]));
  MUXF7 \block_w0_reg_reg[20]_i_1 
       (.I0(\block_w0_reg_reg[20]_0 ),
        .I1(\block_w0_reg[20]_i_3_n_0 ),
        .O(\block_w0_reg_reg[20]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[21] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[21]_i_1_n_0 ),
        .Q(dec_new_block[117]));
  MUXF7 \block_w0_reg_reg[21]_i_1 
       (.I0(\block_w0_reg_reg[21]_0 ),
        .I1(\block_w0_reg[21]_i_3_n_0 ),
        .O(\block_w0_reg_reg[21]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[22] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[22]_i_1_n_0 ),
        .Q(dec_new_block[118]));
  MUXF7 \block_w0_reg_reg[22]_i_1 
       (.I0(\block_w0_reg_reg[22]_0 ),
        .I1(\block_w0_reg[22]_i_3_n_0 ),
        .O(\block_w0_reg_reg[22]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[23] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[23]_i_1_n_0 ),
        .Q(dec_new_block[119]));
  MUXF7 \block_w0_reg_reg[23]_i_1 
       (.I0(\block_w0_reg_reg[23]_0 ),
        .I1(\block_w0_reg[23]_i_3_n_0 ),
        .O(\block_w0_reg_reg[23]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[24] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[24]_i_1_n_0 ),
        .Q(dec_new_block[120]));
  MUXF7 \block_w0_reg_reg[24]_i_1 
       (.I0(\block_w0_reg_reg[24]_0 ),
        .I1(\block_w0_reg[24]_i_3_n_0 ),
        .O(\block_w0_reg_reg[24]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[25] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[25]_i_1_n_0 ),
        .Q(dec_new_block[121]));
  MUXF7 \block_w0_reg_reg[25]_i_1 
       (.I0(\block_w0_reg_reg[25]_0 ),
        .I1(\block_w0_reg[25]_i_3_n_0 ),
        .O(\block_w0_reg_reg[25]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[26] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[26]_i_1_n_0 ),
        .Q(dec_new_block[122]));
  MUXF7 \block_w0_reg_reg[26]_i_1 
       (.I0(\block_w0_reg[26]_i_2__0_n_0 ),
        .I1(\block_w0_reg[26]_i_3_n_0 ),
        .O(\block_w0_reg_reg[26]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[27] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[27]_i_1_n_0 ),
        .Q(dec_new_block[123]));
  MUXF7 \block_w0_reg_reg[27]_i_1 
       (.I0(\block_w0_reg[27]_i_2__0_n_0 ),
        .I1(\block_w0_reg[27]_i_3_n_0 ),
        .O(\block_w0_reg_reg[27]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[28] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[28]_i_1_n_0 ),
        .Q(dec_new_block[124]));
  MUXF7 \block_w0_reg_reg[28]_i_1 
       (.I0(\block_w0_reg_reg[28]_0 ),
        .I1(\block_w0_reg[28]_i_3_n_0 ),
        .O(\block_w0_reg_reg[28]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[29] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[29]_i_1_n_0 ),
        .Q(dec_new_block[125]));
  MUXF7 \block_w0_reg_reg[29]_i_1 
       (.I0(\block_w0_reg_reg[29]_0 ),
        .I1(\block_w0_reg[29]_i_3_n_0 ),
        .O(\block_w0_reg_reg[29]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[2] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[2]_i_1_n_0 ),
        .Q(dec_new_block[98]));
  MUXF7 \block_w0_reg_reg[2]_i_1 
       (.I0(\block_w0_reg_reg[2]_0 ),
        .I1(\block_w0_reg[2]_i_3_n_0 ),
        .O(\block_w0_reg_reg[2]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[30] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[30]_i_1_n_0 ),
        .Q(dec_new_block[126]));
  MUXF7 \block_w0_reg_reg[30]_i_1 
       (.I0(\block_w0_reg_reg[30]_0 ),
        .I1(\block_w0_reg[30]_i_3_n_0 ),
        .O(\block_w0_reg_reg[30]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[31] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[31]_i_2_n_0 ),
        .Q(dec_new_block[127]));
  MUXF7 \block_w0_reg_reg[31]_i_2 
       (.I0(\block_w0_reg_reg[31]_0 ),
        .I1(\block_w0_reg[31]_i_4_n_0 ),
        .O(\block_w0_reg_reg[31]_i_2_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[3] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[3]_i_1_n_0 ),
        .Q(dec_new_block[99]));
  MUXF7 \block_w0_reg_reg[3]_i_1 
       (.I0(\block_w0_reg_reg[3]_0 ),
        .I1(\block_w0_reg[3]_i_3_n_0 ),
        .O(\block_w0_reg_reg[3]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[4] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[4]_i_1_n_0 ),
        .Q(dec_new_block[100]));
  MUXF7 \block_w0_reg_reg[4]_i_1 
       (.I0(\block_w0_reg_reg[4]_0 ),
        .I1(\block_w0_reg[4]_i_3_n_0 ),
        .O(\block_w0_reg_reg[4]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[5] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[5]_i_1_n_0 ),
        .Q(dec_new_block[101]));
  MUXF7 \block_w0_reg_reg[5]_i_1 
       (.I0(\block_w0_reg_reg[5]_0 ),
        .I1(\block_w0_reg[5]_i_3_n_0 ),
        .O(\block_w0_reg_reg[5]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[6] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[6]_i_1_n_0 ),
        .Q(dec_new_block[102]));
  MUXF7 \block_w0_reg_reg[6]_i_1 
       (.I0(\block_w0_reg_reg[6]_0 ),
        .I1(\block_w0_reg[6]_i_3_n_0 ),
        .O(\block_w0_reg_reg[6]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[7] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[7]_i_1_n_0 ),
        .Q(dec_new_block[103]));
  MUXF7 \block_w0_reg_reg[7]_i_1 
       (.I0(\block_w0_reg_reg[7]_0 ),
        .I1(\block_w0_reg[7]_i_3_n_0 ),
        .O(\block_w0_reg_reg[7]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[8] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[8]_i_1_n_0 ),
        .Q(dec_new_block[104]));
  MUXF7 \block_w0_reg_reg[8]_i_1 
       (.I0(\block_w0_reg_reg[8]_0 ),
        .I1(\block_w0_reg[8]_i_3_n_0 ),
        .O(\block_w0_reg_reg[8]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[9] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg_reg[9]_i_1_n_0 ),
        .Q(dec_new_block[105]));
  MUXF7 \block_w0_reg_reg[9]_i_1 
       (.I0(\block_w0_reg_reg[9]_0 ),
        .I1(\block_w0_reg[9]_i_3_n_0 ),
        .O(\block_w0_reg_reg[9]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hBA10BA1044440000)) 
    \block_w1_reg[0]_i_1 
       (.I0(update_type__0),
        .I1(ready_new),
        .I2(\block_w1_reg_reg[0]_0 ),
        .I3(\block_w1_reg_reg[0]_1 ),
        .I4(p_0_in46_in),
        .I5(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w1_reg[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[10]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[9]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[10]),
        .I5(inv_mixcolumns_return0110_out__47[1]),
        .O(\block_w1_reg[10]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w1_reg[11]_i_2__0 
       (.I0(round_key[8]),
        .I1(dec_new_block[75]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w1_reg[11]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[11]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[10]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[11]),
        .I5(inv_mixcolumns_return0110_out__47[2]),
        .O(\block_w1_reg[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[12]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[11]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[12]),
        .I5(inv_mixcolumns_return0110_out__47[3]),
        .O(\block_w1_reg[12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[13]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[12]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[13]),
        .I5(inv_mixcolumns_return0110_out__47[4]),
        .O(\block_w1_reg[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[14]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[13]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[14]),
        .I5(inv_mixcolumns_return0110_out__47[5]),
        .O(\block_w1_reg[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[15]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[14]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[15]),
        .I5(inv_mixcolumns_return0110_out__47[6]),
        .O(\block_w1_reg[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBA10BA1044440000)) 
    \block_w1_reg[16]_i_1 
       (.I0(update_type__0),
        .I1(ready_new),
        .I2(\block_w1_reg_reg[16]_0 ),
        .I3(\block_w1_reg_reg[16]_1 ),
        .I4(op159_in),
        .I5(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w1_reg[16]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[17]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[61]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[17]),
        .I5(inv_mixcolumns_return0213_out__55[0]),
        .O(\block_w1_reg[17]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w1_reg[18]_i_2__0 
       (.I0(dec_new_block[82]),
        .I1(round_key[9]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w1_reg[18]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[18]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[62]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[18]),
        .I5(inv_mixcolumns_return0213_out__55[1]),
        .O(\block_w1_reg[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[19]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[63]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[19]),
        .I5(inv_mixcolumns_return0213_out__55[2]),
        .O(\block_w1_reg[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[1]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[8]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[1]),
        .I5(inv_mixcolumns_return0134_out__63[0]),
        .O(\block_w1_reg[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[20]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[64]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[20]),
        .I5(inv_mixcolumns_return0213_out__55[3]),
        .O(\block_w1_reg[20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[21]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[65]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[21]),
        .I5(inv_mixcolumns_return0213_out__55[4]),
        .O(\block_w1_reg[21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[22]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[66]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[22]),
        .I5(inv_mixcolumns_return0213_out__55[5]),
        .O(\block_w1_reg[22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[23]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[67]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[23]),
        .I5(inv_mixcolumns_return0213_out__55[6]),
        .O(\block_w1_reg[23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[24]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[38]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[24]),
        .I5(inv_mixcolumns_return0188_out__55[0]),
        .O(\block_w1_reg[24]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[25]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[39]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[25]),
        .I5(inv_mixcolumns_return0188_out__55[1]),
        .O(\block_w1_reg[25]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w1_reg[26]_i_2__0 
       (.I0(dec_new_block[90]),
        .I1(round_key[10]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w1_reg[26]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[26]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[40]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[26]),
        .I5(inv_mixcolumns_return0188_out__55[2]),
        .O(\block_w1_reg[26]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w1_reg[27]_i_2__0 
       (.I0(dec_new_block[91]),
        .I1(round_key[11]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w1_reg[27]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[27]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[41]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[27]),
        .I5(inv_mixcolumns_return0188_out__55[3]),
        .O(\block_w1_reg[27]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[28]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[42]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[28]),
        .I5(inv_mixcolumns_return0188_out__55[4]),
        .O(\block_w1_reg[28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[29]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[43]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[29]),
        .I5(inv_mixcolumns_return0188_out__55[5]),
        .O(\block_w1_reg[29]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[2]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[9]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[2]),
        .I5(inv_mixcolumns_return0134_out__63[1]),
        .O(\block_w1_reg[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[30]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[44]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[30]),
        .I5(inv_mixcolumns_return0188_out__55[6]),
        .O(\block_w1_reg[30]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h45446666)) 
    \block_w1_reg[31]_i_1 
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(p_0_in[1]),
        .I3(p_0_in[0]),
        .I4(update_type__0),
        .O(block_w1_we));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[31]_i_4 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[45]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[31]),
        .I5(inv_mixcolumns_return0188_out__55[7]),
        .O(\block_w1_reg[31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[3]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[10]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[3]),
        .I5(inv_mixcolumns_return0134_out__63[2]),
        .O(\block_w1_reg[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[4]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[11]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[4]),
        .I5(inv_mixcolumns_return0134_out__63[3]),
        .O(\block_w1_reg[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[5]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[12]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[5]),
        .I5(inv_mixcolumns_return0134_out__63[4]),
        .O(\block_w1_reg[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[6]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[13]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[6]),
        .I5(inv_mixcolumns_return0134_out__63[5]),
        .O(\block_w1_reg[6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[7]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[14]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[7]),
        .I5(inv_mixcolumns_return0134_out__63[6]),
        .O(\block_w1_reg[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w1_reg[8]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[7]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[8]),
        .I5(inv_mixcolumns_return0110_out__47[0]),
        .O(\block_w1_reg[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBA10BA1044440000)) 
    \block_w1_reg[9]_i_1 
       (.I0(update_type__0),
        .I1(ready_new),
        .I2(\block_w1_reg[9]_i_2__0_n_0 ),
        .I3(\block_w1_reg_reg[9]_0 ),
        .I4(op158_in),
        .I5(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w1_reg[9]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \block_w1_reg[9]_i_2__0 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I1(addroundkey_return[8]),
        .O(\block_w1_reg[9]_i_2__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[0] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[0]_i_1_n_0 ),
        .Q(dec_new_block[64]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[10] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[10]_i_1_n_0 ),
        .Q(dec_new_block[74]));
  MUXF7 \block_w1_reg_reg[10]_i_1 
       (.I0(\block_w1_reg_reg[10]_0 ),
        .I1(\block_w1_reg[10]_i_3_n_0 ),
        .O(\block_w1_reg_reg[10]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[11] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[11]_i_1_n_0 ),
        .Q(dec_new_block[75]));
  MUXF7 \block_w1_reg_reg[11]_i_1 
       (.I0(\block_w1_reg[11]_i_2__0_n_0 ),
        .I1(\block_w1_reg[11]_i_3_n_0 ),
        .O(\block_w1_reg_reg[11]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[12] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[12]_i_1_n_0 ),
        .Q(dec_new_block[76]));
  MUXF7 \block_w1_reg_reg[12]_i_1 
       (.I0(\block_w1_reg_reg[12]_0 ),
        .I1(\block_w1_reg[12]_i_3_n_0 ),
        .O(\block_w1_reg_reg[12]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[13] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[13]_i_1_n_0 ),
        .Q(dec_new_block[77]));
  MUXF7 \block_w1_reg_reg[13]_i_1 
       (.I0(\block_w1_reg_reg[13]_0 ),
        .I1(\block_w1_reg[13]_i_3_n_0 ),
        .O(\block_w1_reg_reg[13]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[14] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[14]_i_1_n_0 ),
        .Q(dec_new_block[78]));
  MUXF7 \block_w1_reg_reg[14]_i_1 
       (.I0(\block_w1_reg_reg[14]_0 ),
        .I1(\block_w1_reg[14]_i_3_n_0 ),
        .O(\block_w1_reg_reg[14]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[15] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[15]_i_1_n_0 ),
        .Q(dec_new_block[79]));
  MUXF7 \block_w1_reg_reg[15]_i_1 
       (.I0(\block_w1_reg_reg[15]_0 ),
        .I1(\block_w1_reg[15]_i_3_n_0 ),
        .O(\block_w1_reg_reg[15]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[16] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[16]_i_1_n_0 ),
        .Q(dec_new_block[80]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[17] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[17]_i_1_n_0 ),
        .Q(dec_new_block[81]));
  MUXF7 \block_w1_reg_reg[17]_i_1 
       (.I0(\block_w1_reg_reg[17]_0 ),
        .I1(\block_w1_reg[17]_i_3_n_0 ),
        .O(\block_w1_reg_reg[17]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[18] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[18]_i_1_n_0 ),
        .Q(dec_new_block[82]));
  MUXF7 \block_w1_reg_reg[18]_i_1 
       (.I0(\block_w1_reg[18]_i_2__0_n_0 ),
        .I1(\block_w1_reg[18]_i_3_n_0 ),
        .O(\block_w1_reg_reg[18]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[19] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[19]_i_1_n_0 ),
        .Q(dec_new_block[83]));
  MUXF7 \block_w1_reg_reg[19]_i_1 
       (.I0(\block_w1_reg_reg[19]_0 ),
        .I1(\block_w1_reg[19]_i_3_n_0 ),
        .O(\block_w1_reg_reg[19]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[1] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[1]_i_1_n_0 ),
        .Q(dec_new_block[65]));
  MUXF7 \block_w1_reg_reg[1]_i_1 
       (.I0(\block_w1_reg_reg[1]_0 ),
        .I1(\block_w1_reg[1]_i_3_n_0 ),
        .O(\block_w1_reg_reg[1]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[20] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[20]_i_1_n_0 ),
        .Q(dec_new_block[84]));
  MUXF7 \block_w1_reg_reg[20]_i_1 
       (.I0(\block_w1_reg_reg[20]_0 ),
        .I1(\block_w1_reg[20]_i_3_n_0 ),
        .O(\block_w1_reg_reg[20]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[21] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[21]_i_1_n_0 ),
        .Q(dec_new_block[85]));
  MUXF7 \block_w1_reg_reg[21]_i_1 
       (.I0(\block_w1_reg_reg[21]_0 ),
        .I1(\block_w1_reg[21]_i_3_n_0 ),
        .O(\block_w1_reg_reg[21]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[22] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[22]_i_1_n_0 ),
        .Q(dec_new_block[86]));
  MUXF7 \block_w1_reg_reg[22]_i_1 
       (.I0(\block_w1_reg_reg[22]_0 ),
        .I1(\block_w1_reg[22]_i_3_n_0 ),
        .O(\block_w1_reg_reg[22]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[23] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[23]_i_1_n_0 ),
        .Q(dec_new_block[87]));
  MUXF7 \block_w1_reg_reg[23]_i_1 
       (.I0(\block_w1_reg_reg[23]_0 ),
        .I1(\block_w1_reg[23]_i_3_n_0 ),
        .O(\block_w1_reg_reg[23]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[24] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[24]_i_1_n_0 ),
        .Q(dec_new_block[88]));
  MUXF7 \block_w1_reg_reg[24]_i_1 
       (.I0(\block_w1_reg_reg[24]_0 ),
        .I1(\block_w1_reg[24]_i_3_n_0 ),
        .O(\block_w1_reg_reg[24]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[25] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[25]_i_1_n_0 ),
        .Q(dec_new_block[89]));
  MUXF7 \block_w1_reg_reg[25]_i_1 
       (.I0(\block_w1_reg_reg[25]_0 ),
        .I1(\block_w1_reg[25]_i_3_n_0 ),
        .O(\block_w1_reg_reg[25]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[26] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[26]_i_1_n_0 ),
        .Q(dec_new_block[90]));
  MUXF7 \block_w1_reg_reg[26]_i_1 
       (.I0(\block_w1_reg[26]_i_2__0_n_0 ),
        .I1(\block_w1_reg[26]_i_3_n_0 ),
        .O(\block_w1_reg_reg[26]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[27] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[27]_i_1_n_0 ),
        .Q(dec_new_block[91]));
  MUXF7 \block_w1_reg_reg[27]_i_1 
       (.I0(\block_w1_reg[27]_i_2__0_n_0 ),
        .I1(\block_w1_reg[27]_i_3_n_0 ),
        .O(\block_w1_reg_reg[27]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[28] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[28]_i_1_n_0 ),
        .Q(dec_new_block[92]));
  MUXF7 \block_w1_reg_reg[28]_i_1 
       (.I0(\block_w1_reg_reg[28]_0 ),
        .I1(\block_w1_reg[28]_i_3_n_0 ),
        .O(\block_w1_reg_reg[28]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[29] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[29]_i_1_n_0 ),
        .Q(dec_new_block[93]));
  MUXF7 \block_w1_reg_reg[29]_i_1 
       (.I0(\block_w1_reg_reg[29]_0 ),
        .I1(\block_w1_reg[29]_i_3_n_0 ),
        .O(\block_w1_reg_reg[29]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[2] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[2]_i_1_n_0 ),
        .Q(dec_new_block[66]));
  MUXF7 \block_w1_reg_reg[2]_i_1 
       (.I0(\block_w1_reg_reg[2]_0 ),
        .I1(\block_w1_reg[2]_i_3_n_0 ),
        .O(\block_w1_reg_reg[2]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[30] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[30]_i_1_n_0 ),
        .Q(dec_new_block[94]));
  MUXF7 \block_w1_reg_reg[30]_i_1 
       (.I0(\block_w1_reg_reg[30]_0 ),
        .I1(\block_w1_reg[30]_i_3_n_0 ),
        .O(\block_w1_reg_reg[30]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[31] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[31]_i_2_n_0 ),
        .Q(dec_new_block[95]));
  MUXF7 \block_w1_reg_reg[31]_i_2 
       (.I0(\block_w1_reg_reg[31]_0 ),
        .I1(\block_w1_reg[31]_i_4_n_0 ),
        .O(\block_w1_reg_reg[31]_i_2_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[3] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[3]_i_1_n_0 ),
        .Q(dec_new_block[67]));
  MUXF7 \block_w1_reg_reg[3]_i_1 
       (.I0(\block_w1_reg_reg[3]_0 ),
        .I1(\block_w1_reg[3]_i_3_n_0 ),
        .O(\block_w1_reg_reg[3]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[4] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[4]_i_1_n_0 ),
        .Q(dec_new_block[68]));
  MUXF7 \block_w1_reg_reg[4]_i_1 
       (.I0(\block_w1_reg_reg[4]_0 ),
        .I1(\block_w1_reg[4]_i_3_n_0 ),
        .O(\block_w1_reg_reg[4]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[5] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[5]_i_1_n_0 ),
        .Q(dec_new_block[69]));
  MUXF7 \block_w1_reg_reg[5]_i_1 
       (.I0(\block_w1_reg_reg[5]_0 ),
        .I1(\block_w1_reg[5]_i_3_n_0 ),
        .O(\block_w1_reg_reg[5]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[6] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[6]_i_1_n_0 ),
        .Q(dec_new_block[70]));
  MUXF7 \block_w1_reg_reg[6]_i_1 
       (.I0(\block_w1_reg_reg[6]_0 ),
        .I1(\block_w1_reg[6]_i_3_n_0 ),
        .O(\block_w1_reg_reg[6]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[7] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[7]_i_1_n_0 ),
        .Q(dec_new_block[71]));
  MUXF7 \block_w1_reg_reg[7]_i_1 
       (.I0(\block_w1_reg_reg[7]_0 ),
        .I1(\block_w1_reg[7]_i_3_n_0 ),
        .O(\block_w1_reg_reg[7]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[8] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg_reg[8]_i_1_n_0 ),
        .Q(dec_new_block[72]));
  MUXF7 \block_w1_reg_reg[8]_i_1 
       (.I0(\block_w1_reg_reg[8]_0 ),
        .I1(\block_w1_reg[8]_i_3_n_0 ),
        .O(\block_w1_reg_reg[8]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[9] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[9]_i_1_n_0 ),
        .Q(dec_new_block[73]));
  LUT6 #(
    .INIT(64'hBA10BA1044440000)) 
    \block_w2_reg[0]_i_1 
       (.I0(update_type__0),
        .I1(ready_new),
        .I2(\block_w2_reg_reg[0]_0 ),
        .I3(\block_w2_reg_reg[0]_1 ),
        .I4(p_0_in38_in),
        .I5(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(p_0_in__0[0]));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[10]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[55]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[10]),
        .I5(inv_mixcolumns_return0206_out__55[1]),
        .O(\block_w2_reg[10]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w2_reg[11]_i_2__0 
       (.I0(round_key[4]),
        .I1(dec_new_block[43]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w2_reg[11]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[11]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[56]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[11]),
        .I5(inv_mixcolumns_return0206_out__55[2]),
        .O(\block_w2_reg[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[12]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[57]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[12]),
        .I5(inv_mixcolumns_return0206_out__55[3]),
        .O(\block_w2_reg[12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[13]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[58]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[13]),
        .I5(inv_mixcolumns_return0206_out__55[4]),
        .O(\block_w2_reg[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[14]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[59]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[14]),
        .I5(inv_mixcolumns_return0206_out__55[5]),
        .O(\block_w2_reg[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[15]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[60]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[15]),
        .I5(inv_mixcolumns_return0206_out__55[6]),
        .O(\block_w2_reg[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBA10BA1044440000)) 
    \block_w2_reg[16]_i_1 
       (.I0(update_type__0),
        .I1(ready_new),
        .I2(\block_w2_reg_reg[16]_0 ),
        .I3(\block_w2_reg_reg[16]_1 ),
        .I4(op127_in),
        .I5(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(p_0_in__0[16]));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[17]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[37]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[17]),
        .I5(inv_mixcolumns_return0181_out__58[0]),
        .O(\block_w2_reg[17]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w2_reg[18]_i_2__0 
       (.I0(dec_new_block[50]),
        .I1(round_key[5]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w2_reg[18]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[18]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[38]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[18]),
        .I5(inv_mixcolumns_return0181_out__58[1]),
        .O(\block_w2_reg[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[19]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[39]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[19]),
        .I5(inv_mixcolumns_return0181_out__58[2]),
        .O(\block_w2_reg[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[1]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[0]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[1]),
        .I5(inv_mixcolumns_return0__55[0]),
        .O(\block_w2_reg[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[20]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[40]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[20]),
        .I5(inv_mixcolumns_return0181_out__58[3]),
        .O(\block_w2_reg[20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[21]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[41]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[21]),
        .I5(inv_mixcolumns_return0181_out__58[4]),
        .O(\block_w2_reg[21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[22]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[42]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[22]),
        .I5(inv_mixcolumns_return0181_out__58[5]),
        .O(\block_w2_reg[22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[23]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[43]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[23]),
        .I5(inv_mixcolumns_return0181_out__58[6]),
        .O(\block_w2_reg[23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[24]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[22]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[24]),
        .I5(inv_mixcolumns_return0156_out__63[0]),
        .O(\block_w2_reg[24]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[25]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[23]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[25]),
        .I5(inv_mixcolumns_return0156_out__63[1]),
        .O(\block_w2_reg[25]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w2_reg[26]_i_2__0 
       (.I0(dec_new_block[58]),
        .I1(round_key[6]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w2_reg[26]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[26]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[24]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[26]),
        .I5(inv_mixcolumns_return0156_out__63[2]),
        .O(\block_w2_reg[26]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w2_reg[27]_i_2__0 
       (.I0(dec_new_block[59]),
        .I1(round_key[7]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w2_reg[27]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[27]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[25]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[27]),
        .I5(inv_mixcolumns_return0156_out__63[3]),
        .O(\block_w2_reg[27]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[28]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[26]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[28]),
        .I5(inv_mixcolumns_return0156_out__63[4]),
        .O(\block_w2_reg[28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[29]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[27]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[29]),
        .I5(inv_mixcolumns_return0156_out__63[5]),
        .O(\block_w2_reg[29]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[2]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[1]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[2]),
        .I5(inv_mixcolumns_return0__55[1]),
        .O(\block_w2_reg[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[30]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[28]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[30]),
        .I5(inv_mixcolumns_return0156_out__63[6]),
        .O(\block_w2_reg[30]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h45664466)) 
    \block_w2_reg[31]_i_1 
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(p_0_in[0]),
        .I3(update_type__0),
        .I4(p_0_in[1]),
        .O(block_w2_we));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[31]_i_4 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[29]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[31]),
        .I5(inv_mixcolumns_return0156_out__63[7]),
        .O(\block_w2_reg[31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[3]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[2]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[3]),
        .I5(inv_mixcolumns_return0__55[2]),
        .O(\block_w2_reg[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[4]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[3]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[4]),
        .I5(inv_mixcolumns_return0__55[3]),
        .O(\block_w2_reg[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[5]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[4]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[5]),
        .I5(inv_mixcolumns_return0__55[4]),
        .O(\block_w2_reg[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[6]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[5]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[6]),
        .I5(inv_mixcolumns_return0__55[5]),
        .O(\block_w2_reg[6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[7]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(addroundkey_return[6]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[7]),
        .I5(inv_mixcolumns_return0__55[6]),
        .O(\block_w2_reg[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w2_reg[8]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[53]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[8]),
        .I5(inv_mixcolumns_return0206_out__55[0]),
        .O(\block_w2_reg[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBA10BA1044440000)) 
    \block_w2_reg[9]_i_1 
       (.I0(update_type__0),
        .I1(ready_new),
        .I2(\block_w2_reg[9]_i_2_n_0 ),
        .I3(\block_w2_reg_reg[9]_0 ),
        .I4(op126_in),
        .I5(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(p_0_in__0[9]));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \block_w2_reg[9]_i_2 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I1(p_0_out[54]),
        .O(\block_w2_reg[9]_i_2_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[0] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[0]),
        .Q(dec_new_block[32]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[10] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[10]),
        .Q(dec_new_block[42]));
  MUXF7 \block_w2_reg_reg[10]_i_1 
       (.I0(\block_w2_reg_reg[10]_0 ),
        .I1(\block_w2_reg[10]_i_3_n_0 ),
        .O(p_0_in__0[10]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[11] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[11]),
        .Q(dec_new_block[43]));
  MUXF7 \block_w2_reg_reg[11]_i_1 
       (.I0(\block_w2_reg[11]_i_2__0_n_0 ),
        .I1(\block_w2_reg[11]_i_3_n_0 ),
        .O(p_0_in__0[11]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[12] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[12]),
        .Q(dec_new_block[44]));
  MUXF7 \block_w2_reg_reg[12]_i_1 
       (.I0(\block_w2_reg_reg[12]_0 ),
        .I1(\block_w2_reg[12]_i_3_n_0 ),
        .O(p_0_in__0[12]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[13] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[13]),
        .Q(dec_new_block[45]));
  MUXF7 \block_w2_reg_reg[13]_i_1 
       (.I0(\block_w2_reg_reg[13]_0 ),
        .I1(\block_w2_reg[13]_i_3_n_0 ),
        .O(p_0_in__0[13]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[14] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[14]),
        .Q(dec_new_block[46]));
  MUXF7 \block_w2_reg_reg[14]_i_1 
       (.I0(\block_w2_reg_reg[14]_0 ),
        .I1(\block_w2_reg[14]_i_3_n_0 ),
        .O(p_0_in__0[14]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[15] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[15]),
        .Q(dec_new_block[47]));
  MUXF7 \block_w2_reg_reg[15]_i_1 
       (.I0(\block_w2_reg_reg[15]_0 ),
        .I1(\block_w2_reg[15]_i_3_n_0 ),
        .O(p_0_in__0[15]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[16] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[16]),
        .Q(dec_new_block[48]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[17] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[17]),
        .Q(dec_new_block[49]));
  MUXF7 \block_w2_reg_reg[17]_i_1 
       (.I0(\block_w2_reg_reg[17]_0 ),
        .I1(\block_w2_reg[17]_i_3_n_0 ),
        .O(p_0_in__0[17]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[18] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[18]),
        .Q(dec_new_block[50]));
  MUXF7 \block_w2_reg_reg[18]_i_1 
       (.I0(\block_w2_reg[18]_i_2__0_n_0 ),
        .I1(\block_w2_reg[18]_i_3_n_0 ),
        .O(p_0_in__0[18]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[19] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[19]),
        .Q(dec_new_block[51]));
  MUXF7 \block_w2_reg_reg[19]_i_1 
       (.I0(\block_w2_reg_reg[19]_0 ),
        .I1(\block_w2_reg[19]_i_3_n_0 ),
        .O(p_0_in__0[19]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[1] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[1]),
        .Q(dec_new_block[33]));
  MUXF7 \block_w2_reg_reg[1]_i_1 
       (.I0(\block_w2_reg_reg[1]_0 ),
        .I1(\block_w2_reg[1]_i_3_n_0 ),
        .O(p_0_in__0[1]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[20] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[20]),
        .Q(dec_new_block[52]));
  MUXF7 \block_w2_reg_reg[20]_i_1 
       (.I0(\block_w2_reg_reg[20]_0 ),
        .I1(\block_w2_reg[20]_i_3_n_0 ),
        .O(p_0_in__0[20]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[21] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[21]),
        .Q(dec_new_block[53]));
  MUXF7 \block_w2_reg_reg[21]_i_1 
       (.I0(\block_w2_reg_reg[21]_0 ),
        .I1(\block_w2_reg[21]_i_3_n_0 ),
        .O(p_0_in__0[21]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[22] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[22]),
        .Q(dec_new_block[54]));
  MUXF7 \block_w2_reg_reg[22]_i_1 
       (.I0(\block_w2_reg_reg[22]_0 ),
        .I1(\block_w2_reg[22]_i_3_n_0 ),
        .O(p_0_in__0[22]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[23] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[23]),
        .Q(dec_new_block[55]));
  MUXF7 \block_w2_reg_reg[23]_i_1 
       (.I0(\block_w2_reg_reg[23]_0 ),
        .I1(\block_w2_reg[23]_i_3_n_0 ),
        .O(p_0_in__0[23]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[24] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[24]),
        .Q(dec_new_block[56]));
  MUXF7 \block_w2_reg_reg[24]_i_1 
       (.I0(\block_w2_reg_reg[24]_0 ),
        .I1(\block_w2_reg[24]_i_3_n_0 ),
        .O(p_0_in__0[24]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[25] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[25]),
        .Q(dec_new_block[57]));
  MUXF7 \block_w2_reg_reg[25]_i_1 
       (.I0(\block_w2_reg_reg[25]_0 ),
        .I1(\block_w2_reg[25]_i_3_n_0 ),
        .O(p_0_in__0[25]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[26] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[26]),
        .Q(dec_new_block[58]));
  MUXF7 \block_w2_reg_reg[26]_i_1 
       (.I0(\block_w2_reg[26]_i_2__0_n_0 ),
        .I1(\block_w2_reg[26]_i_3_n_0 ),
        .O(p_0_in__0[26]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[27] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[27]),
        .Q(dec_new_block[59]));
  MUXF7 \block_w2_reg_reg[27]_i_1 
       (.I0(\block_w2_reg[27]_i_2__0_n_0 ),
        .I1(\block_w2_reg[27]_i_3_n_0 ),
        .O(p_0_in__0[27]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[28] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[28]),
        .Q(dec_new_block[60]));
  MUXF7 \block_w2_reg_reg[28]_i_1 
       (.I0(\block_w2_reg_reg[28]_0 ),
        .I1(\block_w2_reg[28]_i_3_n_0 ),
        .O(p_0_in__0[28]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[29] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[29]),
        .Q(dec_new_block[61]));
  MUXF7 \block_w2_reg_reg[29]_i_1 
       (.I0(\block_w2_reg_reg[29]_0 ),
        .I1(\block_w2_reg[29]_i_3_n_0 ),
        .O(p_0_in__0[29]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[2] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[2]),
        .Q(dec_new_block[34]));
  MUXF7 \block_w2_reg_reg[2]_i_1 
       (.I0(\block_w2_reg_reg[2]_0 ),
        .I1(\block_w2_reg[2]_i_3_n_0 ),
        .O(p_0_in__0[2]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[30] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[30]),
        .Q(dec_new_block[62]));
  MUXF7 \block_w2_reg_reg[30]_i_1 
       (.I0(\block_w2_reg_reg[30]_0 ),
        .I1(\block_w2_reg[30]_i_3_n_0 ),
        .O(p_0_in__0[30]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[31] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[31]),
        .Q(dec_new_block[63]));
  MUXF7 \block_w2_reg_reg[31]_i_2 
       (.I0(\block_w2_reg_reg[31]_0 ),
        .I1(\block_w2_reg[31]_i_4_n_0 ),
        .O(p_0_in__0[31]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[3] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[3]),
        .Q(dec_new_block[35]));
  MUXF7 \block_w2_reg_reg[3]_i_1 
       (.I0(\block_w2_reg_reg[3]_0 ),
        .I1(\block_w2_reg[3]_i_3_n_0 ),
        .O(p_0_in__0[3]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[4] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[4]),
        .Q(dec_new_block[36]));
  MUXF7 \block_w2_reg_reg[4]_i_1 
       (.I0(\block_w2_reg_reg[4]_0 ),
        .I1(\block_w2_reg[4]_i_3_n_0 ),
        .O(p_0_in__0[4]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[5] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[5]),
        .Q(dec_new_block[37]));
  MUXF7 \block_w2_reg_reg[5]_i_1 
       (.I0(\block_w2_reg_reg[5]_0 ),
        .I1(\block_w2_reg[5]_i_3_n_0 ),
        .O(p_0_in__0[5]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[6] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[6]),
        .Q(dec_new_block[38]));
  MUXF7 \block_w2_reg_reg[6]_i_1 
       (.I0(\block_w2_reg_reg[6]_0 ),
        .I1(\block_w2_reg[6]_i_3_n_0 ),
        .O(p_0_in__0[6]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[7] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[7]),
        .Q(dec_new_block[39]));
  MUXF7 \block_w2_reg_reg[7]_i_1 
       (.I0(\block_w2_reg_reg[7]_0 ),
        .I1(\block_w2_reg[7]_i_3_n_0 ),
        .O(p_0_in__0[7]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[8] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[8]),
        .Q(dec_new_block[40]));
  MUXF7 \block_w2_reg_reg[8]_i_1 
       (.I0(\block_w2_reg_reg[8]_0 ),
        .I1(\block_w2_reg[8]_i_3_n_0 ),
        .O(p_0_in__0[8]),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[9] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[9]),
        .Q(dec_new_block[41]));
  LUT6 #(
    .INIT(64'hBA10BA1044440000)) 
    \block_w3_reg[0]_i_1 
       (.I0(update_type__0),
        .I1(ready_new),
        .I2(\block_w3_reg_reg[0]_0 ),
        .I3(\block_w3_reg_reg[0]_1 ),
        .I4(p_0_in31_in),
        .I5(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w3_reg[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[10]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[32]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[10]),
        .I5(inv_mixcolumns_return0174_out__63[2]),
        .O(\block_w3_reg[10]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w3_reg[11]_i_2__0 
       (.I0(round_key[0]),
        .I1(dec_new_block[11]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w3_reg[11]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[11]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[33]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[11]),
        .I5(inv_mixcolumns_return0174_out__63[3]),
        .O(\block_w3_reg[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[12]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[34]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[12]),
        .I5(inv_mixcolumns_return0174_out__63[4]),
        .O(\block_w3_reg[12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[13]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[35]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[13]),
        .I5(inv_mixcolumns_return0174_out__63[5]),
        .O(\block_w3_reg[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[14]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[36]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[14]),
        .I5(inv_mixcolumns_return0174_out__63[6]),
        .O(\block_w3_reg[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w3_reg[15]_i_13 
       (.I0(dec_new_block[79]),
        .I1(dec_new_block[111]),
        .I2(dec_new_block[15]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[47]),
        .O(tmp_sboxw[15]));
  LUT4 #(
    .INIT(16'h1000)) 
    \block_w3_reg[15]_i_14 
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[14]),
        .O(tmp_sboxw_0[14]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w3_reg[15]_i_15 
       (.I0(dec_new_block[78]),
        .I1(dec_new_block[110]),
        .I2(dec_new_block[14]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[46]),
        .O(tmp_sboxw[14]));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[15]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[37]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[15]),
        .I5(inv_mixcolumns_return0174_out__63[7]),
        .O(\block_w3_reg[15]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \block_w3_reg[15]_i_8 
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[15]),
        .O(tmp_sboxw_0[15]));
  LUT6 #(
    .INIT(64'hBA10BA1044440000)) 
    \block_w3_reg[16]_i_1 
       (.I0(update_type__0),
        .I1(ready_new),
        .I2(\block_w3_reg_reg[16]_0 ),
        .I3(\block_w3_reg_reg[16]_1 ),
        .I4(op96_in),
        .I5(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w3_reg[16]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \block_w3_reg[16]_i_5 
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .O(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[17]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[15]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[17]),
        .I5(inv_mixcolumns_return0149_out__55[0]),
        .O(\block_w3_reg[17]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w3_reg[18]_i_2__0 
       (.I0(dec_new_block[18]),
        .I1(round_key[1]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w3_reg[18]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[18]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[16]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[18]),
        .I5(inv_mixcolumns_return0149_out__55[1]),
        .O(\block_w3_reg[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[19]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[17]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[19]),
        .I5(inv_mixcolumns_return0149_out__55[2]),
        .O(\block_w3_reg[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[1]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[46]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[1]),
        .I5(inv_mixcolumns_return0198_out__63[0]),
        .O(\block_w3_reg[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[20]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[18]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[20]),
        .I5(inv_mixcolumns_return0149_out__55[3]),
        .O(\block_w3_reg[20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[21]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[19]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[21]),
        .I5(inv_mixcolumns_return0149_out__55[4]),
        .O(\block_w3_reg[21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[22]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[20]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[22]),
        .I5(inv_mixcolumns_return0149_out__55[5]),
        .O(\block_w3_reg[22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w3_reg[23]_i_13 
       (.I0(dec_new_block[87]),
        .I1(dec_new_block[119]),
        .I2(dec_new_block[23]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[55]),
        .O(tmp_sboxw[23]));
  LUT4 #(
    .INIT(16'h1000)) 
    \block_w3_reg[23]_i_14 
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[22]),
        .O(tmp_sboxw_0[22]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w3_reg[23]_i_15 
       (.I0(dec_new_block[86]),
        .I1(dec_new_block[118]),
        .I2(dec_new_block[22]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[54]),
        .O(tmp_sboxw[22]));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[23]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[21]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[23]),
        .I5(inv_mixcolumns_return0149_out__55[6]),
        .O(\block_w3_reg[23]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \block_w3_reg[23]_i_8 
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[23]),
        .O(tmp_sboxw_0[23]));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[24]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[0]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[24]),
        .I5(inv_mixcolumns_return0124_out__47[0]),
        .O(\block_w3_reg[24]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[25]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[1]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[25]),
        .I5(inv_mixcolumns_return0124_out__47[1]),
        .O(\block_w3_reg[25]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w3_reg[26]_i_2__0 
       (.I0(dec_new_block[26]),
        .I1(round_key[2]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w3_reg[26]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[26]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[2]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[26]),
        .I5(inv_mixcolumns_return0124_out__47[2]),
        .O(\block_w3_reg[26]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \block_w3_reg[27]_i_2__0 
       (.I0(dec_new_block[27]),
        .I1(round_key[3]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .O(\block_w3_reg[27]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[27]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[3]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[27]),
        .I5(inv_mixcolumns_return0124_out__47[3]),
        .O(\block_w3_reg[27]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[28]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[4]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[28]),
        .I5(inv_mixcolumns_return0124_out__47[4]),
        .O(\block_w3_reg[28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[29]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[5]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[29]),
        .I5(inv_mixcolumns_return0124_out__47[5]),
        .O(\block_w3_reg[29]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[2]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[47]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[2]),
        .I5(inv_mixcolumns_return0198_out__63[1]),
        .O(\block_w3_reg[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[30]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[6]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[30]),
        .I5(inv_mixcolumns_return0124_out__47[6]),
        .O(\block_w3_reg[30]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h54446666)) 
    \block_w3_reg[31]_i_1 
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(p_0_in[1]),
        .I3(p_0_in[0]),
        .I4(update_type__0),
        .O(block_w3_we));
  LUT4 #(
    .INIT(16'h1000)) 
    \block_w3_reg[31]_i_10__0 
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[31]),
        .O(tmp_sboxw_0[31]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w3_reg[31]_i_15 
       (.I0(dec_new_block[95]),
        .I1(dec_new_block[127]),
        .I2(dec_new_block[31]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[63]),
        .O(tmp_sboxw[31]));
  LUT4 #(
    .INIT(16'h1000)) 
    \block_w3_reg[31]_i_16 
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[30]),
        .O(tmp_sboxw_0[30]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w3_reg[31]_i_17 
       (.I0(dec_new_block[94]),
        .I1(dec_new_block[126]),
        .I2(dec_new_block[30]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[62]),
        .O(tmp_sboxw[30]));
  LUT2 #(
    .INIT(4'hB)) 
    \block_w3_reg[31]_i_3__0 
       (.I0(update_type__0),
        .I1(ready_new),
        .O(\block_w3_reg[31]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[31]_i_5 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[7]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[31]),
        .I5(inv_mixcolumns_return0124_out__47[7]),
        .O(\block_w3_reg[31]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[3]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[48]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[3]),
        .I5(inv_mixcolumns_return0198_out__63[2]),
        .O(\block_w3_reg[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[4]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[49]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[4]),
        .I5(inv_mixcolumns_return0198_out__63[3]),
        .O(\block_w3_reg[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[5]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[50]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[5]),
        .I5(inv_mixcolumns_return0198_out__63[4]),
        .O(\block_w3_reg[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[6]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[51]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[6]),
        .I5(inv_mixcolumns_return0198_out__63[5]),
        .O(\block_w3_reg[6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w3_reg[7]_i_13 
       (.I0(dec_new_block[71]),
        .I1(dec_new_block[103]),
        .I2(dec_new_block[7]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[39]),
        .O(tmp_sboxw[7]));
  LUT4 #(
    .INIT(16'h1000)) 
    \block_w3_reg[7]_i_14 
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[6]),
        .O(tmp_sboxw_0[6]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w3_reg[7]_i_15 
       (.I0(dec_new_block[70]),
        .I1(dec_new_block[102]),
        .I2(dec_new_block[6]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[38]),
        .O(tmp_sboxw[6]));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[7]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[52]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[7]),
        .I5(inv_mixcolumns_return0198_out__63[6]),
        .O(\block_w3_reg[7]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \block_w3_reg[7]_i_8 
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[7]),
        .O(tmp_sboxw_0[7]));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[8]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[30]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(new_sboxw[8]),
        .I5(inv_mixcolumns_return0174_out__63[0]),
        .O(\block_w3_reg[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA80A0800A800080)) 
    \block_w3_reg[9]_i_3 
       (.I0(\FSM_sequential_dec_ctrl_reg_reg[1]_0 ),
        .I1(p_0_out[31]),
        .I2(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I3(update_type__0),
        .I4(\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11 [1]),
        .I5(inv_mixcolumns_return0174_out__63[1]),
        .O(\block_w3_reg[9]_i_3_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[0] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[0]_i_1_n_0 ),
        .Q(dec_new_block[0]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[10] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[10]_i_1_n_0 ),
        .Q(dec_new_block[10]));
  MUXF7 \block_w3_reg_reg[10]_i_1 
       (.I0(\block_w3_reg_reg[10]_0 ),
        .I1(\block_w3_reg[10]_i_3_n_0 ),
        .O(\block_w3_reg_reg[10]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[11] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[11]_i_1_n_0 ),
        .Q(dec_new_block[11]));
  MUXF7 \block_w3_reg_reg[11]_i_1 
       (.I0(\block_w3_reg[11]_i_2__0_n_0 ),
        .I1(\block_w3_reg[11]_i_3_n_0 ),
        .O(\block_w3_reg_reg[11]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[12] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[12]_i_1_n_0 ),
        .Q(dec_new_block[12]));
  MUXF7 \block_w3_reg_reg[12]_i_1 
       (.I0(\block_w3_reg_reg[12]_0 ),
        .I1(\block_w3_reg[12]_i_3_n_0 ),
        .O(\block_w3_reg_reg[12]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[13] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[13]_i_1_n_0 ),
        .Q(dec_new_block[13]));
  MUXF7 \block_w3_reg_reg[13]_i_1 
       (.I0(\block_w3_reg_reg[13]_0 ),
        .I1(\block_w3_reg[13]_i_3_n_0 ),
        .O(\block_w3_reg_reg[13]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[14] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[14]_i_1_n_0 ),
        .Q(dec_new_block[14]));
  MUXF7 \block_w3_reg_reg[14]_i_1 
       (.I0(\block_w3_reg_reg[14]_0 ),
        .I1(\block_w3_reg[14]_i_3_n_0 ),
        .O(\block_w3_reg_reg[14]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[15] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[15]_i_1_n_0 ),
        .Q(dec_new_block[15]));
  MUXF7 \block_w3_reg_reg[15]_i_1 
       (.I0(\block_w3_reg_reg[15]_0 ),
        .I1(\block_w3_reg[15]_i_3_n_0 ),
        .O(\block_w3_reg_reg[15]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[16] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[16]_i_1_n_0 ),
        .Q(dec_new_block[16]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[17] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[17]_i_1_n_0 ),
        .Q(dec_new_block[17]));
  MUXF7 \block_w3_reg_reg[17]_i_1 
       (.I0(\block_w3_reg_reg[17]_0 ),
        .I1(\block_w3_reg[17]_i_3_n_0 ),
        .O(\block_w3_reg_reg[17]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[18] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[18]_i_1_n_0 ),
        .Q(dec_new_block[18]));
  MUXF7 \block_w3_reg_reg[18]_i_1 
       (.I0(\block_w3_reg[18]_i_2__0_n_0 ),
        .I1(\block_w3_reg[18]_i_3_n_0 ),
        .O(\block_w3_reg_reg[18]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[19] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[19]_i_1_n_0 ),
        .Q(dec_new_block[19]));
  MUXF7 \block_w3_reg_reg[19]_i_1 
       (.I0(\block_w3_reg_reg[19]_0 ),
        .I1(\block_w3_reg[19]_i_3_n_0 ),
        .O(\block_w3_reg_reg[19]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[1] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[1]_i_1_n_0 ),
        .Q(dec_new_block[1]));
  MUXF7 \block_w3_reg_reg[1]_i_1 
       (.I0(\block_w3_reg_reg[1]_0 ),
        .I1(\block_w3_reg[1]_i_3_n_0 ),
        .O(\block_w3_reg_reg[1]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[20] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[20]_i_1_n_0 ),
        .Q(dec_new_block[20]));
  MUXF7 \block_w3_reg_reg[20]_i_1 
       (.I0(\block_w3_reg_reg[20]_0 ),
        .I1(\block_w3_reg[20]_i_3_n_0 ),
        .O(\block_w3_reg_reg[20]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[21] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[21]_i_1_n_0 ),
        .Q(dec_new_block[21]));
  MUXF7 \block_w3_reg_reg[21]_i_1 
       (.I0(\block_w3_reg_reg[21]_0 ),
        .I1(\block_w3_reg[21]_i_3_n_0 ),
        .O(\block_w3_reg_reg[21]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[22] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[22]_i_1_n_0 ),
        .Q(dec_new_block[22]));
  MUXF7 \block_w3_reg_reg[22]_i_1 
       (.I0(\block_w3_reg_reg[22]_0 ),
        .I1(\block_w3_reg[22]_i_3_n_0 ),
        .O(\block_w3_reg_reg[22]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[23] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[23]_i_1_n_0 ),
        .Q(dec_new_block[23]));
  MUXF7 \block_w3_reg_reg[23]_i_1 
       (.I0(\block_w3_reg_reg[23]_0 ),
        .I1(\block_w3_reg[23]_i_3_n_0 ),
        .O(\block_w3_reg_reg[23]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[24] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[24]_i_1_n_0 ),
        .Q(dec_new_block[24]));
  MUXF7 \block_w3_reg_reg[24]_i_1 
       (.I0(\block_w3_reg_reg[24]_0 ),
        .I1(\block_w3_reg[24]_i_3_n_0 ),
        .O(\block_w3_reg_reg[24]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[25] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[25]_i_1_n_0 ),
        .Q(dec_new_block[25]));
  MUXF7 \block_w3_reg_reg[25]_i_1 
       (.I0(\block_w3_reg_reg[25]_0 ),
        .I1(\block_w3_reg[25]_i_3_n_0 ),
        .O(\block_w3_reg_reg[25]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[26] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[26]_i_1_n_0 ),
        .Q(dec_new_block[26]));
  MUXF7 \block_w3_reg_reg[26]_i_1 
       (.I0(\block_w3_reg[26]_i_2__0_n_0 ),
        .I1(\block_w3_reg[26]_i_3_n_0 ),
        .O(\block_w3_reg_reg[26]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[27] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[27]_i_1_n_0 ),
        .Q(dec_new_block[27]));
  MUXF7 \block_w3_reg_reg[27]_i_1 
       (.I0(\block_w3_reg[27]_i_2__0_n_0 ),
        .I1(\block_w3_reg[27]_i_3_n_0 ),
        .O(\block_w3_reg_reg[27]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[28] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[28]_i_1_n_0 ),
        .Q(dec_new_block[28]));
  MUXF7 \block_w3_reg_reg[28]_i_1 
       (.I0(\block_w3_reg_reg[28]_0 ),
        .I1(\block_w3_reg[28]_i_3_n_0 ),
        .O(\block_w3_reg_reg[28]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[29] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[29]_i_1_n_0 ),
        .Q(dec_new_block[29]));
  MUXF7 \block_w3_reg_reg[29]_i_1 
       (.I0(\block_w3_reg_reg[29]_0 ),
        .I1(\block_w3_reg[29]_i_3_n_0 ),
        .O(\block_w3_reg_reg[29]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[2] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[2]_i_1_n_0 ),
        .Q(dec_new_block[2]));
  MUXF7 \block_w3_reg_reg[2]_i_1 
       (.I0(\block_w3_reg_reg[2]_0 ),
        .I1(\block_w3_reg[2]_i_3_n_0 ),
        .O(\block_w3_reg_reg[2]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[30] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[30]_i_1_n_0 ),
        .Q(dec_new_block[30]));
  MUXF7 \block_w3_reg_reg[30]_i_1 
       (.I0(\block_w3_reg_reg[30]_0 ),
        .I1(\block_w3_reg[30]_i_3_n_0 ),
        .O(\block_w3_reg_reg[30]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[31] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[31]_i_2_n_0 ),
        .Q(dec_new_block[31]));
  MUXF7 \block_w3_reg_reg[31]_i_2 
       (.I0(\block_w3_reg_reg[31]_0 ),
        .I1(\block_w3_reg[31]_i_5_n_0 ),
        .O(\block_w3_reg_reg[31]_i_2_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[3] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[3]_i_1_n_0 ),
        .Q(dec_new_block[3]));
  MUXF7 \block_w3_reg_reg[3]_i_1 
       (.I0(\block_w3_reg_reg[3]_0 ),
        .I1(\block_w3_reg[3]_i_3_n_0 ),
        .O(\block_w3_reg_reg[3]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[4] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[4]_i_1_n_0 ),
        .Q(dec_new_block[4]));
  MUXF7 \block_w3_reg_reg[4]_i_1 
       (.I0(\block_w3_reg_reg[4]_0 ),
        .I1(\block_w3_reg[4]_i_3_n_0 ),
        .O(\block_w3_reg_reg[4]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[5] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[5]_i_1_n_0 ),
        .Q(dec_new_block[5]));
  MUXF7 \block_w3_reg_reg[5]_i_1 
       (.I0(\block_w3_reg_reg[5]_0 ),
        .I1(\block_w3_reg[5]_i_3_n_0 ),
        .O(\block_w3_reg_reg[5]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[6] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[6]_i_1_n_0 ),
        .Q(dec_new_block[6]));
  MUXF7 \block_w3_reg_reg[6]_i_1 
       (.I0(\block_w3_reg_reg[6]_0 ),
        .I1(\block_w3_reg[6]_i_3_n_0 ),
        .O(\block_w3_reg_reg[6]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[7] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[7]_i_1_n_0 ),
        .Q(dec_new_block[7]));
  MUXF7 \block_w3_reg_reg[7]_i_1 
       (.I0(\block_w3_reg_reg[7]_0 ),
        .I1(\block_w3_reg[7]_i_3_n_0 ),
        .O(\block_w3_reg_reg[7]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[8] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[8]_i_1_n_0 ),
        .Q(dec_new_block[8]));
  MUXF7 \block_w3_reg_reg[8]_i_1 
       (.I0(\block_w3_reg_reg[8]_0 ),
        .I1(\block_w3_reg[8]_i_3_n_0 ),
        .O(\block_w3_reg_reg[8]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[9] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg_reg[9]_i_1_n_0 ),
        .Q(dec_new_block[9]));
  MUXF7 \block_w3_reg_reg[9]_i_1 
       (.I0(\block_w3_reg_reg[9]_0 ),
        .I1(\block_w3_reg[9]_i_3_n_0 ),
        .O(\block_w3_reg_reg[9]_i_1_n_0 ),
        .S(\block_w3_reg[31]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hFA244CC2C4F6F54A)) 
    g0_b0
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g0_b0_n_0));
  LUT6 #(
    .INIT(64'hFA244CC2C4F6F54A)) 
    g0_b0__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g0_b0__0_n_0));
  LUT6 #(
    .INIT(64'hFA244CC2C4F6F54A)) 
    g0_b0__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g0_b0__1_n_0));
  LUT6 #(
    .INIT(64'hFA244CC2C4F6F54A)) 
    g0_b0__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g0_b0__2_n_0));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_1
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[24]),
        .O(tmp_sboxw_0[24]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_10
       (.I0(dec_new_block[64]),
        .I1(dec_new_block[96]),
        .I2(dec_new_block[0]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[32]),
        .O(tmp_sboxw[0]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_10__0
       (.I0(dec_new_block[75]),
        .I1(dec_new_block[107]),
        .I2(dec_new_block[11]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[43]),
        .O(tmp_sboxw[11]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_10__1
       (.I0(dec_new_block[83]),
        .I1(dec_new_block[115]),
        .I2(dec_new_block[19]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[51]),
        .O(tmp_sboxw[19]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_10__2
       (.I0(dec_new_block[91]),
        .I1(dec_new_block[123]),
        .I2(dec_new_block[27]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[59]),
        .O(tmp_sboxw[27]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_11
       (.I0(dec_new_block[65]),
        .I1(dec_new_block[97]),
        .I2(dec_new_block[1]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[33]),
        .O(tmp_sboxw[1]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_11__0
       (.I0(dec_new_block[76]),
        .I1(dec_new_block[108]),
        .I2(dec_new_block[12]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[44]),
        .O(tmp_sboxw[12]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_11__1
       (.I0(dec_new_block[84]),
        .I1(dec_new_block[116]),
        .I2(dec_new_block[20]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[52]),
        .O(tmp_sboxw[20]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_11__2
       (.I0(dec_new_block[92]),
        .I1(dec_new_block[124]),
        .I2(dec_new_block[28]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[60]),
        .O(tmp_sboxw[28]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_12
       (.I0(dec_new_block[66]),
        .I1(dec_new_block[98]),
        .I2(dec_new_block[2]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[34]),
        .O(tmp_sboxw[2]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_12__0
       (.I0(dec_new_block[77]),
        .I1(dec_new_block[109]),
        .I2(dec_new_block[13]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[45]),
        .O(tmp_sboxw[13]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_12__1
       (.I0(dec_new_block[85]),
        .I1(dec_new_block[117]),
        .I2(dec_new_block[21]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[53]),
        .O(tmp_sboxw[21]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_12__2
       (.I0(dec_new_block[93]),
        .I1(dec_new_block[125]),
        .I2(dec_new_block[29]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[61]),
        .O(tmp_sboxw[29]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_13
       (.I0(dec_new_block[67]),
        .I1(dec_new_block[99]),
        .I2(dec_new_block[3]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[35]),
        .O(tmp_sboxw[3]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_14
       (.I0(dec_new_block[68]),
        .I1(dec_new_block[100]),
        .I2(dec_new_block[4]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[36]),
        .O(tmp_sboxw[4]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_15
       (.I0(dec_new_block[69]),
        .I1(dec_new_block[101]),
        .I2(dec_new_block[5]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[37]),
        .O(tmp_sboxw[5]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_1__0
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[16]),
        .O(tmp_sboxw_0[16]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_1__1
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[8]),
        .O(tmp_sboxw_0[8]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_1__2
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[0]),
        .O(tmp_sboxw_0[0]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_2
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[25]),
        .O(tmp_sboxw_0[25]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_2__0
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[17]),
        .O(tmp_sboxw_0[17]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_2__1
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[9]),
        .O(tmp_sboxw_0[9]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_2__2
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[1]),
        .O(tmp_sboxw_0[1]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_3
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[26]),
        .O(tmp_sboxw_0[26]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_3__0
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[18]),
        .O(tmp_sboxw_0[18]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_3__1
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[10]),
        .O(tmp_sboxw_0[10]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_3__2
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[2]),
        .O(tmp_sboxw_0[2]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_4
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[27]),
        .O(tmp_sboxw_0[27]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_4__0
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[19]),
        .O(tmp_sboxw_0[19]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_4__1
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[11]),
        .O(tmp_sboxw_0[11]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_4__2
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[3]),
        .O(tmp_sboxw_0[3]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_5
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[28]),
        .O(tmp_sboxw_0[28]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_5__0
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[20]),
        .O(tmp_sboxw_0[20]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_5__1
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[12]),
        .O(tmp_sboxw_0[12]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_5__2
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[4]),
        .O(tmp_sboxw_0[4]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_6
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[29]),
        .O(tmp_sboxw_0[29]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_6__0
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[21]),
        .O(tmp_sboxw_0[21]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_6__1
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[13]),
        .O(tmp_sboxw_0[13]));
  LUT4 #(
    .INIT(16'h1000)) 
    g0_b0_i_6__2
       (.I0(ready_new),
        .I1(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ),
        .I2(update_type__0),
        .I3(tmp_sboxw[5]),
        .O(tmp_sboxw_0[5]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    g0_b0_i_7
       (.I0(dec_ctrl_reg),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[3]),
        .I5(sword_ctr_rst),
        .O(ready_new));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_7__0
       (.I0(dec_new_block[72]),
        .I1(dec_new_block[104]),
        .I2(dec_new_block[8]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[40]),
        .O(tmp_sboxw[8]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_7__1
       (.I0(dec_new_block[80]),
        .I1(dec_new_block[112]),
        .I2(dec_new_block[16]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[48]),
        .O(tmp_sboxw[16]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_7__2
       (.I0(dec_new_block[88]),
        .I1(dec_new_block[120]),
        .I2(dec_new_block[24]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[56]),
        .O(tmp_sboxw[24]));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA2)) 
    g0_b0_i_8
       (.I0(sword_ctr_rst),
        .I1(dec_ctrl_reg),
        .I2(Q[2]),
        .I3(Q[1]),
        .I4(Q[0]),
        .I5(Q[3]),
        .O(\FSM_sequential_dec_ctrl_reg_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_8__0
       (.I0(dec_new_block[73]),
        .I1(dec_new_block[105]),
        .I2(dec_new_block[9]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[41]),
        .O(tmp_sboxw[9]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_8__1
       (.I0(dec_new_block[81]),
        .I1(dec_new_block[113]),
        .I2(dec_new_block[17]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[49]),
        .O(tmp_sboxw[17]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_8__2
       (.I0(dec_new_block[89]),
        .I1(dec_new_block[121]),
        .I2(dec_new_block[25]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[57]),
        .O(tmp_sboxw[25]));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA2)) 
    g0_b0_i_9
       (.I0(dec_ctrl_reg),
        .I1(sword_ctr_rst),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(Q[1]),
        .I5(Q[2]),
        .O(update_type__0));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_9__0
       (.I0(dec_new_block[74]),
        .I1(dec_new_block[106]),
        .I2(dec_new_block[10]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[42]),
        .O(tmp_sboxw[10]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_9__1
       (.I0(dec_new_block[82]),
        .I1(dec_new_block[114]),
        .I2(dec_new_block[18]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[50]),
        .O(tmp_sboxw[18]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_9__2
       (.I0(dec_new_block[90]),
        .I1(dec_new_block[122]),
        .I2(dec_new_block[26]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(dec_new_block[58]),
        .O(tmp_sboxw[26]));
  LUT6 #(
    .INIT(64'h278AF97AA6FAED25)) 
    g0_b1
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g0_b1_n_0));
  LUT6 #(
    .INIT(64'h278AF97AA6FAED25)) 
    g0_b1__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g0_b1__0_n_0));
  LUT6 #(
    .INIT(64'h278AF97AA6FAED25)) 
    g0_b1__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g0_b1__1_n_0));
  LUT6 #(
    .INIT(64'h278AF97AA6FAED25)) 
    g0_b1__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g0_b1__2_n_0));
  LUT6 #(
    .INIT(64'h914A87953BE14968)) 
    g0_b2
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g0_b2_n_0));
  LUT6 #(
    .INIT(64'h914A87953BE14968)) 
    g0_b2__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g0_b2__0_n_0));
  LUT6 #(
    .INIT(64'h914A87953BE14968)) 
    g0_b2__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g0_b2__1_n_0));
  LUT6 #(
    .INIT(64'h914A87953BE14968)) 
    g0_b2__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g0_b2__2_n_0));
  LUT6 #(
    .INIT(64'h3A33AB82E2758986)) 
    g0_b3
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g0_b3_n_0));
  LUT6 #(
    .INIT(64'h3A33AB82E2758986)) 
    g0_b3__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g0_b3__0_n_0));
  LUT6 #(
    .INIT(64'h3A33AB82E2758986)) 
    g0_b3__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g0_b3__1_n_0));
  LUT6 #(
    .INIT(64'h3A33AB82E2758986)) 
    g0_b3__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g0_b3__2_n_0));
  LUT6 #(
    .INIT(64'h43A0248F2155E9B9)) 
    g0_b4
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g0_b4_n_0));
  LUT6 #(
    .INIT(64'h43A0248F2155E9B9)) 
    g0_b4__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g0_b4__0_n_0));
  LUT6 #(
    .INIT(64'h43A0248F2155E9B9)) 
    g0_b4__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g0_b4__1_n_0));
  LUT6 #(
    .INIT(64'h43A0248F2155E9B9)) 
    g0_b4__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g0_b4__2_n_0));
  LUT6 #(
    .INIT(64'h95DE21DA4167A5F4)) 
    g0_b5
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g0_b5_n_0));
  LUT6 #(
    .INIT(64'h95DE21DA4167A5F4)) 
    g0_b5__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g0_b5__0_n_0));
  LUT6 #(
    .INIT(64'h95DE21DA4167A5F4)) 
    g0_b5__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g0_b5__1_n_0));
  LUT6 #(
    .INIT(64'h95DE21DA4167A5F4)) 
    g0_b5__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g0_b5__2_n_0));
  LUT6 #(
    .INIT(64'h5B28F323FC43E20D)) 
    g0_b6
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g0_b6_n_0));
  LUT6 #(
    .INIT(64'h5B28F323FC43E20D)) 
    g0_b6__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g0_b6__0_n_0));
  LUT6 #(
    .INIT(64'h5B28F323FC43E20D)) 
    g0_b6__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g0_b6__1_n_0));
  LUT6 #(
    .INIT(64'h5B28F323FC43E20D)) 
    g0_b6__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g0_b6__2_n_0));
  LUT6 #(
    .INIT(64'h64A46534F2DAFD48)) 
    g0_b7
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g0_b7_n_0));
  LUT6 #(
    .INIT(64'h64A46534F2DAFD48)) 
    g0_b7__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g0_b7__0_n_0));
  LUT6 #(
    .INIT(64'h64A46534F2DAFD48)) 
    g0_b7__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g0_b7__1_n_0));
  LUT6 #(
    .INIT(64'h64A46534F2DAFD48)) 
    g0_b7__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g0_b7__2_n_0));
  LUT6 #(
    .INIT(64'hBF6869447A703000)) 
    g1_b0
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g1_b0_n_0));
  LUT6 #(
    .INIT(64'hBF6869447A703000)) 
    g1_b0__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g1_b0__0_n_0));
  LUT6 #(
    .INIT(64'hBF6869447A703000)) 
    g1_b0__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g1_b0__1_n_0));
  LUT6 #(
    .INIT(64'hBF6869447A703000)) 
    g1_b0__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g1_b0__2_n_0));
  LUT6 #(
    .INIT(64'hEAFCA1C41D80C095)) 
    g1_b1
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g1_b1_n_0));
  LUT6 #(
    .INIT(64'hEAFCA1C41D80C095)) 
    g1_b1__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g1_b1__0_n_0));
  LUT6 #(
    .INIT(64'hEAFCA1C41D80C095)) 
    g1_b1__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g1_b1__1_n_0));
  LUT6 #(
    .INIT(64'hEAFCA1C41D80C095)) 
    g1_b1__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g1_b1__2_n_0));
  LUT6 #(
    .INIT(64'h066ECB30FF317F9C)) 
    g1_b2
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g1_b2_n_0));
  LUT6 #(
    .INIT(64'h066ECB30FF317F9C)) 
    g1_b2__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g1_b2__0_n_0));
  LUT6 #(
    .INIT(64'h066ECB30FF317F9C)) 
    g1_b2__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g1_b2__1_n_0));
  LUT6 #(
    .INIT(64'h066ECB30FF317F9C)) 
    g1_b2__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g1_b2__2_n_0));
  LUT6 #(
    .INIT(64'hC67E14B661F51C62)) 
    g1_b3
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g1_b3_n_0));
  LUT6 #(
    .INIT(64'hC67E14B661F51C62)) 
    g1_b3__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g1_b3__0_n_0));
  LUT6 #(
    .INIT(64'hC67E14B661F51C62)) 
    g1_b3__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g1_b3__1_n_0));
  LUT6 #(
    .INIT(64'hC67E14B661F51C62)) 
    g1_b3__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g1_b3__2_n_0));
  LUT6 #(
    .INIT(64'h242535634BDAD5C7)) 
    g1_b4
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g1_b4_n_0));
  LUT6 #(
    .INIT(64'h242535634BDAD5C7)) 
    g1_b4__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g1_b4__0_n_0));
  LUT6 #(
    .INIT(64'h242535634BDAD5C7)) 
    g1_b4__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g1_b4__1_n_0));
  LUT6 #(
    .INIT(64'h242535634BDAD5C7)) 
    g1_b4__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g1_b4__2_n_0));
  LUT6 #(
    .INIT(64'h862233241073622F)) 
    g1_b5
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g1_b5_n_0));
  LUT6 #(
    .INIT(64'h862233241073622F)) 
    g1_b5__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g1_b5__0_n_0));
  LUT6 #(
    .INIT(64'h862233241073622F)) 
    g1_b5__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g1_b5__1_n_0));
  LUT6 #(
    .INIT(64'h862233241073622F)) 
    g1_b5__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g1_b5__2_n_0));
  LUT6 #(
    .INIT(64'h811147420DBF3D2F)) 
    g1_b6
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g1_b6_n_0));
  LUT6 #(
    .INIT(64'h811147420DBF3D2F)) 
    g1_b6__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g1_b6__0_n_0));
  LUT6 #(
    .INIT(64'h811147420DBF3D2F)) 
    g1_b6__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g1_b6__1_n_0));
  LUT6 #(
    .INIT(64'h811147420DBF3D2F)) 
    g1_b6__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g1_b6__2_n_0));
  LUT6 #(
    .INIT(64'h47193377F0F0CB56)) 
    g1_b7
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g1_b7_n_0));
  LUT6 #(
    .INIT(64'h47193377F0F0CB56)) 
    g1_b7__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g1_b7__0_n_0));
  LUT6 #(
    .INIT(64'h47193377F0F0CB56)) 
    g1_b7__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g1_b7__1_n_0));
  LUT6 #(
    .INIT(64'h47193377F0F0CB56)) 
    g1_b7__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g1_b7__2_n_0));
  LUT6 #(
    .INIT(64'h224883FB66F0853E)) 
    g2_b0
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g2_b0_n_0));
  LUT6 #(
    .INIT(64'h224883FB66F0853E)) 
    g2_b0__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g2_b0__0_n_0));
  LUT6 #(
    .INIT(64'h224883FB66F0853E)) 
    g2_b0__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g2_b0__1_n_0));
  LUT6 #(
    .INIT(64'h224883FB66F0853E)) 
    g2_b0__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g2_b0__2_n_0));
  LUT6 #(
    .INIT(64'h4B3EDF05C519CFB1)) 
    g2_b1
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g2_b1_n_0));
  LUT6 #(
    .INIT(64'h4B3EDF05C519CFB1)) 
    g2_b1__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g2_b1__0_n_0));
  LUT6 #(
    .INIT(64'h4B3EDF05C519CFB1)) 
    g2_b1__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g2_b1__1_n_0));
  LUT6 #(
    .INIT(64'h4B3EDF05C519CFB1)) 
    g2_b1__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g2_b1__2_n_0));
  LUT6 #(
    .INIT(64'hA8174B51F4F76D70)) 
    g2_b2
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g2_b2_n_0));
  LUT6 #(
    .INIT(64'hA8174B51F4F76D70)) 
    g2_b2__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g2_b2__0_n_0));
  LUT6 #(
    .INIT(64'hA8174B51F4F76D70)) 
    g2_b2__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g2_b2__1_n_0));
  LUT6 #(
    .INIT(64'hA8174B51F4F76D70)) 
    g2_b2__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g2_b2__2_n_0));
  LUT6 #(
    .INIT(64'h7B4DF9B4DA220CD1)) 
    g2_b3
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g2_b3_n_0));
  LUT6 #(
    .INIT(64'h7B4DF9B4DA220CD1)) 
    g2_b3__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g2_b3__0_n_0));
  LUT6 #(
    .INIT(64'h7B4DF9B4DA220CD1)) 
    g2_b3__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g2_b3__1_n_0));
  LUT6 #(
    .INIT(64'h7B4DF9B4DA220CD1)) 
    g2_b3__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g2_b3__2_n_0));
  LUT6 #(
    .INIT(64'hDB67E21E7645B347)) 
    g2_b4
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g2_b4_n_0));
  LUT6 #(
    .INIT(64'hDB67E21E7645B347)) 
    g2_b4__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g2_b4__0_n_0));
  LUT6 #(
    .INIT(64'hDB67E21E7645B347)) 
    g2_b4__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g2_b4__1_n_0));
  LUT6 #(
    .INIT(64'hDB67E21E7645B347)) 
    g2_b4__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g2_b4__2_n_0));
  LUT6 #(
    .INIT(64'h98C5572AAF7EF2A1)) 
    g2_b5
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g2_b5_n_0));
  LUT6 #(
    .INIT(64'h98C5572AAF7EF2A1)) 
    g2_b5__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g2_b5__0_n_0));
  LUT6 #(
    .INIT(64'h98C5572AAF7EF2A1)) 
    g2_b5__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g2_b5__1_n_0));
  LUT6 #(
    .INIT(64'h98C5572AAF7EF2A1)) 
    g2_b5__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g2_b5__2_n_0));
  LUT6 #(
    .INIT(64'hFE7B054BEB14DEF8)) 
    g2_b6
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g2_b6_n_0));
  LUT6 #(
    .INIT(64'hFE7B054BEB14DEF8)) 
    g2_b6__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g2_b6__0_n_0));
  LUT6 #(
    .INIT(64'hFE7B054BEB14DEF8)) 
    g2_b6__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g2_b6__1_n_0));
  LUT6 #(
    .INIT(64'hFE7B054BEB14DEF8)) 
    g2_b6__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g2_b6__2_n_0));
  LUT6 #(
    .INIT(64'hAF3152C24BB37FC2)) 
    g2_b7
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g2_b7_n_0));
  LUT6 #(
    .INIT(64'hAF3152C24BB37FC2)) 
    g2_b7__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g2_b7__0_n_0));
  LUT6 #(
    .INIT(64'hAF3152C24BB37FC2)) 
    g2_b7__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g2_b7__1_n_0));
  LUT6 #(
    .INIT(64'hAF3152C24BB37FC2)) 
    g2_b7__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g2_b7__2_n_0));
  LUT6 #(
    .INIT(64'hBB23F64CBBBE99EB)) 
    g3_b0
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g3_b0_n_0));
  LUT6 #(
    .INIT(64'hBB23F64CBBBE99EB)) 
    g3_b0__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g3_b0__0_n_0));
  LUT6 #(
    .INIT(64'hBB23F64CBBBE99EB)) 
    g3_b0__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g3_b0__1_n_0));
  LUT6 #(
    .INIT(64'hBB23F64CBBBE99EB)) 
    g3_b0__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g3_b0__2_n_0));
  LUT6 #(
    .INIT(64'h08FB36349C449269)) 
    g3_b1
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g3_b1_n_0));
  LUT6 #(
    .INIT(64'h08FB36349C449269)) 
    g3_b1__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g3_b1__0_n_0));
  LUT6 #(
    .INIT(64'h08FB36349C449269)) 
    g3_b1__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g3_b1__1_n_0));
  LUT6 #(
    .INIT(64'h08FB36349C449269)) 
    g3_b1__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g3_b1__2_n_0));
  LUT6 #(
    .INIT(64'hD4ED0858CBA4D063)) 
    g3_b2
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g3_b2_n_0));
  LUT6 #(
    .INIT(64'hD4ED0858CBA4D063)) 
    g3_b2__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g3_b2__0_n_0));
  LUT6 #(
    .INIT(64'hD4ED0858CBA4D063)) 
    g3_b2__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g3_b2__1_n_0));
  LUT6 #(
    .INIT(64'hD4ED0858CBA4D063)) 
    g3_b2__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g3_b2__2_n_0));
  LUT6 #(
    .INIT(64'hC21A4F3CEDDCC817)) 
    g3_b3
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g3_b3_n_0));
  LUT6 #(
    .INIT(64'hC21A4F3CEDDCC817)) 
    g3_b3__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g3_b3__0_n_0));
  LUT6 #(
    .INIT(64'hC21A4F3CEDDCC817)) 
    g3_b3__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g3_b3__1_n_0));
  LUT6 #(
    .INIT(64'hC21A4F3CEDDCC817)) 
    g3_b3__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g3_b3__2_n_0));
  LUT6 #(
    .INIT(64'h94796CC45C368F8B)) 
    g3_b4
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g3_b4_n_0));
  LUT6 #(
    .INIT(64'h94796CC45C368F8B)) 
    g3_b4__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g3_b4__0_n_0));
  LUT6 #(
    .INIT(64'h94796CC45C368F8B)) 
    g3_b4__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g3_b4__1_n_0));
  LUT6 #(
    .INIT(64'h94796CC45C368F8B)) 
    g3_b4__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g3_b4__2_n_0));
  LUT6 #(
    .INIT(64'hABBA8EF7872D518C)) 
    g3_b5
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g3_b5_n_0));
  LUT6 #(
    .INIT(64'hABBA8EF7872D518C)) 
    g3_b5__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g3_b5__0_n_0));
  LUT6 #(
    .INIT(64'hABBA8EF7872D518C)) 
    g3_b5__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g3_b5__1_n_0));
  LUT6 #(
    .INIT(64'hABBA8EF7872D518C)) 
    g3_b5__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g3_b5__2_n_0));
  LUT6 #(
    .INIT(64'h9B68A34AA647C842)) 
    g3_b6
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g3_b6_n_0));
  LUT6 #(
    .INIT(64'h9B68A34AA647C842)) 
    g3_b6__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g3_b6__0_n_0));
  LUT6 #(
    .INIT(64'h9B68A34AA647C842)) 
    g3_b6__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g3_b6__1_n_0));
  LUT6 #(
    .INIT(64'h9B68A34AA647C842)) 
    g3_b6__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g3_b6__2_n_0));
  LUT6 #(
    .INIT(64'h015057D3FA286156)) 
    g3_b7
       (.I0(tmp_sboxw_0[0]),
        .I1(tmp_sboxw_0[1]),
        .I2(tmp_sboxw_0[2]),
        .I3(tmp_sboxw_0[3]),
        .I4(tmp_sboxw_0[4]),
        .I5(tmp_sboxw_0[5]),
        .O(g3_b7_n_0));
  LUT6 #(
    .INIT(64'h015057D3FA286156)) 
    g3_b7__0
       (.I0(tmp_sboxw_0[8]),
        .I1(tmp_sboxw_0[9]),
        .I2(tmp_sboxw_0[10]),
        .I3(tmp_sboxw_0[11]),
        .I4(tmp_sboxw_0[12]),
        .I5(tmp_sboxw_0[13]),
        .O(g3_b7__0_n_0));
  LUT6 #(
    .INIT(64'h015057D3FA286156)) 
    g3_b7__1
       (.I0(tmp_sboxw_0[16]),
        .I1(tmp_sboxw_0[17]),
        .I2(tmp_sboxw_0[18]),
        .I3(tmp_sboxw_0[19]),
        .I4(tmp_sboxw_0[20]),
        .I5(tmp_sboxw_0[21]),
        .O(g3_b7__1_n_0));
  LUT6 #(
    .INIT(64'h015057D3FA286156)) 
    g3_b7__2
       (.I0(tmp_sboxw_0[24]),
        .I1(tmp_sboxw_0[25]),
        .I2(tmp_sboxw_0[26]),
        .I3(tmp_sboxw_0[27]),
        .I4(tmp_sboxw_0[28]),
        .I5(tmp_sboxw_0[29]),
        .O(g3_b7__2_n_0));
  switch_elements_aes_inv_sbox inv_sbox_inst
       (.\block_w3_reg_reg[0]_i_8_0 (g0_b0_n_0),
        .\block_w3_reg_reg[0]_i_8_1 (g1_b0_n_0),
        .\block_w3_reg_reg[0]_i_8_2 (g2_b0_n_0),
        .\block_w3_reg_reg[0]_i_8_3 (g3_b0_n_0),
        .\block_w3_reg_reg[1]_i_5_0 (g0_b1_n_0),
        .\block_w3_reg_reg[1]_i_5_1 (g1_b1_n_0),
        .\block_w3_reg_reg[1]_i_5_2 (g2_b1_n_0),
        .\block_w3_reg_reg[1]_i_5_3 (g3_b1_n_0),
        .\block_w3_reg_reg[2]_i_6_0 (g0_b2_n_0),
        .\block_w3_reg_reg[2]_i_6_1 (g1_b2_n_0),
        .\block_w3_reg_reg[2]_i_6_2 (g2_b2_n_0),
        .\block_w3_reg_reg[2]_i_6_3 (g3_b2_n_0),
        .\block_w3_reg_reg[3]_i_5_0 (g0_b3_n_0),
        .\block_w3_reg_reg[3]_i_5_1 (g1_b3_n_0),
        .\block_w3_reg_reg[3]_i_5_2 (g2_b3_n_0),
        .\block_w3_reg_reg[3]_i_5_3 (g3_b3_n_0),
        .\block_w3_reg_reg[4]_i_5_0 (g0_b4_n_0),
        .\block_w3_reg_reg[4]_i_5_1 (g1_b4_n_0),
        .\block_w3_reg_reg[4]_i_5_2 (g2_b4_n_0),
        .\block_w3_reg_reg[4]_i_5_3 (g3_b4_n_0),
        .\block_w3_reg_reg[5]_i_6_0 (g0_b5_n_0),
        .\block_w3_reg_reg[5]_i_6_1 (g1_b5_n_0),
        .\block_w3_reg_reg[5]_i_6_2 (g2_b5_n_0),
        .\block_w3_reg_reg[5]_i_6_3 (g3_b5_n_0),
        .\block_w3_reg_reg[6]_i_6_0 (g0_b6_n_0),
        .\block_w3_reg_reg[6]_i_6_1 (g1_b6_n_0),
        .\block_w3_reg_reg[6]_i_6_2 (g2_b6_n_0),
        .\block_w3_reg_reg[6]_i_6_3 (g3_b6_n_0),
        .\block_w3_reg_reg[7]_i_6_0 (g0_b7_n_0),
        .\block_w3_reg_reg[7]_i_6_1 (g1_b7_n_0),
        .\block_w3_reg_reg[7]_i_6_2 (g2_b7_n_0),
        .\block_w3_reg_reg[7]_i_6_3 (g3_b7_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_0 (g0_b2__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_1 (g1_b2__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_2 (g2_b2__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_3 (g3_b2__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_0 (g0_b3__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_1 (g1_b3__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_2 (g2_b3__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_3 (g3_b3__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_0 (g0_b4__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_1 (g1_b4__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_2 (g2_b4__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_3 (g3_b4__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_0 (g0_b5__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_1 (g1_b5__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_2 (g2_b5__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_3 (g3_b5__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_0 (g0_b6__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_1 (g1_b6__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_2 (g2_b6__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_3 (g3_b6__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_0 (g0_b7__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_1 (g1_b7__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_2 (g2_b7__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_3 (g3_b7__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_0 (g0_b0__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_1 (g1_b0__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_2 (g2_b0__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_3 (g3_b0__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_0 (g0_b1__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_1 (g1_b1__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_2 (g2_b1__0_n_0),
        .\inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_3 (g3_b1__0_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11_0 (\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11 ),
        .\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_0 (g0_b0__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_1 (g1_b0__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_2 (g2_b0__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_3 (g3_b0__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_0 (g0_b1__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_1 (g1_b1__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_2 (g2_b1__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_3 (g3_b1__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_0 (g0_b2__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_1 (g1_b2__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_2 (g2_b2__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_3 (g3_b2__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_0 (g0_b3__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_1 (g1_b3__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_2 (g2_b3__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_3 (g3_b3__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_0 (g0_b4__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_1 (g1_b4__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_2 (g2_b4__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_3 (g3_b4__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_0 (g0_b5__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_1 (g1_b5__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_2 (g2_b5__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_3 (g3_b5__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_0 (g0_b6__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_1 (g1_b6__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_2 (g2_b6__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_3 (g3_b6__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_0 (g0_b7__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_1 (g1_b7__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_2 (g2_b7__1_n_0),
        .\inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_3 (g3_b7__1_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_0 (g0_b0__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_1 (g1_b0__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_2 (g2_b0__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_3 (g3_b0__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_0 (g0_b1__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_1 (g1_b1__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_2 (g2_b1__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_3 (g3_b1__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_0 (g0_b2__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_1 (g1_b2__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_2 (g2_b2__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_3 (g3_b2__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_0 (g0_b3__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_1 (g1_b3__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_2 (g2_b3__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_3 (g3_b3__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_0 (g0_b4__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_1 (g1_b4__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_2 (g2_b4__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_3 (g3_b4__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_0 (g0_b5__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_1 (g1_b5__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_2 (g2_b5__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_3 (g3_b5__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_0 (g0_b6__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_1 (g1_b6__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_2 (g2_b6__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_3 (g3_b6__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_0 (g0_b7__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_1 (g1_b7__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_2 (g2_b7__2_n_0),
        .\inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_3 (g3_b7__2_n_0),
        .new_sboxw({new_sboxw[31:17],new_sboxw[15:10],new_sboxw[8:1]}),
        .tmp_sboxw_0({tmp_sboxw_0[31:30],tmp_sboxw_0[23:22],tmp_sboxw_0[15:14],tmp_sboxw_0[7:6]}));
  LUT6 #(
    .INIT(64'hFFFFFCFF44440000)) 
    ready_reg_i_1__0
       (.I0(ready_reg_i_2_n_0),
        .I1(sword_ctr_rst),
        .I2(p_1_in[1]),
        .I3(p_1_in[0]),
        .I4(dec_ctrl_reg),
        .I5(dec_ready),
        .O(ready_reg_i_1__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    ready_reg_i_2
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(Q[3]),
        .O(ready_reg_i_2_n_0));
  FDPE #(
    .INIT(1'b1)) 
    ready_reg_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(ready_reg_i_1__0_n_0),
        .PRE(rst_i),
        .Q(dec_ready));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT4 #(
    .INIT(16'h0800)) 
    \round_ctr_reg[0]_i_1__1 
       (.I0(p_0_in[0]),
        .I1(p_0_in[1]),
        .I2(Q[0]),
        .I3(dec_ctrl_reg),
        .O(round_ctr_new[0]));
  LUT6 #(
    .INIT(64'hF8F0F0F8F0F0F0F0)) 
    \round_ctr_reg[1]_i_1__1 
       (.I0(p_0_in[0]),
        .I1(p_0_in[1]),
        .I2(round_ctr_set__1),
        .I3(Q[0]),
        .I4(Q[1]),
        .I5(dec_ctrl_reg),
        .O(round_ctr_new[1]));
  LUT6 #(
    .INIT(64'hB888B888B88888B8)) 
    \round_ctr_reg[2]_i_1__1 
       (.I0(p_1_in[2]),
        .I1(round_ctr_set__1),
        .I2(round_ctr_dec__1),
        .I3(Q[2]),
        .I4(Q[0]),
        .I5(Q[1]),
        .O(round_ctr_new[2]));
  LUT6 #(
    .INIT(64'h00000000F2020202)) 
    \round_ctr_reg[3]_i_1__1 
       (.I0(p_1_in[0]),
        .I1(p_1_in[1]),
        .I2(dec_ctrl_reg),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(sword_ctr_rst),
        .O(round_ctr_we));
  LUT6 #(
    .INIT(64'hFFFEAAABAAAAAAAA)) 
    \round_ctr_reg[3]_i_2__1 
       (.I0(round_ctr_set__1),
        .I1(Q[2]),
        .I2(Q[0]),
        .I3(Q[1]),
        .I4(Q[3]),
        .I5(round_ctr_dec__1),
        .O(round_ctr_new[3]));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \round_ctr_reg[3]_i_3__0 
       (.I0(p_1_in[1]),
        .I1(p_1_in[0]),
        .I2(sword_ctr_rst),
        .I3(dec_ctrl_reg),
        .O(round_ctr_set__1));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT4 #(
    .INIT(16'h4000)) 
    \round_ctr_reg[3]_i_4 
       (.I0(sword_ctr_rst),
        .I1(p_0_in[0]),
        .I2(p_0_in[1]),
        .I3(dec_ctrl_reg),
        .O(round_ctr_dec__1));
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[0] 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(round_ctr_new[0]),
        .Q(Q[0]));
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[1] 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(round_ctr_new[1]),
        .Q(Q[1]));
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[2] 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(round_ctr_new[2]),
        .Q(Q[2]));
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[3] 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(round_ctr_new[3]),
        .Q(Q[3]));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \sword_ctr_reg[0]_i_1__0 
       (.I0(p_0_in[0]),
        .I1(dec_ctrl_reg),
        .I2(sword_ctr_rst),
        .O(sword_ctr_new[0]));
  LUT2 #(
    .INIT(4'hE)) 
    \sword_ctr_reg[1]_i_1__0 
       (.I0(sword_ctr_rst),
        .I1(dec_ctrl_reg),
        .O(sword_ctr_we));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT4 #(
    .INIT(16'h0060)) 
    \sword_ctr_reg[1]_i_2__0 
       (.I0(p_0_in[0]),
        .I1(p_0_in[1]),
        .I2(dec_ctrl_reg),
        .I3(sword_ctr_rst),
        .O(sword_ctr_new[1]));
  FDCE #(
    .INIT(1'b0)) 
    \sword_ctr_reg_reg[0] 
       (.C(clk_i),
        .CE(sword_ctr_we),
        .CLR(rst_i),
        .D(sword_ctr_new[0]),
        .Q(p_0_in[0]));
  FDCE #(
    .INIT(1'b0)) 
    \sword_ctr_reg_reg[1] 
       (.C(clk_i),
        .CE(sword_ctr_we),
        .CLR(rst_i),
        .D(sword_ctr_new[1]),
        .Q(p_0_in[1]));
endmodule

(* ORIG_REF_NAME = "aes_encipher_block" *) 
module switch_elements_aes_encipher_block
   (\round_ctr_reg_reg[1]_0 ,
    \round_ctr_reg_reg[1]_1 ,
    muxed_round_nr,
    \prev_key1_reg_reg[31] ,
    p_19_in,
    \prev_key1_reg_reg[0] ,
    \prev_key1_reg_reg[0]_0 ,
    \prev_key1_reg_reg[0]_1 ,
    \prev_key1_reg_reg[0]_2 ,
    \prev_key1_reg_reg[0]_3 ,
    \prev_key1_reg_reg[0]_4 ,
    \prev_key1_reg_reg[0]_5 ,
    \prev_key1_reg_reg[0]_6 ,
    \prev_key1_reg_reg[0]_7 ,
    \prev_key1_reg_reg[0]_8 ,
    \prev_key1_reg_reg[0]_9 ,
    \prev_key1_reg_reg[0]_10 ,
    \prev_key1_reg_reg[0]_11 ,
    \prev_key1_reg_reg[0]_12 ,
    \prev_key1_reg_reg[0]_13 ,
    \prev_key1_reg_reg[0]_14 ,
    \prev_key1_reg_reg[0]_15 ,
    \prev_key1_reg_reg[0]_16 ,
    \prev_key1_reg_reg[0]_17 ,
    \prev_key1_reg_reg[0]_18 ,
    \prev_key1_reg_reg[0]_19 ,
    \prev_key1_reg_reg[0]_20 ,
    \prev_key1_reg_reg[0]_21 ,
    \prev_key1_reg_reg[0]_22 ,
    \prev_key1_reg_reg[0]_23 ,
    \prev_key1_reg_reg[0]_24 ,
    \prev_key1_reg_reg[0]_25 ,
    \prev_key1_reg_reg[0]_26 ,
    \prev_key1_reg_reg[0]_27 ,
    \prev_key1_reg_reg[0]_28 ,
    \prev_key1_reg_reg[0]_29 ,
    \prev_key1_reg_reg[0]_30 ,
    \prev_key1_reg_reg[8] ,
    \prev_key1_reg_reg[8]_0 ,
    \prev_key1_reg_reg[8]_1 ,
    \prev_key1_reg_reg[8]_2 ,
    \prev_key1_reg_reg[8]_3 ,
    \prev_key1_reg_reg[8]_4 ,
    \prev_key1_reg_reg[8]_5 ,
    \prev_key1_reg_reg[8]_6 ,
    \prev_key1_reg_reg[8]_7 ,
    \prev_key1_reg_reg[8]_8 ,
    \prev_key1_reg_reg[8]_9 ,
    \prev_key1_reg_reg[8]_10 ,
    \prev_key1_reg_reg[8]_11 ,
    \prev_key1_reg_reg[8]_12 ,
    \prev_key1_reg_reg[8]_13 ,
    \prev_key1_reg_reg[8]_14 ,
    \prev_key1_reg_reg[8]_15 ,
    \prev_key1_reg_reg[8]_16 ,
    \prev_key1_reg_reg[8]_17 ,
    \prev_key1_reg_reg[8]_18 ,
    \prev_key1_reg_reg[8]_19 ,
    \prev_key1_reg_reg[8]_20 ,
    \prev_key1_reg_reg[8]_21 ,
    \prev_key1_reg_reg[8]_22 ,
    \prev_key1_reg_reg[8]_23 ,
    \prev_key1_reg_reg[8]_24 ,
    \prev_key1_reg_reg[8]_25 ,
    \prev_key1_reg_reg[8]_26 ,
    \prev_key1_reg_reg[8]_27 ,
    \prev_key1_reg_reg[8]_28 ,
    \prev_key1_reg_reg[8]_29 ,
    \prev_key1_reg_reg[8]_30 ,
    \prev_key1_reg_reg[16] ,
    \prev_key1_reg_reg[16]_0 ,
    \prev_key1_reg_reg[16]_1 ,
    \prev_key1_reg_reg[16]_2 ,
    \prev_key1_reg_reg[16]_3 ,
    \prev_key1_reg_reg[16]_4 ,
    \prev_key1_reg_reg[16]_5 ,
    \prev_key1_reg_reg[16]_6 ,
    \prev_key1_reg_reg[16]_7 ,
    \prev_key1_reg_reg[16]_8 ,
    \prev_key1_reg_reg[16]_9 ,
    \prev_key1_reg_reg[16]_10 ,
    \prev_key1_reg_reg[16]_11 ,
    \prev_key1_reg_reg[16]_12 ,
    \prev_key1_reg_reg[16]_13 ,
    \prev_key1_reg_reg[16]_14 ,
    \prev_key1_reg_reg[16]_15 ,
    \prev_key1_reg_reg[16]_16 ,
    \prev_key1_reg_reg[16]_17 ,
    \prev_key1_reg_reg[16]_18 ,
    \prev_key1_reg_reg[16]_19 ,
    \prev_key1_reg_reg[16]_20 ,
    \prev_key1_reg_reg[16]_21 ,
    \prev_key1_reg_reg[16]_22 ,
    \prev_key1_reg_reg[16]_23 ,
    \prev_key1_reg_reg[16]_24 ,
    \prev_key1_reg_reg[16]_25 ,
    \prev_key1_reg_reg[16]_26 ,
    \prev_key1_reg_reg[16]_27 ,
    \prev_key1_reg_reg[16]_28 ,
    \prev_key1_reg_reg[16]_29 ,
    \prev_key1_reg_reg[16]_30 ,
    \prev_key1_reg_reg[24] ,
    \prev_key1_reg_reg[24]_0 ,
    \prev_key1_reg_reg[24]_1 ,
    \prev_key1_reg_reg[24]_2 ,
    \prev_key1_reg_reg[24]_3 ,
    \prev_key1_reg_reg[24]_4 ,
    \prev_key1_reg_reg[24]_5 ,
    \prev_key1_reg_reg[24]_6 ,
    \prev_key1_reg_reg[24]_7 ,
    \prev_key1_reg_reg[24]_8 ,
    \prev_key1_reg_reg[24]_9 ,
    \prev_key1_reg_reg[24]_10 ,
    \prev_key1_reg_reg[24]_11 ,
    \prev_key1_reg_reg[24]_12 ,
    \prev_key1_reg_reg[24]_13 ,
    \prev_key1_reg_reg[24]_14 ,
    \prev_key1_reg_reg[24]_15 ,
    \prev_key1_reg_reg[24]_16 ,
    \prev_key1_reg_reg[24]_17 ,
    \prev_key1_reg_reg[24]_18 ,
    \prev_key1_reg_reg[24]_19 ,
    \prev_key1_reg_reg[24]_20 ,
    \prev_key1_reg_reg[24]_21 ,
    \prev_key1_reg_reg[24]_22 ,
    \prev_key1_reg_reg[24]_23 ,
    \prev_key1_reg_reg[24]_24 ,
    \prev_key1_reg_reg[24]_25 ,
    \prev_key1_reg_reg[24]_26 ,
    \prev_key1_reg_reg[24]_27 ,
    \prev_key1_reg_reg[24]_28 ,
    \prev_key1_reg_reg[24]_29 ,
    \prev_key1_reg_reg[24]_30 ,
    next_reg_reg,
    E,
    enc_ready,
    D,
    \round_ctr_reg_reg[3]_0 ,
    \round_ctr_reg_reg[3]_1 ,
    \round_ctr_reg_reg[1]_2 ,
    \round_ctr_reg_reg[1]_3 ,
    \round_ctr_reg_reg[1]_4 ,
    \round_ctr_reg_reg[0]_0 ,
    \round_ctr_reg_reg[0]_1 ,
    \round_ctr_reg_reg[0]_2 ,
    \round_ctr_reg_reg[0]_3 ,
    p_1_in,
    Q,
    init_state,
    round_key,
    new_sboxw,
    \prev_key1_reg[127]_i_5 ,
    result_valid_reg_reg,
    core_valid,
    core_block,
    p_0_out,
    addroundkey_return,
    key_ready,
    dec_ready,
    \block_w2_reg[28]_i_3 ,
    dec_new_block,
    clk_i,
    rst_i);
  output \round_ctr_reg_reg[1]_0 ;
  output \round_ctr_reg_reg[1]_1 ;
  output [3:0]muxed_round_nr;
  output [7:0]\prev_key1_reg_reg[31] ;
  output [7:0]p_19_in;
  output \prev_key1_reg_reg[0] ;
  output \prev_key1_reg_reg[0]_0 ;
  output \prev_key1_reg_reg[0]_1 ;
  output \prev_key1_reg_reg[0]_2 ;
  output \prev_key1_reg_reg[0]_3 ;
  output \prev_key1_reg_reg[0]_4 ;
  output \prev_key1_reg_reg[0]_5 ;
  output \prev_key1_reg_reg[0]_6 ;
  output \prev_key1_reg_reg[0]_7 ;
  output \prev_key1_reg_reg[0]_8 ;
  output \prev_key1_reg_reg[0]_9 ;
  output \prev_key1_reg_reg[0]_10 ;
  output \prev_key1_reg_reg[0]_11 ;
  output \prev_key1_reg_reg[0]_12 ;
  output \prev_key1_reg_reg[0]_13 ;
  output \prev_key1_reg_reg[0]_14 ;
  output \prev_key1_reg_reg[0]_15 ;
  output \prev_key1_reg_reg[0]_16 ;
  output \prev_key1_reg_reg[0]_17 ;
  output \prev_key1_reg_reg[0]_18 ;
  output \prev_key1_reg_reg[0]_19 ;
  output \prev_key1_reg_reg[0]_20 ;
  output \prev_key1_reg_reg[0]_21 ;
  output \prev_key1_reg_reg[0]_22 ;
  output \prev_key1_reg_reg[0]_23 ;
  output \prev_key1_reg_reg[0]_24 ;
  output \prev_key1_reg_reg[0]_25 ;
  output \prev_key1_reg_reg[0]_26 ;
  output \prev_key1_reg_reg[0]_27 ;
  output \prev_key1_reg_reg[0]_28 ;
  output \prev_key1_reg_reg[0]_29 ;
  output \prev_key1_reg_reg[0]_30 ;
  output \prev_key1_reg_reg[8] ;
  output \prev_key1_reg_reg[8]_0 ;
  output \prev_key1_reg_reg[8]_1 ;
  output \prev_key1_reg_reg[8]_2 ;
  output \prev_key1_reg_reg[8]_3 ;
  output \prev_key1_reg_reg[8]_4 ;
  output \prev_key1_reg_reg[8]_5 ;
  output \prev_key1_reg_reg[8]_6 ;
  output \prev_key1_reg_reg[8]_7 ;
  output \prev_key1_reg_reg[8]_8 ;
  output \prev_key1_reg_reg[8]_9 ;
  output \prev_key1_reg_reg[8]_10 ;
  output \prev_key1_reg_reg[8]_11 ;
  output \prev_key1_reg_reg[8]_12 ;
  output \prev_key1_reg_reg[8]_13 ;
  output \prev_key1_reg_reg[8]_14 ;
  output \prev_key1_reg_reg[8]_15 ;
  output \prev_key1_reg_reg[8]_16 ;
  output \prev_key1_reg_reg[8]_17 ;
  output \prev_key1_reg_reg[8]_18 ;
  output \prev_key1_reg_reg[8]_19 ;
  output \prev_key1_reg_reg[8]_20 ;
  output \prev_key1_reg_reg[8]_21 ;
  output \prev_key1_reg_reg[8]_22 ;
  output \prev_key1_reg_reg[8]_23 ;
  output \prev_key1_reg_reg[8]_24 ;
  output \prev_key1_reg_reg[8]_25 ;
  output \prev_key1_reg_reg[8]_26 ;
  output \prev_key1_reg_reg[8]_27 ;
  output \prev_key1_reg_reg[8]_28 ;
  output \prev_key1_reg_reg[8]_29 ;
  output \prev_key1_reg_reg[8]_30 ;
  output \prev_key1_reg_reg[16] ;
  output \prev_key1_reg_reg[16]_0 ;
  output \prev_key1_reg_reg[16]_1 ;
  output \prev_key1_reg_reg[16]_2 ;
  output \prev_key1_reg_reg[16]_3 ;
  output \prev_key1_reg_reg[16]_4 ;
  output \prev_key1_reg_reg[16]_5 ;
  output \prev_key1_reg_reg[16]_6 ;
  output \prev_key1_reg_reg[16]_7 ;
  output \prev_key1_reg_reg[16]_8 ;
  output \prev_key1_reg_reg[16]_9 ;
  output \prev_key1_reg_reg[16]_10 ;
  output \prev_key1_reg_reg[16]_11 ;
  output \prev_key1_reg_reg[16]_12 ;
  output \prev_key1_reg_reg[16]_13 ;
  output \prev_key1_reg_reg[16]_14 ;
  output \prev_key1_reg_reg[16]_15 ;
  output \prev_key1_reg_reg[16]_16 ;
  output \prev_key1_reg_reg[16]_17 ;
  output \prev_key1_reg_reg[16]_18 ;
  output \prev_key1_reg_reg[16]_19 ;
  output \prev_key1_reg_reg[16]_20 ;
  output \prev_key1_reg_reg[16]_21 ;
  output \prev_key1_reg_reg[16]_22 ;
  output \prev_key1_reg_reg[16]_23 ;
  output \prev_key1_reg_reg[16]_24 ;
  output \prev_key1_reg_reg[16]_25 ;
  output \prev_key1_reg_reg[16]_26 ;
  output \prev_key1_reg_reg[16]_27 ;
  output \prev_key1_reg_reg[16]_28 ;
  output \prev_key1_reg_reg[16]_29 ;
  output \prev_key1_reg_reg[16]_30 ;
  output \prev_key1_reg_reg[24] ;
  output \prev_key1_reg_reg[24]_0 ;
  output \prev_key1_reg_reg[24]_1 ;
  output \prev_key1_reg_reg[24]_2 ;
  output \prev_key1_reg_reg[24]_3 ;
  output \prev_key1_reg_reg[24]_4 ;
  output \prev_key1_reg_reg[24]_5 ;
  output \prev_key1_reg_reg[24]_6 ;
  output \prev_key1_reg_reg[24]_7 ;
  output \prev_key1_reg_reg[24]_8 ;
  output \prev_key1_reg_reg[24]_9 ;
  output \prev_key1_reg_reg[24]_10 ;
  output \prev_key1_reg_reg[24]_11 ;
  output \prev_key1_reg_reg[24]_12 ;
  output \prev_key1_reg_reg[24]_13 ;
  output \prev_key1_reg_reg[24]_14 ;
  output \prev_key1_reg_reg[24]_15 ;
  output \prev_key1_reg_reg[24]_16 ;
  output \prev_key1_reg_reg[24]_17 ;
  output \prev_key1_reg_reg[24]_18 ;
  output \prev_key1_reg_reg[24]_19 ;
  output \prev_key1_reg_reg[24]_20 ;
  output \prev_key1_reg_reg[24]_21 ;
  output \prev_key1_reg_reg[24]_22 ;
  output \prev_key1_reg_reg[24]_23 ;
  output \prev_key1_reg_reg[24]_24 ;
  output \prev_key1_reg_reg[24]_25 ;
  output \prev_key1_reg_reg[24]_26 ;
  output \prev_key1_reg_reg[24]_27 ;
  output \prev_key1_reg_reg[24]_28 ;
  output \prev_key1_reg_reg[24]_29 ;
  output \prev_key1_reg_reg[24]_30 ;
  output next_reg_reg;
  output [0:0]E;
  output enc_ready;
  output [127:0]D;
  output \round_ctr_reg_reg[3]_0 ;
  output \round_ctr_reg_reg[3]_1 ;
  output \round_ctr_reg_reg[1]_2 ;
  output \round_ctr_reg_reg[1]_3 ;
  output \round_ctr_reg_reg[1]_4 ;
  output \round_ctr_reg_reg[0]_0 ;
  output \round_ctr_reg_reg[0]_1 ;
  output \round_ctr_reg_reg[0]_2 ;
  output \round_ctr_reg_reg[0]_3 ;
  input [3:0]p_1_in;
  input [31:0]Q;
  input init_state;
  input [127:0]round_key;
  input [31:0]new_sboxw;
  input [7:0]\prev_key1_reg[127]_i_5 ;
  input [1:0]result_valid_reg_reg;
  input core_valid;
  input [79:0]core_block;
  input [29:0]p_0_out;
  input [17:0]addroundkey_return;
  input key_ready;
  input dec_ready;
  input [3:0]\block_w2_reg[28]_i_3 ;
  input [127:0]dec_new_block;
  input clk_i;
  input rst_i;

  wire [127:0]D;
  wire [0:0]E;
  wire \FSM_sequential_enc_ctrl_reg[1]_i_1_n_0 ;
  wire \FSM_sequential_enc_ctrl_reg[1]_i_3_n_0 ;
  wire [31:0]Q;
  wire [124:3]addroundkey0_return__514;
  wire [17:0]addroundkey_return;
  wire \block_w0_reg[0]_i_1__0_n_0 ;
  wire \block_w0_reg[0]_i_2_n_0 ;
  wire \block_w0_reg[10]_i_1_n_0 ;
  wire \block_w0_reg[10]_i_2_n_0 ;
  wire \block_w0_reg[11]_i_1_n_0 ;
  wire \block_w0_reg[11]_i_2_n_0 ;
  wire \block_w0_reg[12]_i_1_n_0 ;
  wire \block_w0_reg[12]_i_2_n_0 ;
  wire \block_w0_reg[13]_i_1_n_0 ;
  wire \block_w0_reg[13]_i_2_n_0 ;
  wire \block_w0_reg[14]_i_1_n_0 ;
  wire \block_w0_reg[14]_i_2_n_0 ;
  wire \block_w0_reg[15]_i_1_n_0 ;
  wire \block_w0_reg[15]_i_2_n_0 ;
  wire \block_w0_reg[16]_i_1__0_n_0 ;
  wire \block_w0_reg[16]_i_2_n_0 ;
  wire \block_w0_reg[17]_i_1_n_0 ;
  wire \block_w0_reg[17]_i_2_n_0 ;
  wire \block_w0_reg[17]_i_4_n_0 ;
  wire \block_w0_reg[18]_i_1_n_0 ;
  wire \block_w0_reg[18]_i_2_n_0 ;
  wire \block_w0_reg[19]_i_1_n_0 ;
  wire \block_w0_reg[19]_i_2_n_0 ;
  wire \block_w0_reg[1]_i_1_n_0 ;
  wire \block_w0_reg[1]_i_2_n_0 ;
  wire \block_w0_reg[1]_i_4_n_0 ;
  wire \block_w0_reg[20]_i_1_n_0 ;
  wire \block_w0_reg[20]_i_2_n_0 ;
  wire \block_w0_reg[20]_i_4__0_n_0 ;
  wire \block_w0_reg[20]_i_5_n_0 ;
  wire \block_w0_reg[21]_i_1_n_0 ;
  wire \block_w0_reg[21]_i_2_n_0 ;
  wire \block_w0_reg[22]_i_1_n_0 ;
  wire \block_w0_reg[22]_i_2_n_0 ;
  wire \block_w0_reg[23]_i_1_n_0 ;
  wire \block_w0_reg[23]_i_2_n_0 ;
  wire \block_w0_reg[24]_i_1_n_0 ;
  wire \block_w0_reg[24]_i_2_n_0 ;
  wire \block_w0_reg[25]_i_1_n_0 ;
  wire \block_w0_reg[25]_i_2_n_0 ;
  wire \block_w0_reg[25]_i_4__0_n_0 ;
  wire \block_w0_reg[25]_i_5__0_n_0 ;
  wire \block_w0_reg[26]_i_1_n_0 ;
  wire \block_w0_reg[26]_i_2_n_0 ;
  wire \block_w0_reg[27]_i_1_n_0 ;
  wire \block_w0_reg[27]_i_2_n_0 ;
  wire \block_w0_reg[27]_i_9_n_0 ;
  wire \block_w0_reg[28]_i_1_n_0 ;
  wire \block_w0_reg[28]_i_2_n_0 ;
  wire \block_w0_reg[28]_i_9_n_0 ;
  wire \block_w0_reg[29]_i_1_n_0 ;
  wire \block_w0_reg[29]_i_2_n_0 ;
  wire \block_w0_reg[2]_i_1_n_0 ;
  wire \block_w0_reg[2]_i_2_n_0 ;
  wire \block_w0_reg[30]_i_1_n_0 ;
  wire \block_w0_reg[30]_i_2_n_0 ;
  wire \block_w0_reg[31]_i_2_n_0 ;
  wire \block_w0_reg[31]_i_3_n_0 ;
  wire \block_w0_reg[3]_i_1_n_0 ;
  wire \block_w0_reg[3]_i_2_n_0 ;
  wire \block_w0_reg[4]_i_1_n_0 ;
  wire \block_w0_reg[4]_i_2_n_0 ;
  wire \block_w0_reg[4]_i_4__0_n_0 ;
  wire \block_w0_reg[4]_i_5_n_0 ;
  wire \block_w0_reg[5]_i_1_n_0 ;
  wire \block_w0_reg[5]_i_2_n_0 ;
  wire \block_w0_reg[6]_i_1_n_0 ;
  wire \block_w0_reg[6]_i_2_n_0 ;
  wire \block_w0_reg[7]_i_1_n_0 ;
  wire \block_w0_reg[7]_i_2_n_0 ;
  wire \block_w0_reg[8]_i_1_n_0 ;
  wire \block_w0_reg[8]_i_2_n_0 ;
  wire \block_w0_reg[9]_i_1_n_0 ;
  wire \block_w0_reg[9]_i_2_n_0 ;
  wire \block_w0_reg[9]_i_4__0_n_0 ;
  wire \block_w0_reg[9]_i_5_n_0 ;
  wire block_w0_we;
  wire \block_w1_reg[0]_i_1__0_n_0 ;
  wire \block_w1_reg[0]_i_2_n_0 ;
  wire \block_w1_reg[10]_i_1_n_0 ;
  wire \block_w1_reg[10]_i_2_n_0 ;
  wire \block_w1_reg[11]_i_1_n_0 ;
  wire \block_w1_reg[11]_i_2_n_0 ;
  wire \block_w1_reg[12]_i_1_n_0 ;
  wire \block_w1_reg[12]_i_2_n_0 ;
  wire \block_w1_reg[13]_i_1_n_0 ;
  wire \block_w1_reg[13]_i_2_n_0 ;
  wire \block_w1_reg[14]_i_1_n_0 ;
  wire \block_w1_reg[14]_i_2_n_0 ;
  wire \block_w1_reg[15]_i_1_n_0 ;
  wire \block_w1_reg[15]_i_2_n_0 ;
  wire \block_w1_reg[16]_i_1__0_n_0 ;
  wire \block_w1_reg[16]_i_2_n_0 ;
  wire \block_w1_reg[17]_i_1_n_0 ;
  wire \block_w1_reg[17]_i_2_n_0 ;
  wire \block_w1_reg[17]_i_4_n_0 ;
  wire \block_w1_reg[18]_i_1_n_0 ;
  wire \block_w1_reg[18]_i_2_n_0 ;
  wire \block_w1_reg[19]_i_1_n_0 ;
  wire \block_w1_reg[19]_i_2_n_0 ;
  wire \block_w1_reg[1]_i_1_n_0 ;
  wire \block_w1_reg[1]_i_2_n_0 ;
  wire \block_w1_reg[1]_i_4_n_0 ;
  wire \block_w1_reg[20]_i_1_n_0 ;
  wire \block_w1_reg[20]_i_2_n_0 ;
  wire \block_w1_reg[20]_i_4__0_n_0 ;
  wire \block_w1_reg[20]_i_5__0_n_0 ;
  wire \block_w1_reg[21]_i_1_n_0 ;
  wire \block_w1_reg[21]_i_2_n_0 ;
  wire \block_w1_reg[22]_i_1_n_0 ;
  wire \block_w1_reg[22]_i_2_n_0 ;
  wire \block_w1_reg[23]_i_1_n_0 ;
  wire \block_w1_reg[23]_i_2_n_0 ;
  wire \block_w1_reg[24]_i_1_n_0 ;
  wire \block_w1_reg[24]_i_2_n_0 ;
  wire \block_w1_reg[25]_i_1_n_0 ;
  wire \block_w1_reg[25]_i_2_n_0 ;
  wire \block_w1_reg[25]_i_4__0_n_0 ;
  wire \block_w1_reg[25]_i_5__0_n_0 ;
  wire \block_w1_reg[26]_i_1_n_0 ;
  wire \block_w1_reg[26]_i_2_n_0 ;
  wire \block_w1_reg[27]_i_1_n_0 ;
  wire \block_w1_reg[27]_i_2_n_0 ;
  wire \block_w1_reg[27]_i_9_n_0 ;
  wire \block_w1_reg[28]_i_1_n_0 ;
  wire \block_w1_reg[28]_i_2_n_0 ;
  wire \block_w1_reg[28]_i_9_n_0 ;
  wire \block_w1_reg[29]_i_1_n_0 ;
  wire \block_w1_reg[29]_i_2_n_0 ;
  wire \block_w1_reg[2]_i_1_n_0 ;
  wire \block_w1_reg[2]_i_2_n_0 ;
  wire \block_w1_reg[30]_i_1_n_0 ;
  wire \block_w1_reg[30]_i_2_n_0 ;
  wire \block_w1_reg[31]_i_2_n_0 ;
  wire \block_w1_reg[31]_i_3_n_0 ;
  wire \block_w1_reg[3]_i_1_n_0 ;
  wire \block_w1_reg[3]_i_2_n_0 ;
  wire \block_w1_reg[4]_i_1_n_0 ;
  wire \block_w1_reg[4]_i_2_n_0 ;
  wire \block_w1_reg[4]_i_4__0_n_0 ;
  wire \block_w1_reg[4]_i_5_n_0 ;
  wire \block_w1_reg[5]_i_1_n_0 ;
  wire \block_w1_reg[5]_i_2_n_0 ;
  wire \block_w1_reg[6]_i_1_n_0 ;
  wire \block_w1_reg[6]_i_2_n_0 ;
  wire \block_w1_reg[7]_i_1_n_0 ;
  wire \block_w1_reg[7]_i_2_n_0 ;
  wire \block_w1_reg[8]_i_1_n_0 ;
  wire \block_w1_reg[8]_i_2_n_0 ;
  wire \block_w1_reg[9]_i_1__0_n_0 ;
  wire \block_w1_reg[9]_i_2_n_0 ;
  wire \block_w1_reg[9]_i_4__0_n_0 ;
  wire \block_w1_reg[9]_i_5__0_n_0 ;
  wire block_w1_we;
  wire \block_w2_reg[0]_i_2_n_0 ;
  wire \block_w2_reg[10]_i_2_n_0 ;
  wire \block_w2_reg[11]_i_2_n_0 ;
  wire \block_w2_reg[12]_i_2_n_0 ;
  wire \block_w2_reg[13]_i_2_n_0 ;
  wire \block_w2_reg[14]_i_2_n_0 ;
  wire \block_w2_reg[15]_i_2_n_0 ;
  wire \block_w2_reg[16]_i_2_n_0 ;
  wire \block_w2_reg[17]_i_2_n_0 ;
  wire \block_w2_reg[17]_i_4_n_0 ;
  wire \block_w2_reg[18]_i_2_n_0 ;
  wire \block_w2_reg[19]_i_2_n_0 ;
  wire \block_w2_reg[1]_i_2_n_0 ;
  wire \block_w2_reg[1]_i_4_n_0 ;
  wire \block_w2_reg[20]_i_2_n_0 ;
  wire \block_w2_reg[20]_i_4__0_n_0 ;
  wire \block_w2_reg[20]_i_5__0_n_0 ;
  wire \block_w2_reg[21]_i_2_n_0 ;
  wire \block_w2_reg[22]_i_2_n_0 ;
  wire \block_w2_reg[23]_i_2_n_0 ;
  wire \block_w2_reg[24]_i_2_n_0 ;
  wire \block_w2_reg[25]_i_2_n_0 ;
  wire \block_w2_reg[25]_i_4__0_n_0 ;
  wire \block_w2_reg[25]_i_5__0_n_0 ;
  wire \block_w2_reg[26]_i_2_n_0 ;
  wire \block_w2_reg[27]_i_11_n_0 ;
  wire \block_w2_reg[27]_i_2_n_0 ;
  wire \block_w2_reg[28]_i_10_n_0 ;
  wire \block_w2_reg[28]_i_2_n_0 ;
  wire [3:0]\block_w2_reg[28]_i_3 ;
  wire \block_w2_reg[29]_i_2_n_0 ;
  wire \block_w2_reg[2]_i_2_n_0 ;
  wire \block_w2_reg[30]_i_2_n_0 ;
  wire \block_w2_reg[31]_i_6_n_0 ;
  wire \block_w2_reg[31]_i_8_n_0 ;
  wire \block_w2_reg[3]_i_2_n_0 ;
  wire \block_w2_reg[4]_i_2_n_0 ;
  wire \block_w2_reg[4]_i_4__0_n_0 ;
  wire \block_w2_reg[4]_i_5_n_0 ;
  wire \block_w2_reg[5]_i_2_n_0 ;
  wire \block_w2_reg[6]_i_2_n_0 ;
  wire \block_w2_reg[7]_i_2_n_0 ;
  wire \block_w2_reg[8]_i_2_n_0 ;
  wire \block_w2_reg[9]_i_2__0_n_0 ;
  wire \block_w2_reg[9]_i_4__0_n_0 ;
  wire \block_w2_reg[9]_i_5__0_n_0 ;
  wire block_w2_we;
  wire \block_w3_reg[0]_i_1__0_n_0 ;
  wire \block_w3_reg[0]_i_2_n_0 ;
  wire \block_w3_reg[10]_i_1_n_0 ;
  wire \block_w3_reg[10]_i_2_n_0 ;
  wire \block_w3_reg[11]_i_1_n_0 ;
  wire \block_w3_reg[11]_i_2_n_0 ;
  wire \block_w3_reg[12]_i_1_n_0 ;
  wire \block_w3_reg[12]_i_2_n_0 ;
  wire \block_w3_reg[13]_i_1_n_0 ;
  wire \block_w3_reg[13]_i_2_n_0 ;
  wire \block_w3_reg[14]_i_1_n_0 ;
  wire \block_w3_reg[14]_i_2_n_0 ;
  wire \block_w3_reg[15]_i_1_n_0 ;
  wire \block_w3_reg[15]_i_2_n_0 ;
  wire \block_w3_reg[16]_i_1__0_n_0 ;
  wire \block_w3_reg[16]_i_2_n_0 ;
  wire \block_w3_reg[17]_i_1_n_0 ;
  wire \block_w3_reg[17]_i_2_n_0 ;
  wire \block_w3_reg[17]_i_4_n_0 ;
  wire \block_w3_reg[18]_i_1_n_0 ;
  wire \block_w3_reg[18]_i_2_n_0 ;
  wire \block_w3_reg[19]_i_1_n_0 ;
  wire \block_w3_reg[19]_i_2_n_0 ;
  wire \block_w3_reg[19]_i_9__0_n_0 ;
  wire \block_w3_reg[1]_i_1_n_0 ;
  wire \block_w3_reg[1]_i_2_n_0 ;
  wire \block_w3_reg[1]_i_4_n_0 ;
  wire \block_w3_reg[20]_i_1_n_0 ;
  wire \block_w3_reg[20]_i_2_n_0 ;
  wire \block_w3_reg[20]_i_4__0_n_0 ;
  wire \block_w3_reg[20]_i_5_n_0 ;
  wire \block_w3_reg[21]_i_1_n_0 ;
  wire \block_w3_reg[21]_i_2_n_0 ;
  wire \block_w3_reg[22]_i_1_n_0 ;
  wire \block_w3_reg[22]_i_2_n_0 ;
  wire \block_w3_reg[23]_i_1_n_0 ;
  wire \block_w3_reg[23]_i_2_n_0 ;
  wire \block_w3_reg[24]_i_1_n_0 ;
  wire \block_w3_reg[24]_i_2_n_0 ;
  wire \block_w3_reg[25]_i_1_n_0 ;
  wire \block_w3_reg[25]_i_2_n_0 ;
  wire \block_w3_reg[25]_i_4__0_n_0 ;
  wire \block_w3_reg[25]_i_5_n_0 ;
  wire \block_w3_reg[26]_i_1_n_0 ;
  wire \block_w3_reg[26]_i_2_n_0 ;
  wire \block_w3_reg[27]_i_1_n_0 ;
  wire \block_w3_reg[27]_i_2_n_0 ;
  wire \block_w3_reg[27]_i_9__0_n_0 ;
  wire \block_w3_reg[28]_i_1_n_0 ;
  wire \block_w3_reg[28]_i_2_n_0 ;
  wire \block_w3_reg[28]_i_9__0_n_0 ;
  wire \block_w3_reg[29]_i_1_n_0 ;
  wire \block_w3_reg[29]_i_2_n_0 ;
  wire \block_w3_reg[2]_i_1_n_0 ;
  wire \block_w3_reg[2]_i_2_n_0 ;
  wire \block_w3_reg[30]_i_1_n_0 ;
  wire \block_w3_reg[30]_i_2_n_0 ;
  wire \block_w3_reg[31]_i_2_n_0 ;
  wire \block_w3_reg[31]_i_3_n_0 ;
  wire \block_w3_reg[3]_i_1_n_0 ;
  wire \block_w3_reg[3]_i_2_n_0 ;
  wire \block_w3_reg[4]_i_1_n_0 ;
  wire \block_w3_reg[4]_i_2_n_0 ;
  wire \block_w3_reg[4]_i_4__0_n_0 ;
  wire \block_w3_reg[4]_i_5_n_0 ;
  wire \block_w3_reg[5]_i_1_n_0 ;
  wire \block_w3_reg[5]_i_2_n_0 ;
  wire \block_w3_reg[6]_i_1_n_0 ;
  wire \block_w3_reg[6]_i_2_n_0 ;
  wire \block_w3_reg[7]_i_1_n_0 ;
  wire \block_w3_reg[7]_i_2_n_0 ;
  wire \block_w3_reg[8]_i_1_n_0 ;
  wire \block_w3_reg[8]_i_2_n_0 ;
  wire \block_w3_reg[9]_i_1_n_0 ;
  wire \block_w3_reg[9]_i_2_n_0 ;
  wire \block_w3_reg[9]_i_4__0_n_0 ;
  wire \block_w3_reg[9]_i_5_n_0 ;
  wire block_w3_we;
  wire clk_i;
  wire [79:0]core_block;
  wire core_valid;
  wire [127:0]dec_new_block;
  wire dec_ready;
  wire [1:0]enc_ctrl_new;
  wire [1:1]enc_ctrl_reg;
  wire [127:0]enc_new_block;
  wire enc_ready;
  wire [3:0]enc_round_nr;
  wire init_state;
  wire key_ready;
  wire [7:0]mixcolumns_return0;
  wire [7:0]mixcolumns_return022_out;
  wire [7:0]mixcolumns_return025_out;
  wire [7:0]mixcolumns_return028_out;
  wire [7:0]mixcolumns_return034_out;
  wire [7:0]mixcolumns_return038_out;
  wire [7:0]mixcolumns_return041_out;
  wire [7:0]mixcolumns_return044_out;
  wire [7:0]mixcolumns_return050_out;
  wire [7:0]mixcolumns_return054_out;
  wire [7:0]mixcolumns_return057_out;
  wire [7:0]mixcolumns_return060_out;
  wire [7:0]mixcolumns_return066_out;
  wire [7:0]mixcolumns_return070_out;
  wire [7:0]mixcolumns_return073_out;
  wire [7:0]mixcolumns_return076_out;
  wire muxed_ready;
  wire [3:0]muxed_round_nr;
  wire [29:0]muxed_sboxw;
  wire [31:0]muxed_sboxw__0;
  wire [31:0]new_sboxw;
  wire next_reg_reg;
  wire [1:0]p_0_in;
  wire [31:0]p_0_in__0;
  wire [29:0]p_0_out;
  wire [7:0]p_19_in;
  wire [3:0]p_1_in;
  wire [7:0]\prev_key1_reg[127]_i_5 ;
  wire \prev_key1_reg_reg[0] ;
  wire \prev_key1_reg_reg[0]_0 ;
  wire \prev_key1_reg_reg[0]_1 ;
  wire \prev_key1_reg_reg[0]_10 ;
  wire \prev_key1_reg_reg[0]_11 ;
  wire \prev_key1_reg_reg[0]_12 ;
  wire \prev_key1_reg_reg[0]_13 ;
  wire \prev_key1_reg_reg[0]_14 ;
  wire \prev_key1_reg_reg[0]_15 ;
  wire \prev_key1_reg_reg[0]_16 ;
  wire \prev_key1_reg_reg[0]_17 ;
  wire \prev_key1_reg_reg[0]_18 ;
  wire \prev_key1_reg_reg[0]_19 ;
  wire \prev_key1_reg_reg[0]_2 ;
  wire \prev_key1_reg_reg[0]_20 ;
  wire \prev_key1_reg_reg[0]_21 ;
  wire \prev_key1_reg_reg[0]_22 ;
  wire \prev_key1_reg_reg[0]_23 ;
  wire \prev_key1_reg_reg[0]_24 ;
  wire \prev_key1_reg_reg[0]_25 ;
  wire \prev_key1_reg_reg[0]_26 ;
  wire \prev_key1_reg_reg[0]_27 ;
  wire \prev_key1_reg_reg[0]_28 ;
  wire \prev_key1_reg_reg[0]_29 ;
  wire \prev_key1_reg_reg[0]_3 ;
  wire \prev_key1_reg_reg[0]_30 ;
  wire \prev_key1_reg_reg[0]_4 ;
  wire \prev_key1_reg_reg[0]_5 ;
  wire \prev_key1_reg_reg[0]_6 ;
  wire \prev_key1_reg_reg[0]_7 ;
  wire \prev_key1_reg_reg[0]_8 ;
  wire \prev_key1_reg_reg[0]_9 ;
  wire \prev_key1_reg_reg[16] ;
  wire \prev_key1_reg_reg[16]_0 ;
  wire \prev_key1_reg_reg[16]_1 ;
  wire \prev_key1_reg_reg[16]_10 ;
  wire \prev_key1_reg_reg[16]_11 ;
  wire \prev_key1_reg_reg[16]_12 ;
  wire \prev_key1_reg_reg[16]_13 ;
  wire \prev_key1_reg_reg[16]_14 ;
  wire \prev_key1_reg_reg[16]_15 ;
  wire \prev_key1_reg_reg[16]_16 ;
  wire \prev_key1_reg_reg[16]_17 ;
  wire \prev_key1_reg_reg[16]_18 ;
  wire \prev_key1_reg_reg[16]_19 ;
  wire \prev_key1_reg_reg[16]_2 ;
  wire \prev_key1_reg_reg[16]_20 ;
  wire \prev_key1_reg_reg[16]_21 ;
  wire \prev_key1_reg_reg[16]_22 ;
  wire \prev_key1_reg_reg[16]_23 ;
  wire \prev_key1_reg_reg[16]_24 ;
  wire \prev_key1_reg_reg[16]_25 ;
  wire \prev_key1_reg_reg[16]_26 ;
  wire \prev_key1_reg_reg[16]_27 ;
  wire \prev_key1_reg_reg[16]_28 ;
  wire \prev_key1_reg_reg[16]_29 ;
  wire \prev_key1_reg_reg[16]_3 ;
  wire \prev_key1_reg_reg[16]_30 ;
  wire \prev_key1_reg_reg[16]_4 ;
  wire \prev_key1_reg_reg[16]_5 ;
  wire \prev_key1_reg_reg[16]_6 ;
  wire \prev_key1_reg_reg[16]_7 ;
  wire \prev_key1_reg_reg[16]_8 ;
  wire \prev_key1_reg_reg[16]_9 ;
  wire \prev_key1_reg_reg[24] ;
  wire \prev_key1_reg_reg[24]_0 ;
  wire \prev_key1_reg_reg[24]_1 ;
  wire \prev_key1_reg_reg[24]_10 ;
  wire \prev_key1_reg_reg[24]_11 ;
  wire \prev_key1_reg_reg[24]_12 ;
  wire \prev_key1_reg_reg[24]_13 ;
  wire \prev_key1_reg_reg[24]_14 ;
  wire \prev_key1_reg_reg[24]_15 ;
  wire \prev_key1_reg_reg[24]_16 ;
  wire \prev_key1_reg_reg[24]_17 ;
  wire \prev_key1_reg_reg[24]_18 ;
  wire \prev_key1_reg_reg[24]_19 ;
  wire \prev_key1_reg_reg[24]_2 ;
  wire \prev_key1_reg_reg[24]_20 ;
  wire \prev_key1_reg_reg[24]_21 ;
  wire \prev_key1_reg_reg[24]_22 ;
  wire \prev_key1_reg_reg[24]_23 ;
  wire \prev_key1_reg_reg[24]_24 ;
  wire \prev_key1_reg_reg[24]_25 ;
  wire \prev_key1_reg_reg[24]_26 ;
  wire \prev_key1_reg_reg[24]_27 ;
  wire \prev_key1_reg_reg[24]_28 ;
  wire \prev_key1_reg_reg[24]_29 ;
  wire \prev_key1_reg_reg[24]_3 ;
  wire \prev_key1_reg_reg[24]_30 ;
  wire \prev_key1_reg_reg[24]_4 ;
  wire \prev_key1_reg_reg[24]_5 ;
  wire \prev_key1_reg_reg[24]_6 ;
  wire \prev_key1_reg_reg[24]_7 ;
  wire \prev_key1_reg_reg[24]_8 ;
  wire \prev_key1_reg_reg[24]_9 ;
  wire [7:0]\prev_key1_reg_reg[31] ;
  wire \prev_key1_reg_reg[8] ;
  wire \prev_key1_reg_reg[8]_0 ;
  wire \prev_key1_reg_reg[8]_1 ;
  wire \prev_key1_reg_reg[8]_10 ;
  wire \prev_key1_reg_reg[8]_11 ;
  wire \prev_key1_reg_reg[8]_12 ;
  wire \prev_key1_reg_reg[8]_13 ;
  wire \prev_key1_reg_reg[8]_14 ;
  wire \prev_key1_reg_reg[8]_15 ;
  wire \prev_key1_reg_reg[8]_16 ;
  wire \prev_key1_reg_reg[8]_17 ;
  wire \prev_key1_reg_reg[8]_18 ;
  wire \prev_key1_reg_reg[8]_19 ;
  wire \prev_key1_reg_reg[8]_2 ;
  wire \prev_key1_reg_reg[8]_20 ;
  wire \prev_key1_reg_reg[8]_21 ;
  wire \prev_key1_reg_reg[8]_22 ;
  wire \prev_key1_reg_reg[8]_23 ;
  wire \prev_key1_reg_reg[8]_24 ;
  wire \prev_key1_reg_reg[8]_25 ;
  wire \prev_key1_reg_reg[8]_26 ;
  wire \prev_key1_reg_reg[8]_27 ;
  wire \prev_key1_reg_reg[8]_28 ;
  wire \prev_key1_reg_reg[8]_29 ;
  wire \prev_key1_reg_reg[8]_3 ;
  wire \prev_key1_reg_reg[8]_30 ;
  wire \prev_key1_reg_reg[8]_4 ;
  wire \prev_key1_reg_reg[8]_5 ;
  wire \prev_key1_reg_reg[8]_6 ;
  wire \prev_key1_reg_reg[8]_7 ;
  wire \prev_key1_reg_reg[8]_8 ;
  wire \prev_key1_reg_reg[8]_9 ;
  wire ready_new;
  wire ready_reg_i_1_n_0;
  wire ready_reg_i_2__0_n_0;
  wire [1:0]result_valid_reg_reg;
  wire round_ctr_inc;
  wire [3:0]round_ctr_new;
  wire \round_ctr_reg_reg[0]_0 ;
  wire \round_ctr_reg_reg[0]_1 ;
  wire \round_ctr_reg_reg[0]_2 ;
  wire \round_ctr_reg_reg[0]_3 ;
  wire \round_ctr_reg_reg[1]_0 ;
  wire \round_ctr_reg_reg[1]_1 ;
  wire \round_ctr_reg_reg[1]_2 ;
  wire \round_ctr_reg_reg[1]_3 ;
  wire \round_ctr_reg_reg[1]_4 ;
  wire \round_ctr_reg_reg[3]_0 ;
  wire \round_ctr_reg_reg[3]_1 ;
  wire round_ctr_rst__1;
  wire round_ctr_we;
  wire [127:0]round_key;
  wire rst_i;
  wire [1:0]sword_ctr_new;
  wire sword_ctr_we;
  wire [1:0]update_type__0;

  LUT6 #(
    .INIT(64'h00F0FFEE00F000EE)) 
    \FSM_sequential_aes_core_ctrl_reg[1]_i_1 
       (.I0(p_1_in[0]),
        .I1(p_1_in[1]),
        .I2(muxed_ready),
        .I3(result_valid_reg_reg[0]),
        .I4(result_valid_reg_reg[1]),
        .I5(key_ready),
        .O(E));
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \FSM_sequential_aes_core_ctrl_reg[1]_i_3 
       (.I0(enc_ready),
        .I1(p_1_in[2]),
        .I2(dec_ready),
        .O(muxed_ready));
  LUT6 #(
    .INIT(64'h00000000F8080808)) 
    \FSM_sequential_enc_ctrl_reg[0]_i_1 
       (.I0(p_1_in[1]),
        .I1(p_1_in[2]),
        .I2(enc_ctrl_reg),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(round_ctr_inc),
        .O(enc_ctrl_new[0]));
  LUT6 #(
    .INIT(64'hFFEAAAEAAAEAAAEA)) 
    \FSM_sequential_enc_ctrl_reg[1]_i_1 
       (.I0(round_ctr_inc),
        .I1(p_1_in[1]),
        .I2(p_1_in[2]),
        .I3(enc_ctrl_reg),
        .I4(p_0_in[1]),
        .I5(p_0_in[0]),
        .O(\FSM_sequential_enc_ctrl_reg[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT5 #(
    .INIT(32'hB8888888)) 
    \FSM_sequential_enc_ctrl_reg[1]_i_2 
       (.I0(\FSM_sequential_enc_ctrl_reg[1]_i_3_n_0 ),
        .I1(round_ctr_inc),
        .I2(p_0_in[1]),
        .I3(p_0_in[0]),
        .I4(enc_ctrl_reg),
        .O(enc_ctrl_new[1]));
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT5 #(
    .INIT(32'h5DDFFFFF)) 
    \FSM_sequential_enc_ctrl_reg[1]_i_3 
       (.I0(enc_round_nr[3]),
        .I1(p_1_in[3]),
        .I2(enc_round_nr[2]),
        .I3(enc_round_nr[1]),
        .I4(enc_ctrl_reg),
        .O(\FSM_sequential_enc_ctrl_reg[1]_i_3_n_0 ));
  (* FSM_ENCODED_STATES = "CTRL_INIT:01,CTRL_MAIN:11,CTRL_IDLE:00,CTRL_SBOX:10" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_enc_ctrl_reg_reg[0] 
       (.C(clk_i),
        .CE(\FSM_sequential_enc_ctrl_reg[1]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enc_ctrl_new[0]),
        .Q(round_ctr_inc));
  (* FSM_ENCODED_STATES = "CTRL_INIT:01,CTRL_MAIN:11,CTRL_IDLE:00,CTRL_SBOX:10" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_enc_ctrl_reg_reg[1] 
       (.C(clk_i),
        .CE(\FSM_sequential_enc_ctrl_reg[1]_i_1_n_0 ),
        .CLR(rst_i),
        .D(enc_ctrl_new[1]),
        .Q(enc_ctrl_reg));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[0]_i_1__0 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[0]_i_2_n_0 ),
        .I3(enc_new_block[0]),
        .I4(round_key[96]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[0]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[0]_i_2 
       (.I0(mixcolumns_return066_out[0]),
        .I1(new_sboxw[0]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[60]),
        .I5(round_key[96]),
        .O(\block_w0_reg[0]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[0]_i_4__0 
       (.I0(enc_new_block[80]),
        .I1(enc_new_block[7]),
        .I2(enc_new_block[127]),
        .I3(enc_new_block[40]),
        .I4(enc_new_block[120]),
        .O(mixcolumns_return066_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[10]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[10]_i_2_n_0 ),
        .I3(enc_new_block[42]),
        .I4(round_key[106]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[10]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[10]_i_2 
       (.I0(mixcolumns_return070_out[2]),
        .I1(new_sboxw[10]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[66]),
        .I5(round_key[106]),
        .O(\block_w0_reg[10]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[10]_i_4__0 
       (.I0(enc_new_block[82]),
        .I1(enc_new_block[1]),
        .I2(enc_new_block[41]),
        .I3(enc_new_block[2]),
        .I4(enc_new_block[122]),
        .O(mixcolumns_return070_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[11]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[11]_i_2_n_0 ),
        .I3(enc_new_block[43]),
        .I4(round_key[107]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[11]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w0_reg[11]_i_2 
       (.I0(addroundkey0_return__514[107]),
        .I1(new_sboxw[11]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[22]),
        .O(\block_w0_reg[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[11]_i_4 
       (.I0(\block_w0_reg[28]_i_9_n_0 ),
        .I1(\block_w0_reg[9]_i_4__0_n_0 ),
        .I2(enc_new_block[2]),
        .I3(round_key[107]),
        .I4(enc_new_block[42]),
        .I5(enc_new_block[3]),
        .O(addroundkey0_return__514[107]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[12]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[12]_i_2_n_0 ),
        .I3(enc_new_block[44]),
        .I4(round_key[108]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[12]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w0_reg[12]_i_2 
       (.I0(addroundkey0_return__514[108]),
        .I1(new_sboxw[12]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[23]),
        .O(\block_w0_reg[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[12]_i_4 
       (.I0(\block_w0_reg[27]_i_9_n_0 ),
        .I1(\block_w0_reg[9]_i_4__0_n_0 ),
        .I2(enc_new_block[124]),
        .I3(round_key[108]),
        .I4(enc_new_block[4]),
        .I5(enc_new_block[84]),
        .O(addroundkey0_return__514[108]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[13]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[13]_i_2_n_0 ),
        .I3(enc_new_block[45]),
        .I4(round_key[109]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[13]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[13]_i_2 
       (.I0(mixcolumns_return070_out[5]),
        .I1(new_sboxw[13]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[67]),
        .I5(round_key[109]),
        .O(\block_w0_reg[13]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[13]_i_4__0 
       (.I0(enc_new_block[85]),
        .I1(enc_new_block[4]),
        .I2(enc_new_block[44]),
        .I3(enc_new_block[5]),
        .I4(enc_new_block[125]),
        .O(mixcolumns_return070_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[14]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[14]_i_2_n_0 ),
        .I3(enc_new_block[46]),
        .I4(round_key[110]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[14]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[14]_i_2 
       (.I0(mixcolumns_return070_out[6]),
        .I1(new_sboxw[14]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[68]),
        .I5(round_key[110]),
        .O(\block_w0_reg[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[14]_i_4__0 
       (.I0(enc_new_block[86]),
        .I1(enc_new_block[5]),
        .I2(enc_new_block[45]),
        .I3(enc_new_block[6]),
        .I4(enc_new_block[126]),
        .O(mixcolumns_return070_out[6]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[15]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[15]_i_2_n_0 ),
        .I3(enc_new_block[47]),
        .I4(round_key[111]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[15]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[15]_i_2 
       (.I0(mixcolumns_return070_out[7]),
        .I1(new_sboxw[15]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[69]),
        .I5(round_key[111]),
        .O(\block_w0_reg[15]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[15]_i_4__0 
       (.I0(enc_new_block[87]),
        .I1(enc_new_block[6]),
        .I2(enc_new_block[46]),
        .I3(enc_new_block[7]),
        .I4(enc_new_block[127]),
        .O(mixcolumns_return070_out[7]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[16]_i_1__0 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[16]_i_2_n_0 ),
        .I3(enc_new_block[80]),
        .I4(round_key[112]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[16]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[16]_i_2 
       (.I0(mixcolumns_return073_out[0]),
        .I1(new_sboxw[16]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[70]),
        .I5(round_key[112]),
        .O(\block_w0_reg[16]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[16]_i_4__0 
       (.I0(enc_new_block[120]),
        .I1(enc_new_block[87]),
        .I2(enc_new_block[0]),
        .I3(enc_new_block[40]),
        .I4(enc_new_block[47]),
        .O(mixcolumns_return073_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[17]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[17]_i_2_n_0 ),
        .I3(enc_new_block[81]),
        .I4(round_key[113]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[17]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w0_reg[17]_i_2 
       (.I0(\block_w0_reg[20]_i_4__0_n_0 ),
        .I1(\block_w0_reg[17]_i_4_n_0 ),
        .I2(new_sboxw[17]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[24]),
        .O(\block_w0_reg[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[17]_i_4 
       (.I0(enc_new_block[1]),
        .I1(enc_new_block[80]),
        .I2(enc_new_block[121]),
        .I3(round_key[113]),
        .I4(enc_new_block[40]),
        .I5(enc_new_block[41]),
        .O(\block_w0_reg[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[18]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[18]_i_2_n_0 ),
        .I3(enc_new_block[82]),
        .I4(round_key[114]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[18]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[18]_i_2 
       (.I0(mixcolumns_return073_out[2]),
        .I1(new_sboxw[18]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[71]),
        .I5(round_key[114]),
        .O(\block_w0_reg[18]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[18]_i_4__0 
       (.I0(enc_new_block[122]),
        .I1(enc_new_block[81]),
        .I2(enc_new_block[2]),
        .I3(enc_new_block[42]),
        .I4(enc_new_block[41]),
        .O(mixcolumns_return073_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[19]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[19]_i_2_n_0 ),
        .I3(enc_new_block[83]),
        .I4(round_key[115]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[19]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w0_reg[19]_i_2 
       (.I0(addroundkey0_return__514[115]),
        .I1(new_sboxw[19]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[25]),
        .O(\block_w0_reg[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[19]_i_4 
       (.I0(\block_w0_reg[20]_i_4__0_n_0 ),
        .I1(\block_w0_reg[27]_i_9_n_0 ),
        .I2(enc_new_block[123]),
        .I3(round_key[115]),
        .I4(enc_new_block[82]),
        .I5(enc_new_block[42]),
        .O(addroundkey0_return__514[115]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[1]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[1]_i_2_n_0 ),
        .I3(enc_new_block[1]),
        .I4(round_key[97]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w0_reg[1]_i_2 
       (.I0(\block_w0_reg[4]_i_4__0_n_0 ),
        .I1(\block_w0_reg[1]_i_4_n_0 ),
        .I2(new_sboxw[1]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[18]),
        .O(\block_w0_reg[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[1]_i_4 
       (.I0(enc_new_block[41]),
        .I1(enc_new_block[81]),
        .I2(enc_new_block[120]),
        .I3(round_key[97]),
        .I4(enc_new_block[121]),
        .I5(enc_new_block[0]),
        .O(\block_w0_reg[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[20]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[20]_i_2_n_0 ),
        .I3(enc_new_block[84]),
        .I4(round_key[116]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[20]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w0_reg[20]_i_2 
       (.I0(\block_w0_reg[20]_i_4__0_n_0 ),
        .I1(\block_w0_reg[20]_i_5_n_0 ),
        .I2(new_sboxw[20]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[26]),
        .O(\block_w0_reg[20]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[20]_i_4__0 
       (.I0(enc_new_block[87]),
        .I1(enc_new_block[47]),
        .O(\block_w0_reg[20]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[20]_i_5 
       (.I0(enc_new_block[44]),
        .I1(enc_new_block[4]),
        .I2(enc_new_block[43]),
        .I3(round_key[116]),
        .I4(enc_new_block[124]),
        .I5(enc_new_block[83]),
        .O(\block_w0_reg[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[21]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[21]_i_2_n_0 ),
        .I3(enc_new_block[85]),
        .I4(round_key[117]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[21]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[21]_i_2 
       (.I0(mixcolumns_return073_out[5]),
        .I1(new_sboxw[21]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[72]),
        .I5(round_key[117]),
        .O(\block_w0_reg[21]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[21]_i_4__0 
       (.I0(enc_new_block[125]),
        .I1(enc_new_block[84]),
        .I2(enc_new_block[5]),
        .I3(enc_new_block[45]),
        .I4(enc_new_block[44]),
        .O(mixcolumns_return073_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[22]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[22]_i_2_n_0 ),
        .I3(enc_new_block[86]),
        .I4(round_key[118]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[22]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[22]_i_2 
       (.I0(mixcolumns_return073_out[6]),
        .I1(new_sboxw[22]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[73]),
        .I5(round_key[118]),
        .O(\block_w0_reg[22]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[22]_i_4__0 
       (.I0(enc_new_block[126]),
        .I1(enc_new_block[85]),
        .I2(enc_new_block[6]),
        .I3(enc_new_block[46]),
        .I4(enc_new_block[45]),
        .O(mixcolumns_return073_out[6]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[23]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[23]_i_2_n_0 ),
        .I3(enc_new_block[87]),
        .I4(round_key[119]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[23]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[23]_i_2 
       (.I0(mixcolumns_return073_out[7]),
        .I1(new_sboxw[23]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[74]),
        .I5(round_key[119]),
        .O(\block_w0_reg[23]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[23]_i_4__0 
       (.I0(enc_new_block[127]),
        .I1(enc_new_block[86]),
        .I2(enc_new_block[7]),
        .I3(enc_new_block[47]),
        .I4(enc_new_block[46]),
        .O(mixcolumns_return073_out[7]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[24]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[24]_i_2_n_0 ),
        .I3(enc_new_block[120]),
        .I4(round_key[120]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[24]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[24]_i_2 
       (.I0(mixcolumns_return076_out[0]),
        .I1(new_sboxw[24]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[75]),
        .I5(round_key[120]),
        .O(\block_w0_reg[24]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[24]_i_4__0 
       (.I0(enc_new_block[127]),
        .I1(enc_new_block[87]),
        .I2(enc_new_block[0]),
        .I3(enc_new_block[40]),
        .I4(enc_new_block[80]),
        .O(mixcolumns_return076_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[25]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[25]_i_2_n_0 ),
        .I3(enc_new_block[121]),
        .I4(round_key[121]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[25]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w0_reg[25]_i_2 
       (.I0(\block_w0_reg[25]_i_4__0_n_0 ),
        .I1(\block_w0_reg[25]_i_5__0_n_0 ),
        .I2(new_sboxw[25]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[27]),
        .O(\block_w0_reg[25]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[25]_i_4__0 
       (.I0(enc_new_block[87]),
        .I1(enc_new_block[127]),
        .O(\block_w0_reg[25]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[25]_i_5__0 
       (.I0(enc_new_block[1]),
        .I1(enc_new_block[80]),
        .I2(enc_new_block[120]),
        .I3(round_key[121]),
        .I4(enc_new_block[81]),
        .I5(enc_new_block[41]),
        .O(\block_w0_reg[25]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[26]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[26]_i_2_n_0 ),
        .I3(enc_new_block[122]),
        .I4(round_key[122]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[26]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[26]_i_2 
       (.I0(mixcolumns_return076_out[2]),
        .I1(new_sboxw[26]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[76]),
        .I5(round_key[122]),
        .O(\block_w0_reg[26]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[26]_i_4__0 
       (.I0(enc_new_block[121]),
        .I1(enc_new_block[81]),
        .I2(enc_new_block[2]),
        .I3(enc_new_block[42]),
        .I4(enc_new_block[82]),
        .O(mixcolumns_return076_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[27]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[27]_i_2_n_0 ),
        .I3(enc_new_block[123]),
        .I4(round_key[123]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[27]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w0_reg[27]_i_2 
       (.I0(addroundkey0_return__514[123]),
        .I1(new_sboxw[27]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[28]),
        .O(\block_w0_reg[27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[27]_i_4__0 
       (.I0(\block_w0_reg[27]_i_9_n_0 ),
        .I1(\block_w0_reg[25]_i_4__0_n_0 ),
        .I2(enc_new_block[122]),
        .I3(round_key[123]),
        .I4(enc_new_block[82]),
        .I5(enc_new_block[83]),
        .O(addroundkey0_return__514[123]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[27]_i_9 
       (.I0(enc_new_block[3]),
        .I1(enc_new_block[43]),
        .O(\block_w0_reg[27]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[28]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[28]_i_2_n_0 ),
        .I3(enc_new_block[124]),
        .I4(round_key[124]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[28]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w0_reg[28]_i_2 
       (.I0(addroundkey0_return__514[124]),
        .I1(new_sboxw[28]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[29]),
        .O(\block_w0_reg[28]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[28]_i_4 
       (.I0(\block_w0_reg[28]_i_9_n_0 ),
        .I1(\block_w0_reg[25]_i_4__0_n_0 ),
        .I2(enc_new_block[44]),
        .I3(round_key[124]),
        .I4(enc_new_block[4]),
        .I5(enc_new_block[84]),
        .O(addroundkey0_return__514[124]));
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[28]_i_9 
       (.I0(enc_new_block[83]),
        .I1(enc_new_block[123]),
        .O(\block_w0_reg[28]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[29]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[29]_i_2_n_0 ),
        .I3(enc_new_block[125]),
        .I4(round_key[125]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[29]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[29]_i_2 
       (.I0(mixcolumns_return076_out[5]),
        .I1(new_sboxw[29]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[77]),
        .I5(round_key[125]),
        .O(\block_w0_reg[29]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[29]_i_4__0 
       (.I0(enc_new_block[124]),
        .I1(enc_new_block[84]),
        .I2(enc_new_block[5]),
        .I3(enc_new_block[45]),
        .I4(enc_new_block[85]),
        .O(mixcolumns_return076_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[2]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[2]_i_2_n_0 ),
        .I3(enc_new_block[2]),
        .I4(round_key[98]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[2]_i_2 
       (.I0(mixcolumns_return066_out[2]),
        .I1(new_sboxw[2]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[61]),
        .I5(round_key[98]),
        .O(\block_w0_reg[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[2]_i_4__0 
       (.I0(enc_new_block[82]),
        .I1(enc_new_block[1]),
        .I2(enc_new_block[121]),
        .I3(enc_new_block[42]),
        .I4(enc_new_block[122]),
        .O(mixcolumns_return066_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[30]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[30]_i_2_n_0 ),
        .I3(enc_new_block[126]),
        .I4(round_key[126]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[30]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[30]_i_2 
       (.I0(mixcolumns_return076_out[6]),
        .I1(new_sboxw[30]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[78]),
        .I5(round_key[126]),
        .O(\block_w0_reg[30]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[30]_i_4__0 
       (.I0(enc_new_block[125]),
        .I1(enc_new_block[85]),
        .I2(enc_new_block[6]),
        .I3(enc_new_block[46]),
        .I4(enc_new_block[86]),
        .O(mixcolumns_return076_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w0_reg[31]_i_10 
       (.I0(enc_round_nr[1]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [1]),
        .O(muxed_round_nr[1]));
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w0_reg[31]_i_11 
       (.I0(enc_round_nr[0]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [0]),
        .O(muxed_round_nr[0]));
  LUT5 #(
    .INIT(32'h46464656)) 
    \block_w0_reg[31]_i_1__0 
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(update_type__0[1]),
        .I3(p_0_in[0]),
        .I4(p_0_in[1]),
        .O(block_w0_we));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[31]_i_2 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[31]_i_3_n_0 ),
        .I3(enc_new_block[127]),
        .I4(round_key[127]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[31]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[31]_i_3 
       (.I0(mixcolumns_return076_out[7]),
        .I1(new_sboxw[31]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[79]),
        .I5(round_key[127]),
        .O(\block_w0_reg[31]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[31]_i_5__0 
       (.I0(enc_new_block[126]),
        .I1(enc_new_block[86]),
        .I2(enc_new_block[7]),
        .I3(enc_new_block[47]),
        .I4(enc_new_block[87]),
        .O(mixcolumns_return076_out[7]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[3]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[3]_i_2_n_0 ),
        .I3(enc_new_block[3]),
        .I4(round_key[99]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[3]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w0_reg[3]_i_2 
       (.I0(addroundkey0_return__514[99]),
        .I1(new_sboxw[3]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[19]),
        .O(\block_w0_reg[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[3]_i_4 
       (.I0(\block_w0_reg[28]_i_9_n_0 ),
        .I1(\block_w0_reg[4]_i_4__0_n_0 ),
        .I2(enc_new_block[122]),
        .I3(round_key[99]),
        .I4(enc_new_block[43]),
        .I5(enc_new_block[2]),
        .O(addroundkey0_return__514[99]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[4]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[4]_i_2_n_0 ),
        .I3(enc_new_block[4]),
        .I4(round_key[100]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w0_reg[4]_i_2 
       (.I0(\block_w0_reg[4]_i_4__0_n_0 ),
        .I1(\block_w0_reg[4]_i_5_n_0 ),
        .I2(new_sboxw[4]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[20]),
        .O(\block_w0_reg[4]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[4]_i_4__0 
       (.I0(enc_new_block[7]),
        .I1(enc_new_block[127]),
        .O(\block_w0_reg[4]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[4]_i_5 
       (.I0(enc_new_block[44]),
        .I1(enc_new_block[84]),
        .I2(enc_new_block[123]),
        .I3(round_key[100]),
        .I4(enc_new_block[124]),
        .I5(enc_new_block[3]),
        .O(\block_w0_reg[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[5]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[5]_i_2_n_0 ),
        .I3(enc_new_block[5]),
        .I4(round_key[101]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[5]_i_2 
       (.I0(mixcolumns_return066_out[5]),
        .I1(new_sboxw[5]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[62]),
        .I5(round_key[101]),
        .O(\block_w0_reg[5]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[5]_i_4__0 
       (.I0(enc_new_block[85]),
        .I1(enc_new_block[4]),
        .I2(enc_new_block[124]),
        .I3(enc_new_block[45]),
        .I4(enc_new_block[125]),
        .O(mixcolumns_return066_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[6]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[6]_i_2_n_0 ),
        .I3(enc_new_block[6]),
        .I4(round_key[102]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[6]_i_2 
       (.I0(mixcolumns_return066_out[6]),
        .I1(new_sboxw[6]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[63]),
        .I5(round_key[102]),
        .O(\block_w0_reg[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[6]_i_4__0 
       (.I0(enc_new_block[86]),
        .I1(enc_new_block[5]),
        .I2(enc_new_block[125]),
        .I3(enc_new_block[46]),
        .I4(enc_new_block[126]),
        .O(mixcolumns_return066_out[6]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[7]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[7]_i_2_n_0 ),
        .I3(enc_new_block[7]),
        .I4(round_key[103]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[7]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[7]_i_2 
       (.I0(mixcolumns_return066_out[7]),
        .I1(new_sboxw[7]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[64]),
        .I5(round_key[103]),
        .O(\block_w0_reg[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[7]_i_4__0 
       (.I0(enc_new_block[87]),
        .I1(enc_new_block[6]),
        .I2(enc_new_block[126]),
        .I3(enc_new_block[47]),
        .I4(enc_new_block[127]),
        .O(mixcolumns_return066_out[7]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[8]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[8]_i_2_n_0 ),
        .I3(enc_new_block[40]),
        .I4(round_key[104]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[8]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w0_reg[8]_i_2 
       (.I0(mixcolumns_return070_out[0]),
        .I1(new_sboxw[8]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[65]),
        .I5(round_key[104]),
        .O(\block_w0_reg[8]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[8]_i_4__0 
       (.I0(enc_new_block[80]),
        .I1(enc_new_block[7]),
        .I2(enc_new_block[47]),
        .I3(enc_new_block[0]),
        .I4(enc_new_block[120]),
        .O(mixcolumns_return070_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w0_reg[9]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w0_reg[9]_i_2_n_0 ),
        .I3(enc_new_block[41]),
        .I4(round_key[105]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w0_reg[9]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w0_reg[9]_i_2 
       (.I0(\block_w0_reg[9]_i_4__0_n_0 ),
        .I1(\block_w0_reg[9]_i_5_n_0 ),
        .I2(new_sboxw[9]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[21]),
        .O(\block_w0_reg[9]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[9]_i_4__0 
       (.I0(enc_new_block[47]),
        .I1(enc_new_block[7]),
        .O(\block_w0_reg[9]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[9]_i_5 
       (.I0(enc_new_block[40]),
        .I1(enc_new_block[1]),
        .I2(enc_new_block[0]),
        .I3(round_key[105]),
        .I4(enc_new_block[81]),
        .I5(enc_new_block[121]),
        .O(\block_w0_reg[9]_i_5_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[0] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[0]_i_1__0_n_0 ),
        .Q(enc_new_block[96]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[10] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[10]_i_1_n_0 ),
        .Q(enc_new_block[106]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[11] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[11]_i_1_n_0 ),
        .Q(enc_new_block[107]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[12] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[12]_i_1_n_0 ),
        .Q(enc_new_block[108]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[13] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[13]_i_1_n_0 ),
        .Q(enc_new_block[109]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[14] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[14]_i_1_n_0 ),
        .Q(enc_new_block[110]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[15] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[15]_i_1_n_0 ),
        .Q(enc_new_block[111]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[16] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[16]_i_1__0_n_0 ),
        .Q(enc_new_block[112]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[17] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[17]_i_1_n_0 ),
        .Q(enc_new_block[113]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[18] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[18]_i_1_n_0 ),
        .Q(enc_new_block[114]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[19] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[19]_i_1_n_0 ),
        .Q(enc_new_block[115]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[1] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[1]_i_1_n_0 ),
        .Q(enc_new_block[97]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[20] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[20]_i_1_n_0 ),
        .Q(enc_new_block[116]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[21] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[21]_i_1_n_0 ),
        .Q(enc_new_block[117]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[22] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[22]_i_1_n_0 ),
        .Q(enc_new_block[118]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[23] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[23]_i_1_n_0 ),
        .Q(enc_new_block[119]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[24] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[24]_i_1_n_0 ),
        .Q(enc_new_block[120]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[25] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[25]_i_1_n_0 ),
        .Q(enc_new_block[121]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[26] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[26]_i_1_n_0 ),
        .Q(enc_new_block[122]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[27] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[27]_i_1_n_0 ),
        .Q(enc_new_block[123]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[28] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[28]_i_1_n_0 ),
        .Q(enc_new_block[124]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[29] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[29]_i_1_n_0 ),
        .Q(enc_new_block[125]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[2] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[2]_i_1_n_0 ),
        .Q(enc_new_block[98]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[30] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[30]_i_1_n_0 ),
        .Q(enc_new_block[126]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[31] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[31]_i_2_n_0 ),
        .Q(enc_new_block[127]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[3] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[3]_i_1_n_0 ),
        .Q(enc_new_block[99]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[4] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[4]_i_1_n_0 ),
        .Q(enc_new_block[100]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[5] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[5]_i_1_n_0 ),
        .Q(enc_new_block[101]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[6] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[6]_i_1_n_0 ),
        .Q(enc_new_block[102]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[7] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[7]_i_1_n_0 ),
        .Q(enc_new_block[103]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[8] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[8]_i_1_n_0 ),
        .Q(enc_new_block[104]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w0_reg_reg[9] 
       (.C(clk_i),
        .CE(block_w0_we),
        .CLR(rst_i),
        .D(\block_w0_reg[9]_i_1_n_0 ),
        .Q(enc_new_block[105]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[0]_i_1__0 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[0]_i_2_n_0 ),
        .I3(enc_new_block[96]),
        .I4(round_key[64]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[0]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[0]_i_2 
       (.I0(mixcolumns_return050_out[0]),
        .I1(new_sboxw[0]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[40]),
        .I5(round_key[64]),
        .O(\block_w1_reg[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[0]_i_4__0 
       (.I0(enc_new_block[103]),
        .I1(enc_new_block[95]),
        .I2(enc_new_block[88]),
        .I3(enc_new_block[48]),
        .I4(enc_new_block[8]),
        .O(mixcolumns_return050_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[10]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[10]_i_2_n_0 ),
        .I3(enc_new_block[10]),
        .I4(round_key[74]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[10]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[10]_i_2 
       (.I0(mixcolumns_return054_out[2]),
        .I1(new_sboxw[10]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[46]),
        .I5(round_key[74]),
        .O(\block_w1_reg[10]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[10]_i_4__0 
       (.I0(enc_new_block[98]),
        .I1(enc_new_block[9]),
        .I2(enc_new_block[90]),
        .I3(enc_new_block[50]),
        .I4(enc_new_block[97]),
        .O(mixcolumns_return054_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[11]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[11]_i_2_n_0 ),
        .I3(enc_new_block[11]),
        .I4(round_key[75]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[11]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w1_reg[11]_i_2 
       (.I0(addroundkey0_return__514[75]),
        .I1(new_sboxw[11]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[13]),
        .O(\block_w1_reg[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[11]_i_4__0 
       (.I0(\block_w1_reg[28]_i_9_n_0 ),
        .I1(\block_w1_reg[9]_i_4__0_n_0 ),
        .I2(enc_new_block[98]),
        .I3(round_key[75]),
        .I4(enc_new_block[10]),
        .I5(enc_new_block[99]),
        .O(addroundkey0_return__514[75]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[12]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[12]_i_2_n_0 ),
        .I3(enc_new_block[12]),
        .I4(round_key[76]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[12]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w1_reg[12]_i_2 
       (.I0(addroundkey0_return__514[76]),
        .I1(new_sboxw[12]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[14]),
        .O(\block_w1_reg[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[12]_i_4 
       (.I0(\block_w1_reg[27]_i_9_n_0 ),
        .I1(\block_w1_reg[9]_i_4__0_n_0 ),
        .I2(enc_new_block[52]),
        .I3(round_key[76]),
        .I4(enc_new_block[100]),
        .I5(enc_new_block[92]),
        .O(addroundkey0_return__514[76]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[13]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[13]_i_2_n_0 ),
        .I3(enc_new_block[13]),
        .I4(round_key[77]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[13]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[13]_i_2 
       (.I0(mixcolumns_return054_out[5]),
        .I1(new_sboxw[13]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[47]),
        .I5(round_key[77]),
        .O(\block_w1_reg[13]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[13]_i_4__0 
       (.I0(enc_new_block[101]),
        .I1(enc_new_block[12]),
        .I2(enc_new_block[93]),
        .I3(enc_new_block[53]),
        .I4(enc_new_block[100]),
        .O(mixcolumns_return054_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[14]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[14]_i_2_n_0 ),
        .I3(enc_new_block[14]),
        .I4(round_key[78]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[14]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[14]_i_2 
       (.I0(mixcolumns_return054_out[6]),
        .I1(new_sboxw[14]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[48]),
        .I5(round_key[78]),
        .O(\block_w1_reg[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[14]_i_4__0 
       (.I0(enc_new_block[102]),
        .I1(enc_new_block[13]),
        .I2(enc_new_block[94]),
        .I3(enc_new_block[54]),
        .I4(enc_new_block[101]),
        .O(mixcolumns_return054_out[6]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[15]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[15]_i_2_n_0 ),
        .I3(enc_new_block[15]),
        .I4(round_key[79]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[15]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[15]_i_2 
       (.I0(mixcolumns_return054_out[7]),
        .I1(new_sboxw[15]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[49]),
        .I5(round_key[79]),
        .O(\block_w1_reg[15]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[15]_i_4__0 
       (.I0(enc_new_block[103]),
        .I1(enc_new_block[14]),
        .I2(enc_new_block[95]),
        .I3(enc_new_block[55]),
        .I4(enc_new_block[102]),
        .O(mixcolumns_return054_out[7]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[16]_i_1__0 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[16]_i_2_n_0 ),
        .I3(enc_new_block[48]),
        .I4(round_key[80]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[16]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[16]_i_2 
       (.I0(mixcolumns_return057_out[0]),
        .I1(new_sboxw[16]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[50]),
        .I5(round_key[80]),
        .O(\block_w1_reg[16]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[16]_i_4__0 
       (.I0(enc_new_block[8]),
        .I1(enc_new_block[15]),
        .I2(enc_new_block[55]),
        .I3(enc_new_block[88]),
        .I4(enc_new_block[96]),
        .O(mixcolumns_return057_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[17]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[17]_i_2_n_0 ),
        .I3(enc_new_block[49]),
        .I4(round_key[81]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[17]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w1_reg[17]_i_2 
       (.I0(\block_w1_reg[20]_i_4__0_n_0 ),
        .I1(\block_w1_reg[17]_i_4_n_0 ),
        .I2(new_sboxw[17]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(addroundkey_return[15]),
        .O(\block_w1_reg[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[17]_i_4 
       (.I0(enc_new_block[8]),
        .I1(enc_new_block[48]),
        .I2(enc_new_block[89]),
        .I3(round_key[81]),
        .I4(enc_new_block[97]),
        .I5(enc_new_block[9]),
        .O(\block_w1_reg[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[18]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[18]_i_2_n_0 ),
        .I3(enc_new_block[50]),
        .I4(round_key[82]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[18]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[18]_i_2 
       (.I0(mixcolumns_return057_out[2]),
        .I1(new_sboxw[18]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[51]),
        .I5(round_key[82]),
        .O(\block_w1_reg[18]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[18]_i_4__0 
       (.I0(enc_new_block[10]),
        .I1(enc_new_block[9]),
        .I2(enc_new_block[49]),
        .I3(enc_new_block[90]),
        .I4(enc_new_block[98]),
        .O(mixcolumns_return057_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[19]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[19]_i_2_n_0 ),
        .I3(enc_new_block[51]),
        .I4(round_key[83]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[19]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w1_reg[19]_i_2 
       (.I0(addroundkey0_return__514[83]),
        .I1(new_sboxw[19]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(addroundkey_return[16]),
        .O(\block_w1_reg[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[19]_i_4 
       (.I0(\block_w1_reg[20]_i_4__0_n_0 ),
        .I1(\block_w1_reg[27]_i_9_n_0 ),
        .I2(enc_new_block[91]),
        .I3(round_key[83]),
        .I4(enc_new_block[50]),
        .I5(enc_new_block[10]),
        .O(addroundkey0_return__514[83]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[1]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[1]_i_2_n_0 ),
        .I3(enc_new_block[97]),
        .I4(round_key[65]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w1_reg[1]_i_2 
       (.I0(\block_w1_reg[4]_i_4__0_n_0 ),
        .I1(\block_w1_reg[1]_i_4_n_0 ),
        .I2(new_sboxw[1]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(addroundkey_return[12]),
        .O(\block_w1_reg[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[1]_i_4 
       (.I0(enc_new_block[96]),
        .I1(enc_new_block[88]),
        .I2(enc_new_block[49]),
        .I3(round_key[65]),
        .I4(enc_new_block[9]),
        .I5(enc_new_block[89]),
        .O(\block_w1_reg[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[20]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[20]_i_2_n_0 ),
        .I3(enc_new_block[52]),
        .I4(round_key[84]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[20]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w1_reg[20]_i_2 
       (.I0(\block_w1_reg[20]_i_4__0_n_0 ),
        .I1(\block_w1_reg[20]_i_5__0_n_0 ),
        .I2(new_sboxw[20]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(addroundkey_return[17]),
        .O(\block_w1_reg[20]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[20]_i_4__0 
       (.I0(enc_new_block[55]),
        .I1(enc_new_block[15]),
        .O(\block_w1_reg[20]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[20]_i_5__0 
       (.I0(enc_new_block[12]),
        .I1(enc_new_block[100]),
        .I2(enc_new_block[51]),
        .I3(round_key[84]),
        .I4(enc_new_block[92]),
        .I5(enc_new_block[11]),
        .O(\block_w1_reg[20]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[21]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[21]_i_2_n_0 ),
        .I3(enc_new_block[53]),
        .I4(round_key[85]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[21]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[21]_i_2 
       (.I0(mixcolumns_return057_out[5]),
        .I1(new_sboxw[21]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[52]),
        .I5(round_key[85]),
        .O(\block_w1_reg[21]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[21]_i_4__0 
       (.I0(enc_new_block[13]),
        .I1(enc_new_block[12]),
        .I2(enc_new_block[52]),
        .I3(enc_new_block[93]),
        .I4(enc_new_block[101]),
        .O(mixcolumns_return057_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[22]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[22]_i_2_n_0 ),
        .I3(enc_new_block[54]),
        .I4(round_key[86]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[22]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[22]_i_2 
       (.I0(mixcolumns_return057_out[6]),
        .I1(new_sboxw[22]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[53]),
        .I5(round_key[86]),
        .O(\block_w1_reg[22]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[22]_i_4__0 
       (.I0(enc_new_block[14]),
        .I1(enc_new_block[13]),
        .I2(enc_new_block[53]),
        .I3(enc_new_block[94]),
        .I4(enc_new_block[102]),
        .O(mixcolumns_return057_out[6]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[23]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[23]_i_2_n_0 ),
        .I3(enc_new_block[55]),
        .I4(round_key[87]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[23]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[23]_i_2 
       (.I0(mixcolumns_return057_out[7]),
        .I1(new_sboxw[23]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[54]),
        .I5(round_key[87]),
        .O(\block_w1_reg[23]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[23]_i_4__0 
       (.I0(enc_new_block[15]),
        .I1(enc_new_block[14]),
        .I2(enc_new_block[54]),
        .I3(enc_new_block[95]),
        .I4(enc_new_block[103]),
        .O(mixcolumns_return057_out[7]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[24]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[24]_i_2_n_0 ),
        .I3(enc_new_block[88]),
        .I4(round_key[88]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[24]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[24]_i_2 
       (.I0(mixcolumns_return060_out[0]),
        .I1(new_sboxw[24]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[55]),
        .I5(round_key[88]),
        .O(\block_w1_reg[24]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[24]_i_4__0 
       (.I0(enc_new_block[55]),
        .I1(enc_new_block[96]),
        .I2(enc_new_block[95]),
        .I3(enc_new_block[8]),
        .I4(enc_new_block[48]),
        .O(mixcolumns_return060_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[25]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[25]_i_2_n_0 ),
        .I3(enc_new_block[89]),
        .I4(round_key[89]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[25]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w1_reg[25]_i_2 
       (.I0(\block_w1_reg[25]_i_4__0_n_0 ),
        .I1(\block_w1_reg[25]_i_5__0_n_0 ),
        .I2(new_sboxw[25]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[15]),
        .O(\block_w1_reg[25]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[25]_i_4__0 
       (.I0(enc_new_block[55]),
        .I1(enc_new_block[95]),
        .O(\block_w1_reg[25]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[25]_i_5__0 
       (.I0(enc_new_block[97]),
        .I1(enc_new_block[48]),
        .I2(enc_new_block[49]),
        .I3(round_key[89]),
        .I4(enc_new_block[88]),
        .I5(enc_new_block[9]),
        .O(\block_w1_reg[25]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[26]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[26]_i_2_n_0 ),
        .I3(enc_new_block[90]),
        .I4(round_key[90]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[26]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[26]_i_2 
       (.I0(mixcolumns_return060_out[2]),
        .I1(new_sboxw[26]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[56]),
        .I5(round_key[90]),
        .O(\block_w1_reg[26]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[26]_i_4__0 
       (.I0(enc_new_block[49]),
        .I1(enc_new_block[98]),
        .I2(enc_new_block[89]),
        .I3(enc_new_block[10]),
        .I4(enc_new_block[50]),
        .O(mixcolumns_return060_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[27]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[27]_i_2_n_0 ),
        .I3(enc_new_block[91]),
        .I4(round_key[91]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[27]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w1_reg[27]_i_2 
       (.I0(addroundkey0_return__514[91]),
        .I1(new_sboxw[27]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[16]),
        .O(\block_w1_reg[27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[27]_i_4__0 
       (.I0(\block_w1_reg[27]_i_9_n_0 ),
        .I1(\block_w1_reg[25]_i_4__0_n_0 ),
        .I2(enc_new_block[51]),
        .I3(round_key[91]),
        .I4(enc_new_block[50]),
        .I5(enc_new_block[90]),
        .O(addroundkey0_return__514[91]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[27]_i_9 
       (.I0(enc_new_block[99]),
        .I1(enc_new_block[11]),
        .O(\block_w1_reg[27]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[28]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[28]_i_2_n_0 ),
        .I3(enc_new_block[92]),
        .I4(round_key[92]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[28]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w1_reg[28]_i_2 
       (.I0(addroundkey0_return__514[92]),
        .I1(new_sboxw[28]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[17]),
        .O(\block_w1_reg[28]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[28]_i_4 
       (.I0(\block_w1_reg[28]_i_9_n_0 ),
        .I1(\block_w1_reg[25]_i_4__0_n_0 ),
        .I2(enc_new_block[52]),
        .I3(round_key[92]),
        .I4(enc_new_block[100]),
        .I5(enc_new_block[12]),
        .O(addroundkey0_return__514[92]));
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[28]_i_9 
       (.I0(enc_new_block[91]),
        .I1(enc_new_block[51]),
        .O(\block_w1_reg[28]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[29]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[29]_i_2_n_0 ),
        .I3(enc_new_block[93]),
        .I4(round_key[93]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[29]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[29]_i_2 
       (.I0(mixcolumns_return060_out[5]),
        .I1(new_sboxw[29]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[57]),
        .I5(round_key[93]),
        .O(\block_w1_reg[29]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[29]_i_4__0 
       (.I0(enc_new_block[52]),
        .I1(enc_new_block[101]),
        .I2(enc_new_block[92]),
        .I3(enc_new_block[13]),
        .I4(enc_new_block[53]),
        .O(mixcolumns_return060_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[2]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[2]_i_2_n_0 ),
        .I3(enc_new_block[98]),
        .I4(round_key[66]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[2]_i_2 
       (.I0(mixcolumns_return050_out[2]),
        .I1(new_sboxw[2]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[41]),
        .I5(round_key[66]),
        .O(\block_w1_reg[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[2]_i_4__0 
       (.I0(enc_new_block[97]),
        .I1(enc_new_block[89]),
        .I2(enc_new_block[90]),
        .I3(enc_new_block[50]),
        .I4(enc_new_block[10]),
        .O(mixcolumns_return050_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[30]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[30]_i_2_n_0 ),
        .I3(enc_new_block[94]),
        .I4(round_key[94]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[30]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[30]_i_2 
       (.I0(mixcolumns_return060_out[6]),
        .I1(new_sboxw[30]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[58]),
        .I5(round_key[94]),
        .O(\block_w1_reg[30]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[30]_i_4__0 
       (.I0(enc_new_block[53]),
        .I1(enc_new_block[102]),
        .I2(enc_new_block[93]),
        .I3(enc_new_block[14]),
        .I4(enc_new_block[54]),
        .O(mixcolumns_return060_out[6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w1_reg[31]_i_10 
       (.I0(enc_round_nr[1]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [1]),
        .O(\round_ctr_reg_reg[1]_2 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w1_reg[31]_i_11 
       (.I0(enc_round_nr[0]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [0]),
        .O(\round_ctr_reg_reg[0]_0 ));
  LUT5 #(
    .INIT(32'h45446666)) 
    \block_w1_reg[31]_i_1__0 
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(p_0_in[1]),
        .I3(p_0_in[0]),
        .I4(update_type__0[1]),
        .O(block_w1_we));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[31]_i_2 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[31]_i_3_n_0 ),
        .I3(enc_new_block[95]),
        .I4(round_key[95]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[31]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[31]_i_3 
       (.I0(mixcolumns_return060_out[7]),
        .I1(new_sboxw[31]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[59]),
        .I5(round_key[95]),
        .O(\block_w1_reg[31]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[31]_i_5__0 
       (.I0(enc_new_block[54]),
        .I1(enc_new_block[103]),
        .I2(enc_new_block[94]),
        .I3(enc_new_block[15]),
        .I4(enc_new_block[55]),
        .O(mixcolumns_return060_out[7]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[3]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[3]_i_2_n_0 ),
        .I3(enc_new_block[99]),
        .I4(round_key[67]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[3]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w1_reg[3]_i_2 
       (.I0(addroundkey0_return__514[67]),
        .I1(new_sboxw[3]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(addroundkey_return[13]),
        .O(\block_w1_reg[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[3]_i_4 
       (.I0(\block_w1_reg[28]_i_9_n_0 ),
        .I1(\block_w1_reg[4]_i_4__0_n_0 ),
        .I2(enc_new_block[11]),
        .I3(round_key[67]),
        .I4(enc_new_block[90]),
        .I5(enc_new_block[98]),
        .O(addroundkey0_return__514[67]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[4]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[4]_i_2_n_0 ),
        .I3(enc_new_block[100]),
        .I4(round_key[68]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w1_reg[4]_i_2 
       (.I0(\block_w1_reg[4]_i_4__0_n_0 ),
        .I1(\block_w1_reg[4]_i_5_n_0 ),
        .I2(new_sboxw[4]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(addroundkey_return[14]),
        .O(\block_w1_reg[4]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[4]_i_4__0 
       (.I0(enc_new_block[95]),
        .I1(enc_new_block[103]),
        .O(\block_w1_reg[4]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[4]_i_5 
       (.I0(enc_new_block[12]),
        .I1(enc_new_block[99]),
        .I2(enc_new_block[91]),
        .I3(round_key[68]),
        .I4(enc_new_block[92]),
        .I5(enc_new_block[52]),
        .O(\block_w1_reg[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[5]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[5]_i_2_n_0 ),
        .I3(enc_new_block[101]),
        .I4(round_key[69]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[5]_i_2 
       (.I0(mixcolumns_return050_out[5]),
        .I1(new_sboxw[5]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[42]),
        .I5(round_key[69]),
        .O(\block_w1_reg[5]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[5]_i_4__0 
       (.I0(enc_new_block[100]),
        .I1(enc_new_block[92]),
        .I2(enc_new_block[93]),
        .I3(enc_new_block[53]),
        .I4(enc_new_block[13]),
        .O(mixcolumns_return050_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[6]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[6]_i_2_n_0 ),
        .I3(enc_new_block[102]),
        .I4(round_key[70]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[6]_i_2 
       (.I0(mixcolumns_return050_out[6]),
        .I1(new_sboxw[6]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[43]),
        .I5(round_key[70]),
        .O(\block_w1_reg[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[6]_i_4__0 
       (.I0(enc_new_block[101]),
        .I1(enc_new_block[93]),
        .I2(enc_new_block[94]),
        .I3(enc_new_block[54]),
        .I4(enc_new_block[14]),
        .O(mixcolumns_return050_out[6]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[7]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[7]_i_2_n_0 ),
        .I3(enc_new_block[103]),
        .I4(round_key[71]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[7]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[7]_i_2 
       (.I0(mixcolumns_return050_out[7]),
        .I1(new_sboxw[7]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[44]),
        .I5(round_key[71]),
        .O(\block_w1_reg[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[7]_i_4__0 
       (.I0(enc_new_block[102]),
        .I1(enc_new_block[94]),
        .I2(enc_new_block[95]),
        .I3(enc_new_block[55]),
        .I4(enc_new_block[15]),
        .O(mixcolumns_return050_out[7]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[8]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[8]_i_2_n_0 ),
        .I3(enc_new_block[8]),
        .I4(round_key[72]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[8]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w1_reg[8]_i_2 
       (.I0(mixcolumns_return054_out[0]),
        .I1(new_sboxw[8]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[45]),
        .I5(round_key[72]),
        .O(\block_w1_reg[8]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[8]_i_4__0 
       (.I0(enc_new_block[96]),
        .I1(enc_new_block[15]),
        .I2(enc_new_block[88]),
        .I3(enc_new_block[48]),
        .I4(enc_new_block[103]),
        .O(mixcolumns_return054_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w1_reg[9]_i_1__0 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w1_reg[9]_i_2_n_0 ),
        .I3(enc_new_block[9]),
        .I4(round_key[73]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w1_reg[9]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w1_reg[9]_i_2 
       (.I0(\block_w1_reg[9]_i_4__0_n_0 ),
        .I1(\block_w1_reg[9]_i_5__0_n_0 ),
        .I2(new_sboxw[9]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[12]),
        .O(\block_w1_reg[9]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[9]_i_4__0 
       (.I0(enc_new_block[15]),
        .I1(enc_new_block[103]),
        .O(\block_w1_reg[9]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[9]_i_5__0 
       (.I0(enc_new_block[97]),
        .I1(enc_new_block[8]),
        .I2(enc_new_block[49]),
        .I3(round_key[73]),
        .I4(enc_new_block[96]),
        .I5(enc_new_block[89]),
        .O(\block_w1_reg[9]_i_5__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[0] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[0]_i_1__0_n_0 ),
        .Q(enc_new_block[64]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[10] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[10]_i_1_n_0 ),
        .Q(enc_new_block[74]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[11] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[11]_i_1_n_0 ),
        .Q(enc_new_block[75]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[12] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[12]_i_1_n_0 ),
        .Q(enc_new_block[76]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[13] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[13]_i_1_n_0 ),
        .Q(enc_new_block[77]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[14] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[14]_i_1_n_0 ),
        .Q(enc_new_block[78]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[15] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[15]_i_1_n_0 ),
        .Q(enc_new_block[79]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[16] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[16]_i_1__0_n_0 ),
        .Q(enc_new_block[80]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[17] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[17]_i_1_n_0 ),
        .Q(enc_new_block[81]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[18] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[18]_i_1_n_0 ),
        .Q(enc_new_block[82]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[19] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[19]_i_1_n_0 ),
        .Q(enc_new_block[83]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[1] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[1]_i_1_n_0 ),
        .Q(enc_new_block[65]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[20] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[20]_i_1_n_0 ),
        .Q(enc_new_block[84]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[21] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[21]_i_1_n_0 ),
        .Q(enc_new_block[85]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[22] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[22]_i_1_n_0 ),
        .Q(enc_new_block[86]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[23] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[23]_i_1_n_0 ),
        .Q(enc_new_block[87]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[24] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[24]_i_1_n_0 ),
        .Q(enc_new_block[88]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[25] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[25]_i_1_n_0 ),
        .Q(enc_new_block[89]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[26] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[26]_i_1_n_0 ),
        .Q(enc_new_block[90]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[27] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[27]_i_1_n_0 ),
        .Q(enc_new_block[91]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[28] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[28]_i_1_n_0 ),
        .Q(enc_new_block[92]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[29] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[29]_i_1_n_0 ),
        .Q(enc_new_block[93]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[2] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[2]_i_1_n_0 ),
        .Q(enc_new_block[66]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[30] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[30]_i_1_n_0 ),
        .Q(enc_new_block[94]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[31] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[31]_i_2_n_0 ),
        .Q(enc_new_block[95]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[3] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[3]_i_1_n_0 ),
        .Q(enc_new_block[67]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[4] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[4]_i_1_n_0 ),
        .Q(enc_new_block[68]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[5] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[5]_i_1_n_0 ),
        .Q(enc_new_block[69]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[6] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[6]_i_1_n_0 ),
        .Q(enc_new_block[70]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[7] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[7]_i_1_n_0 ),
        .Q(enc_new_block[71]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[8] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[8]_i_1_n_0 ),
        .Q(enc_new_block[72]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w1_reg_reg[9] 
       (.C(clk_i),
        .CE(block_w1_we),
        .CLR(rst_i),
        .D(\block_w1_reg[9]_i_1__0_n_0 ),
        .Q(enc_new_block[73]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[0]_i_1__0 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[0]_i_2_n_0 ),
        .I3(enc_new_block[64]),
        .I4(round_key[32]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[0]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[0]_i_2 
       (.I0(mixcolumns_return034_out[0]),
        .I1(new_sboxw[0]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[20]),
        .I5(round_key[32]),
        .O(\block_w2_reg[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[0]_i_4__0 
       (.I0(enc_new_block[104]),
        .I1(enc_new_block[63]),
        .I2(enc_new_block[56]),
        .I3(enc_new_block[16]),
        .I4(enc_new_block[71]),
        .O(mixcolumns_return034_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[10]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[10]_i_2_n_0 ),
        .I3(enc_new_block[106]),
        .I4(round_key[42]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[10]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[10]_i_2 
       (.I0(mixcolumns_return038_out[2]),
        .I1(new_sboxw[10]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[26]),
        .I5(round_key[42]),
        .O(\block_w2_reg[10]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[10]_i_4__0 
       (.I0(enc_new_block[105]),
        .I1(enc_new_block[66]),
        .I2(enc_new_block[58]),
        .I3(enc_new_block[18]),
        .I4(enc_new_block[65]),
        .O(mixcolumns_return038_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[11]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[11]_i_2_n_0 ),
        .I3(enc_new_block[107]),
        .I4(round_key[43]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[11]));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w2_reg[11]_i_2 
       (.I0(addroundkey0_return__514[43]),
        .I1(new_sboxw[11]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(addroundkey_return[10]),
        .O(\block_w2_reg[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[11]_i_4__0 
       (.I0(\block_w2_reg[28]_i_10_n_0 ),
        .I1(\block_w2_reg[9]_i_4__0_n_0 ),
        .I2(enc_new_block[66]),
        .I3(round_key[43]),
        .I4(enc_new_block[106]),
        .I5(enc_new_block[67]),
        .O(addroundkey0_return__514[43]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[12]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[12]_i_2_n_0 ),
        .I3(enc_new_block[108]),
        .I4(round_key[44]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[12]));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w2_reg[12]_i_2 
       (.I0(addroundkey0_return__514[44]),
        .I1(new_sboxw[12]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(addroundkey_return[11]),
        .O(\block_w2_reg[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[12]_i_4 
       (.I0(\block_w2_reg[27]_i_11_n_0 ),
        .I1(\block_w2_reg[9]_i_4__0_n_0 ),
        .I2(enc_new_block[20]),
        .I3(round_key[44]),
        .I4(enc_new_block[68]),
        .I5(enc_new_block[60]),
        .O(addroundkey0_return__514[44]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[13]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[13]_i_2_n_0 ),
        .I3(enc_new_block[109]),
        .I4(round_key[45]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[13]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[13]_i_2 
       (.I0(mixcolumns_return038_out[5]),
        .I1(new_sboxw[13]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[27]),
        .I5(round_key[45]),
        .O(\block_w2_reg[13]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[13]_i_4__0 
       (.I0(enc_new_block[108]),
        .I1(enc_new_block[69]),
        .I2(enc_new_block[61]),
        .I3(enc_new_block[21]),
        .I4(enc_new_block[68]),
        .O(mixcolumns_return038_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[14]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[14]_i_2_n_0 ),
        .I3(enc_new_block[110]),
        .I4(round_key[46]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[14]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[14]_i_2 
       (.I0(mixcolumns_return038_out[6]),
        .I1(new_sboxw[14]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[28]),
        .I5(round_key[46]),
        .O(\block_w2_reg[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[14]_i_4__0 
       (.I0(enc_new_block[109]),
        .I1(enc_new_block[70]),
        .I2(enc_new_block[62]),
        .I3(enc_new_block[22]),
        .I4(enc_new_block[69]),
        .O(mixcolumns_return038_out[6]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[15]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[15]_i_2_n_0 ),
        .I3(enc_new_block[111]),
        .I4(round_key[47]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[15]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w2_reg[15]_i_13 
       (.I0(enc_new_block[79]),
        .I1(enc_new_block[111]),
        .I2(enc_new_block[15]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[47]),
        .O(muxed_sboxw__0[15]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    \block_w2_reg[15]_i_14 
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[14]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[14]),
        .I5(init_state),
        .O(\prev_key1_reg_reg[31] [2]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w2_reg[15]_i_15 
       (.I0(enc_new_block[78]),
        .I1(enc_new_block[110]),
        .I2(enc_new_block[14]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[46]),
        .O(muxed_sboxw__0[14]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[15]_i_2 
       (.I0(mixcolumns_return038_out[7]),
        .I1(new_sboxw[15]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[29]),
        .I5(round_key[47]),
        .O(\block_w2_reg[15]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[15]_i_4__0 
       (.I0(enc_new_block[110]),
        .I1(enc_new_block[71]),
        .I2(enc_new_block[63]),
        .I3(enc_new_block[23]),
        .I4(enc_new_block[70]),
        .O(mixcolumns_return038_out[7]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    \block_w2_reg[15]_i_9 
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[15]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[15]),
        .I5(init_state),
        .O(\prev_key1_reg_reg[31] [3]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[16]_i_1__0 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[16]_i_2_n_0 ),
        .I3(enc_new_block[16]),
        .I4(round_key[48]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[16]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[16]_i_2 
       (.I0(mixcolumns_return041_out[0]),
        .I1(new_sboxw[16]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[30]),
        .I5(round_key[48]),
        .O(\block_w2_reg[16]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[16]_i_4__0 
       (.I0(enc_new_block[23]),
        .I1(enc_new_block[111]),
        .I2(enc_new_block[104]),
        .I3(enc_new_block[64]),
        .I4(enc_new_block[56]),
        .O(mixcolumns_return041_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[17]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[17]_i_2_n_0 ),
        .I3(enc_new_block[17]),
        .I4(round_key[49]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[17]));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w2_reg[17]_i_2 
       (.I0(\block_w2_reg[20]_i_4__0_n_0 ),
        .I1(\block_w2_reg[17]_i_4_n_0 ),
        .I2(new_sboxw[17]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[6]),
        .O(\block_w2_reg[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[17]_i_4 
       (.I0(enc_new_block[65]),
        .I1(enc_new_block[16]),
        .I2(enc_new_block[57]),
        .I3(round_key[49]),
        .I4(enc_new_block[104]),
        .I5(enc_new_block[105]),
        .O(\block_w2_reg[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[18]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[18]_i_2_n_0 ),
        .I3(enc_new_block[18]),
        .I4(round_key[50]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[18]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[18]_i_2 
       (.I0(mixcolumns_return041_out[2]),
        .I1(new_sboxw[18]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[31]),
        .I5(round_key[50]),
        .O(\block_w2_reg[18]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[18]_i_4__0 
       (.I0(enc_new_block[17]),
        .I1(enc_new_block[105]),
        .I2(enc_new_block[106]),
        .I3(enc_new_block[66]),
        .I4(enc_new_block[58]),
        .O(mixcolumns_return041_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[19]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[19]_i_2_n_0 ),
        .I3(enc_new_block[19]),
        .I4(round_key[51]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[19]));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w2_reg[19]_i_2 
       (.I0(addroundkey0_return__514[51]),
        .I1(new_sboxw[19]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[7]),
        .O(\block_w2_reg[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[19]_i_4 
       (.I0(\block_w2_reg[20]_i_4__0_n_0 ),
        .I1(\block_w2_reg[27]_i_11_n_0 ),
        .I2(enc_new_block[59]),
        .I3(round_key[51]),
        .I4(enc_new_block[18]),
        .I5(enc_new_block[106]),
        .O(addroundkey0_return__514[51]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[1]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[1]_i_2_n_0 ),
        .I3(enc_new_block[65]),
        .I4(round_key[33]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[1]));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w2_reg[1]_i_2 
       (.I0(\block_w2_reg[4]_i_4__0_n_0 ),
        .I1(\block_w2_reg[1]_i_4_n_0 ),
        .I2(new_sboxw[1]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[3]),
        .O(\block_w2_reg[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[1]_i_4 
       (.I0(enc_new_block[105]),
        .I1(enc_new_block[56]),
        .I2(enc_new_block[17]),
        .I3(round_key[33]),
        .I4(enc_new_block[64]),
        .I5(enc_new_block[57]),
        .O(\block_w2_reg[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[20]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[20]_i_2_n_0 ),
        .I3(enc_new_block[20]),
        .I4(round_key[52]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[20]));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w2_reg[20]_i_2 
       (.I0(\block_w2_reg[20]_i_4__0_n_0 ),
        .I1(\block_w2_reg[20]_i_5__0_n_0 ),
        .I2(new_sboxw[20]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[8]),
        .O(\block_w2_reg[20]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[20]_i_4__0 
       (.I0(enc_new_block[23]),
        .I1(enc_new_block[111]),
        .O(\block_w2_reg[20]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[20]_i_5__0 
       (.I0(enc_new_block[108]),
        .I1(enc_new_block[68]),
        .I2(enc_new_block[19]),
        .I3(round_key[52]),
        .I4(enc_new_block[60]),
        .I5(enc_new_block[107]),
        .O(\block_w2_reg[20]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[21]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[21]_i_2_n_0 ),
        .I3(enc_new_block[21]),
        .I4(round_key[53]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[21]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[21]_i_2 
       (.I0(mixcolumns_return041_out[5]),
        .I1(new_sboxw[21]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[32]),
        .I5(round_key[53]),
        .O(\block_w2_reg[21]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[21]_i_4__0 
       (.I0(enc_new_block[20]),
        .I1(enc_new_block[108]),
        .I2(enc_new_block[109]),
        .I3(enc_new_block[69]),
        .I4(enc_new_block[61]),
        .O(mixcolumns_return041_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[22]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[22]_i_2_n_0 ),
        .I3(enc_new_block[22]),
        .I4(round_key[54]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[22]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[22]_i_2 
       (.I0(mixcolumns_return041_out[6]),
        .I1(new_sboxw[22]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[33]),
        .I5(round_key[54]),
        .O(\block_w2_reg[22]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[22]_i_4__0 
       (.I0(enc_new_block[21]),
        .I1(enc_new_block[109]),
        .I2(enc_new_block[110]),
        .I3(enc_new_block[70]),
        .I4(enc_new_block[62]),
        .O(mixcolumns_return041_out[6]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[23]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[23]_i_2_n_0 ),
        .I3(enc_new_block[23]),
        .I4(round_key[55]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[23]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w2_reg[23]_i_13 
       (.I0(enc_new_block[87]),
        .I1(enc_new_block[119]),
        .I2(enc_new_block[23]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[55]),
        .O(muxed_sboxw__0[23]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    \block_w2_reg[23]_i_14 
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[22]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[22]),
        .I5(init_state),
        .O(\prev_key1_reg_reg[31] [4]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w2_reg[23]_i_15 
       (.I0(enc_new_block[86]),
        .I1(enc_new_block[118]),
        .I2(enc_new_block[22]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[54]),
        .O(muxed_sboxw__0[22]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[23]_i_2 
       (.I0(mixcolumns_return041_out[7]),
        .I1(new_sboxw[23]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[34]),
        .I5(round_key[55]),
        .O(\block_w2_reg[23]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[23]_i_4__0 
       (.I0(enc_new_block[22]),
        .I1(enc_new_block[110]),
        .I2(enc_new_block[111]),
        .I3(enc_new_block[71]),
        .I4(enc_new_block[63]),
        .O(mixcolumns_return041_out[7]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    \block_w2_reg[23]_i_9 
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[23]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[23]),
        .I5(init_state),
        .O(\prev_key1_reg_reg[31] [5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[24]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[24]_i_2_n_0 ),
        .I3(enc_new_block[56]),
        .I4(round_key[56]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[24]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[24]_i_2 
       (.I0(mixcolumns_return044_out[0]),
        .I1(new_sboxw[24]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[35]),
        .I5(round_key[56]),
        .O(\block_w2_reg[24]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[24]_i_4__0 
       (.I0(enc_new_block[63]),
        .I1(enc_new_block[23]),
        .I2(enc_new_block[104]),
        .I3(enc_new_block[64]),
        .I4(enc_new_block[16]),
        .O(mixcolumns_return044_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[25]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[25]_i_2_n_0 ),
        .I3(enc_new_block[57]),
        .I4(round_key[57]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[25]));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w2_reg[25]_i_2 
       (.I0(\block_w2_reg[25]_i_4__0_n_0 ),
        .I1(\block_w2_reg[25]_i_5__0_n_0 ),
        .I2(new_sboxw[25]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[9]),
        .O(\block_w2_reg[25]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[25]_i_4__0 
       (.I0(enc_new_block[23]),
        .I1(enc_new_block[63]),
        .O(\block_w2_reg[25]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[25]_i_5__0 
       (.I0(enc_new_block[65]),
        .I1(enc_new_block[16]),
        .I2(enc_new_block[17]),
        .I3(round_key[57]),
        .I4(enc_new_block[56]),
        .I5(enc_new_block[105]),
        .O(\block_w2_reg[25]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[26]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[26]_i_2_n_0 ),
        .I3(enc_new_block[58]),
        .I4(round_key[58]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[26]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[26]_i_2 
       (.I0(mixcolumns_return044_out[2]),
        .I1(new_sboxw[26]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[36]),
        .I5(round_key[58]),
        .O(\block_w2_reg[26]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[26]_i_4__0 
       (.I0(enc_new_block[57]),
        .I1(enc_new_block[17]),
        .I2(enc_new_block[106]),
        .I3(enc_new_block[66]),
        .I4(enc_new_block[18]),
        .O(mixcolumns_return044_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[27]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[27]_i_2_n_0 ),
        .I3(enc_new_block[59]),
        .I4(round_key[59]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[27]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[27]_i_11 
       (.I0(enc_new_block[67]),
        .I1(enc_new_block[107]),
        .O(\block_w2_reg[27]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w2_reg[27]_i_2 
       (.I0(addroundkey0_return__514[59]),
        .I1(new_sboxw[27]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[10]),
        .O(\block_w2_reg[27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[27]_i_4__0 
       (.I0(\block_w2_reg[27]_i_11_n_0 ),
        .I1(\block_w2_reg[25]_i_4__0_n_0 ),
        .I2(enc_new_block[19]),
        .I3(round_key[59]),
        .I4(enc_new_block[18]),
        .I5(enc_new_block[58]),
        .O(addroundkey0_return__514[59]));
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w2_reg[27]_i_8 
       (.I0(enc_round_nr[3]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [3]),
        .O(\round_ctr_reg_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[28]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[28]_i_2_n_0 ),
        .I3(enc_new_block[60]),
        .I4(round_key[60]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[28]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[28]_i_10 
       (.I0(enc_new_block[59]),
        .I1(enc_new_block[19]),
        .O(\block_w2_reg[28]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w2_reg[28]_i_2 
       (.I0(addroundkey0_return__514[60]),
        .I1(new_sboxw[28]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[11]),
        .O(\block_w2_reg[28]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[28]_i_4 
       (.I0(\block_w2_reg[28]_i_10_n_0 ),
        .I1(\block_w2_reg[25]_i_4__0_n_0 ),
        .I2(enc_new_block[20]),
        .I3(round_key[60]),
        .I4(enc_new_block[68]),
        .I5(enc_new_block[108]),
        .O(addroundkey0_return__514[60]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[29]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[29]_i_2_n_0 ),
        .I3(enc_new_block[61]),
        .I4(round_key[61]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[29]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[29]_i_2 
       (.I0(mixcolumns_return044_out[5]),
        .I1(new_sboxw[29]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[37]),
        .I5(round_key[61]),
        .O(\block_w2_reg[29]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[29]_i_4__0 
       (.I0(enc_new_block[60]),
        .I1(enc_new_block[20]),
        .I2(enc_new_block[109]),
        .I3(enc_new_block[69]),
        .I4(enc_new_block[21]),
        .O(mixcolumns_return044_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[2]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[2]_i_2_n_0 ),
        .I3(enc_new_block[66]),
        .I4(round_key[34]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[2]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[2]_i_2 
       (.I0(mixcolumns_return034_out[2]),
        .I1(new_sboxw[2]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[21]),
        .I5(round_key[34]),
        .O(\block_w2_reg[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[2]_i_4__0 
       (.I0(enc_new_block[106]),
        .I1(enc_new_block[57]),
        .I2(enc_new_block[58]),
        .I3(enc_new_block[18]),
        .I4(enc_new_block[65]),
        .O(mixcolumns_return034_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[30]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[30]_i_2_n_0 ),
        .I3(enc_new_block[62]),
        .I4(round_key[62]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[30]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[30]_i_2 
       (.I0(mixcolumns_return044_out[6]),
        .I1(new_sboxw[30]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[38]),
        .I5(round_key[62]),
        .O(\block_w2_reg[30]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[30]_i_4__0 
       (.I0(enc_new_block[61]),
        .I1(enc_new_block[21]),
        .I2(enc_new_block[110]),
        .I3(enc_new_block[70]),
        .I4(enc_new_block[22]),
        .O(mixcolumns_return044_out[6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w2_reg[31]_i_12 
       (.I0(enc_round_nr[3]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [3]),
        .O(\round_ctr_reg_reg[3]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w2_reg[31]_i_14 
       (.I0(enc_round_nr[2]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [2]),
        .O(muxed_round_nr[2]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    \block_w2_reg[31]_i_16 
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[31]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[31]),
        .I5(init_state),
        .O(\prev_key1_reg_reg[31] [7]));
  LUT5 #(
    .INIT(32'h45664466)) 
    \block_w2_reg[31]_i_1__0 
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(p_0_in[0]),
        .I3(update_type__0[1]),
        .I4(p_0_in[1]),
        .O(block_w2_we));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[31]_i_2 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[31]_i_6_n_0 ),
        .I3(enc_new_block[63]),
        .I4(round_key[63]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[31]));
  LUT2 #(
    .INIT(4'hB)) 
    \block_w2_reg[31]_i_20 
       (.I0(\round_ctr_reg_reg[1]_1 ),
        .I1(muxed_round_nr[2]),
        .O(\round_ctr_reg_reg[1]_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w2_reg[31]_i_22 
       (.I0(enc_round_nr[1]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [1]),
        .O(\round_ctr_reg_reg[1]_3 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w2_reg[31]_i_23 
       (.I0(enc_round_nr[0]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [0]),
        .O(\round_ctr_reg_reg[0]_1 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w2_reg[31]_i_24 
       (.I0(enc_new_block[95]),
        .I1(enc_new_block[127]),
        .I2(enc_new_block[31]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[63]),
        .O(muxed_sboxw__0[31]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    \block_w2_reg[31]_i_25 
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[30]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[30]),
        .I5(init_state),
        .O(\prev_key1_reg_reg[31] [6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w2_reg[31]_i_26 
       (.I0(enc_round_nr[1]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [1]),
        .O(\round_ctr_reg_reg[1]_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w2_reg[31]_i_27 
       (.I0(enc_round_nr[0]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [0]),
        .O(\round_ctr_reg_reg[0]_2 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w2_reg[31]_i_28 
       (.I0(enc_new_block[94]),
        .I1(enc_new_block[126]),
        .I2(enc_new_block[30]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[62]),
        .O(muxed_sboxw__0[30]));
  LUT6 #(
    .INIT(64'h80A8000000000000)) 
    \block_w2_reg[31]_i_3 
       (.I0(enc_ctrl_reg),
        .I1(enc_round_nr[1]),
        .I2(enc_round_nr[2]),
        .I3(p_1_in[3]),
        .I4(enc_round_nr[3]),
        .I5(round_ctr_inc),
        .O(ready_new));
  LUT6 #(
    .INIT(64'h2AAA222AAAAAAAAA)) 
    \block_w2_reg[31]_i_4__0 
       (.I0(round_ctr_inc),
        .I1(enc_ctrl_reg),
        .I2(enc_round_nr[1]),
        .I3(enc_round_nr[2]),
        .I4(p_1_in[3]),
        .I5(enc_round_nr[3]),
        .O(update_type__0[0]));
  LUT6 #(
    .INIT(64'h2A2AAA2AAA2AAAAA)) 
    \block_w2_reg[31]_i_5__0 
       (.I0(enc_ctrl_reg),
        .I1(round_ctr_inc),
        .I2(enc_round_nr[3]),
        .I3(p_1_in[3]),
        .I4(enc_round_nr[2]),
        .I5(enc_round_nr[1]),
        .O(update_type__0[1]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[31]_i_6 
       (.I0(mixcolumns_return044_out[7]),
        .I1(new_sboxw[31]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[39]),
        .I5(round_key[63]),
        .O(\block_w2_reg[31]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \block_w2_reg[31]_i_8 
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(update_type__0[1]),
        .O(\block_w2_reg[31]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[31]_i_9 
       (.I0(enc_new_block[62]),
        .I1(enc_new_block[22]),
        .I2(enc_new_block[111]),
        .I3(enc_new_block[71]),
        .I4(enc_new_block[23]),
        .O(mixcolumns_return044_out[7]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[3]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[3]_i_2_n_0 ),
        .I3(enc_new_block[67]),
        .I4(round_key[35]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[3]));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w2_reg[3]_i_2 
       (.I0(addroundkey0_return__514[35]),
        .I1(new_sboxw[3]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[4]),
        .O(\block_w2_reg[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[3]_i_4 
       (.I0(\block_w2_reg[28]_i_10_n_0 ),
        .I1(\block_w2_reg[4]_i_4__0_n_0 ),
        .I2(enc_new_block[66]),
        .I3(round_key[35]),
        .I4(enc_new_block[58]),
        .I5(enc_new_block[107]),
        .O(addroundkey0_return__514[35]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[4]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[4]_i_2_n_0 ),
        .I3(enc_new_block[68]),
        .I4(round_key[36]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[4]));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w2_reg[4]_i_2 
       (.I0(\block_w2_reg[4]_i_4__0_n_0 ),
        .I1(\block_w2_reg[4]_i_5_n_0 ),
        .I2(new_sboxw[4]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[5]),
        .O(\block_w2_reg[4]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[4]_i_4__0 
       (.I0(enc_new_block[63]),
        .I1(enc_new_block[71]),
        .O(\block_w2_reg[4]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[4]_i_5 
       (.I0(enc_new_block[67]),
        .I1(enc_new_block[108]),
        .I2(enc_new_block[59]),
        .I3(round_key[36]),
        .I4(enc_new_block[60]),
        .I5(enc_new_block[20]),
        .O(\block_w2_reg[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[5]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[5]_i_2_n_0 ),
        .I3(enc_new_block[69]),
        .I4(round_key[37]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[5]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[5]_i_2 
       (.I0(mixcolumns_return034_out[5]),
        .I1(new_sboxw[5]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[22]),
        .I5(round_key[37]),
        .O(\block_w2_reg[5]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[5]_i_4__0 
       (.I0(enc_new_block[109]),
        .I1(enc_new_block[60]),
        .I2(enc_new_block[61]),
        .I3(enc_new_block[21]),
        .I4(enc_new_block[68]),
        .O(mixcolumns_return034_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[6]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[6]_i_2_n_0 ),
        .I3(enc_new_block[70]),
        .I4(round_key[38]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[6]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[6]_i_2 
       (.I0(mixcolumns_return034_out[6]),
        .I1(new_sboxw[6]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[23]),
        .I5(round_key[38]),
        .O(\block_w2_reg[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[6]_i_4__0 
       (.I0(enc_new_block[110]),
        .I1(enc_new_block[61]),
        .I2(enc_new_block[62]),
        .I3(enc_new_block[22]),
        .I4(enc_new_block[69]),
        .O(mixcolumns_return034_out[6]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[7]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[7]_i_2_n_0 ),
        .I3(enc_new_block[71]),
        .I4(round_key[39]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[7]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w2_reg[7]_i_13 
       (.I0(enc_new_block[71]),
        .I1(enc_new_block[103]),
        .I2(enc_new_block[7]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[39]),
        .O(muxed_sboxw__0[7]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    \block_w2_reg[7]_i_14 
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[6]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[6]),
        .I5(init_state),
        .O(\prev_key1_reg_reg[31] [0]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \block_w2_reg[7]_i_15 
       (.I0(enc_new_block[70]),
        .I1(enc_new_block[102]),
        .I2(enc_new_block[6]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[38]),
        .O(muxed_sboxw__0[6]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[7]_i_2 
       (.I0(mixcolumns_return034_out[7]),
        .I1(new_sboxw[7]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[24]),
        .I5(round_key[39]),
        .O(\block_w2_reg[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[7]_i_4__0 
       (.I0(enc_new_block[111]),
        .I1(enc_new_block[62]),
        .I2(enc_new_block[63]),
        .I3(enc_new_block[23]),
        .I4(enc_new_block[70]),
        .O(mixcolumns_return034_out[7]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    \block_w2_reg[7]_i_9 
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[7]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[7]),
        .I5(init_state),
        .O(\prev_key1_reg_reg[31] [1]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[8]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[8]_i_2_n_0 ),
        .I3(enc_new_block[104]),
        .I4(round_key[40]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[8]));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w2_reg[8]_i_2 
       (.I0(mixcolumns_return038_out[0]),
        .I1(new_sboxw[8]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[25]),
        .I5(round_key[40]),
        .O(\block_w2_reg[8]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[8]_i_4__0 
       (.I0(enc_new_block[111]),
        .I1(enc_new_block[64]),
        .I2(enc_new_block[56]),
        .I3(enc_new_block[16]),
        .I4(enc_new_block[71]),
        .O(mixcolumns_return038_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w2_reg[9]_i_1__0 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w2_reg[9]_i_2__0_n_0 ),
        .I3(enc_new_block[105]),
        .I4(round_key[41]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(p_0_in__0[9]));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w2_reg[9]_i_2__0 
       (.I0(\block_w2_reg[9]_i_4__0_n_0 ),
        .I1(\block_w2_reg[9]_i_5__0_n_0 ),
        .I2(new_sboxw[9]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(addroundkey_return[9]),
        .O(\block_w2_reg[9]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[9]_i_4__0 
       (.I0(enc_new_block[111]),
        .I1(enc_new_block[71]),
        .O(\block_w2_reg[9]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[9]_i_5__0 
       (.I0(enc_new_block[104]),
        .I1(enc_new_block[65]),
        .I2(enc_new_block[17]),
        .I3(round_key[41]),
        .I4(enc_new_block[64]),
        .I5(enc_new_block[57]),
        .O(\block_w2_reg[9]_i_5__0_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[0] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[0]),
        .Q(enc_new_block[32]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[10] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[10]),
        .Q(enc_new_block[42]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[11] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[11]),
        .Q(enc_new_block[43]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[12] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[12]),
        .Q(enc_new_block[44]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[13] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[13]),
        .Q(enc_new_block[45]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[14] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[14]),
        .Q(enc_new_block[46]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[15] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[15]),
        .Q(enc_new_block[47]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[16] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[16]),
        .Q(enc_new_block[48]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[17] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[17]),
        .Q(enc_new_block[49]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[18] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[18]),
        .Q(enc_new_block[50]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[19] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[19]),
        .Q(enc_new_block[51]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[1] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[1]),
        .Q(enc_new_block[33]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[20] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[20]),
        .Q(enc_new_block[52]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[21] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[21]),
        .Q(enc_new_block[53]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[22] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[22]),
        .Q(enc_new_block[54]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[23] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[23]),
        .Q(enc_new_block[55]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[24] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[24]),
        .Q(enc_new_block[56]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[25] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[25]),
        .Q(enc_new_block[57]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[26] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[26]),
        .Q(enc_new_block[58]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[27] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[27]),
        .Q(enc_new_block[59]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[28] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[28]),
        .Q(enc_new_block[60]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[29] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[29]),
        .Q(enc_new_block[61]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[2] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[2]),
        .Q(enc_new_block[34]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[30] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[30]),
        .Q(enc_new_block[62]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[31] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[31]),
        .Q(enc_new_block[63]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[3] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[3]),
        .Q(enc_new_block[35]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[4] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[4]),
        .Q(enc_new_block[36]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[5] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[5]),
        .Q(enc_new_block[37]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[6] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[6]),
        .Q(enc_new_block[38]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[7] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[7]),
        .Q(enc_new_block[39]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[8] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[8]),
        .Q(enc_new_block[40]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w2_reg_reg[9] 
       (.C(clk_i),
        .CE(block_w2_we),
        .CLR(rst_i),
        .D(p_0_in__0[9]),
        .Q(enc_new_block[41]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[0]_i_1__0 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[0]_i_2_n_0 ),
        .I3(enc_new_block[32]),
        .I4(round_key[0]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[0]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[0]_i_2 
       (.I0(mixcolumns_return0[0]),
        .I1(new_sboxw[0]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[0]),
        .I5(round_key[0]),
        .O(\block_w3_reg[0]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[0]_i_4__0 
       (.I0(enc_new_block[39]),
        .I1(enc_new_block[72]),
        .I2(enc_new_block[112]),
        .I3(enc_new_block[24]),
        .I4(enc_new_block[31]),
        .O(mixcolumns_return0[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[10]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[10]_i_2_n_0 ),
        .I3(enc_new_block[74]),
        .I4(round_key[10]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[10]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[10]_i_2 
       (.I0(mixcolumns_return022_out[2]),
        .I1(new_sboxw[10]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[6]),
        .I5(round_key[10]),
        .O(\block_w3_reg[10]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[10]_i_4__0 
       (.I0(enc_new_block[73]),
        .I1(enc_new_block[34]),
        .I2(enc_new_block[114]),
        .I3(enc_new_block[26]),
        .I4(enc_new_block[33]),
        .O(mixcolumns_return022_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[11]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[11]_i_2_n_0 ),
        .I3(enc_new_block[75]),
        .I4(round_key[11]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[11]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w3_reg[11]_i_2 
       (.I0(addroundkey0_return__514[11]),
        .I1(new_sboxw[11]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(addroundkey_return[4]),
        .O(\block_w3_reg[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[11]_i_4 
       (.I0(\block_w3_reg[28]_i_9__0_n_0 ),
        .I1(\block_w3_reg[9]_i_4__0_n_0 ),
        .I2(enc_new_block[34]),
        .I3(round_key[11]),
        .I4(enc_new_block[74]),
        .I5(enc_new_block[35]),
        .O(addroundkey0_return__514[11]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[12]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[12]_i_2_n_0 ),
        .I3(enc_new_block[76]),
        .I4(round_key[12]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[12]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w3_reg[12]_i_2 
       (.I0(addroundkey0_return__514[12]),
        .I1(new_sboxw[12]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(addroundkey_return[5]),
        .O(\block_w3_reg[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[12]_i_4 
       (.I0(\block_w3_reg[19]_i_9__0_n_0 ),
        .I1(\block_w3_reg[9]_i_4__0_n_0 ),
        .I2(enc_new_block[28]),
        .I3(round_key[12]),
        .I4(enc_new_block[36]),
        .I5(enc_new_block[116]),
        .O(addroundkey0_return__514[12]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[13]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[13]_i_2_n_0 ),
        .I3(enc_new_block[77]),
        .I4(round_key[13]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[13]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[13]_i_2 
       (.I0(mixcolumns_return022_out[5]),
        .I1(new_sboxw[13]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[7]),
        .I5(round_key[13]),
        .O(\block_w3_reg[13]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[13]_i_4__0 
       (.I0(enc_new_block[76]),
        .I1(enc_new_block[37]),
        .I2(enc_new_block[117]),
        .I3(enc_new_block[29]),
        .I4(enc_new_block[36]),
        .O(mixcolumns_return022_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[14]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[14]_i_2_n_0 ),
        .I3(enc_new_block[78]),
        .I4(round_key[14]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[14]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[14]_i_2 
       (.I0(mixcolumns_return022_out[6]),
        .I1(new_sboxw[14]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[8]),
        .I5(round_key[14]),
        .O(\block_w3_reg[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[14]_i_4__0 
       (.I0(enc_new_block[77]),
        .I1(enc_new_block[38]),
        .I2(enc_new_block[118]),
        .I3(enc_new_block[30]),
        .I4(enc_new_block[37]),
        .O(mixcolumns_return022_out[6]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[15]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[15]_i_2_n_0 ),
        .I3(enc_new_block[79]),
        .I4(round_key[15]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[15]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[15]_i_2 
       (.I0(mixcolumns_return022_out[7]),
        .I1(new_sboxw[15]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[9]),
        .I5(round_key[15]),
        .O(\block_w3_reg[15]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[15]_i_4__0 
       (.I0(enc_new_block[78]),
        .I1(enc_new_block[39]),
        .I2(enc_new_block[119]),
        .I3(enc_new_block[31]),
        .I4(enc_new_block[38]),
        .O(mixcolumns_return022_out[7]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[16]_i_1__0 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[16]_i_2_n_0 ),
        .I3(enc_new_block[112]),
        .I4(round_key[16]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[16]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[16]_i_2 
       (.I0(mixcolumns_return025_out[0]),
        .I1(new_sboxw[16]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[10]),
        .I5(round_key[16]),
        .O(\block_w3_reg[16]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[16]_i_4__0 
       (.I0(enc_new_block[79]),
        .I1(enc_new_block[24]),
        .I2(enc_new_block[72]),
        .I3(enc_new_block[32]),
        .I4(enc_new_block[119]),
        .O(mixcolumns_return025_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[17]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[17]_i_2_n_0 ),
        .I3(enc_new_block[113]),
        .I4(round_key[17]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[17]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w3_reg[17]_i_2 
       (.I0(\block_w3_reg[20]_i_4__0_n_0 ),
        .I1(\block_w3_reg[17]_i_4_n_0 ),
        .I2(new_sboxw[17]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(addroundkey_return[6]),
        .O(\block_w3_reg[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[17]_i_4 
       (.I0(enc_new_block[33]),
        .I1(enc_new_block[112]),
        .I2(enc_new_block[25]),
        .I3(round_key[17]),
        .I4(enc_new_block[72]),
        .I5(enc_new_block[73]),
        .O(\block_w3_reg[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[18]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[18]_i_2_n_0 ),
        .I3(enc_new_block[114]),
        .I4(round_key[18]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[18]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[18]_i_2 
       (.I0(mixcolumns_return025_out[2]),
        .I1(new_sboxw[18]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[11]),
        .I5(round_key[18]),
        .O(\block_w3_reg[18]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[18]_i_4__0 
       (.I0(enc_new_block[73]),
        .I1(enc_new_block[26]),
        .I2(enc_new_block[74]),
        .I3(enc_new_block[34]),
        .I4(enc_new_block[113]),
        .O(mixcolumns_return025_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[19]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[19]_i_2_n_0 ),
        .I3(enc_new_block[115]),
        .I4(round_key[19]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[19]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w3_reg[19]_i_2 
       (.I0(addroundkey0_return__514[19]),
        .I1(new_sboxw[19]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(addroundkey_return[7]),
        .O(\block_w3_reg[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[19]_i_4 
       (.I0(\block_w3_reg[20]_i_4__0_n_0 ),
        .I1(\block_w3_reg[19]_i_9__0_n_0 ),
        .I2(enc_new_block[27]),
        .I3(round_key[19]),
        .I4(enc_new_block[114]),
        .I5(enc_new_block[74]),
        .O(addroundkey0_return__514[19]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[19]_i_9__0 
       (.I0(enc_new_block[35]),
        .I1(enc_new_block[75]),
        .O(\block_w3_reg[19]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[1]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[1]_i_2_n_0 ),
        .I3(enc_new_block[33]),
        .I4(round_key[1]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w3_reg[1]_i_2 
       (.I0(\block_w3_reg[4]_i_4__0_n_0 ),
        .I1(\block_w3_reg[1]_i_4_n_0 ),
        .I2(new_sboxw[1]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(addroundkey_return[0]),
        .O(\block_w3_reg[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[1]_i_4 
       (.I0(enc_new_block[32]),
        .I1(enc_new_block[73]),
        .I2(enc_new_block[25]),
        .I3(round_key[1]),
        .I4(enc_new_block[24]),
        .I5(enc_new_block[113]),
        .O(\block_w3_reg[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[20]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[20]_i_2_n_0 ),
        .I3(enc_new_block[116]),
        .I4(round_key[20]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[20]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w3_reg[20]_i_2 
       (.I0(\block_w3_reg[20]_i_4__0_n_0 ),
        .I1(\block_w3_reg[20]_i_5_n_0 ),
        .I2(new_sboxw[20]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(addroundkey_return[8]),
        .O(\block_w3_reg[20]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[20]_i_4__0 
       (.I0(enc_new_block[119]),
        .I1(enc_new_block[79]),
        .O(\block_w3_reg[20]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[20]_i_5 
       (.I0(enc_new_block[76]),
        .I1(enc_new_block[36]),
        .I2(enc_new_block[115]),
        .I3(round_key[20]),
        .I4(enc_new_block[28]),
        .I5(enc_new_block[75]),
        .O(\block_w3_reg[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[21]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[21]_i_2_n_0 ),
        .I3(enc_new_block[117]),
        .I4(round_key[21]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[21]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[21]_i_2 
       (.I0(mixcolumns_return025_out[5]),
        .I1(new_sboxw[21]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[12]),
        .I5(round_key[21]),
        .O(\block_w3_reg[21]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[21]_i_4__0 
       (.I0(enc_new_block[76]),
        .I1(enc_new_block[29]),
        .I2(enc_new_block[77]),
        .I3(enc_new_block[37]),
        .I4(enc_new_block[116]),
        .O(mixcolumns_return025_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[22]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[22]_i_2_n_0 ),
        .I3(enc_new_block[118]),
        .I4(round_key[22]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[22]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[22]_i_2 
       (.I0(mixcolumns_return025_out[6]),
        .I1(new_sboxw[22]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[13]),
        .I5(round_key[22]),
        .O(\block_w3_reg[22]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[22]_i_4__0 
       (.I0(enc_new_block[77]),
        .I1(enc_new_block[30]),
        .I2(enc_new_block[78]),
        .I3(enc_new_block[38]),
        .I4(enc_new_block[117]),
        .O(mixcolumns_return025_out[6]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[23]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[23]_i_2_n_0 ),
        .I3(enc_new_block[119]),
        .I4(round_key[23]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[23]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[23]_i_2 
       (.I0(mixcolumns_return025_out[7]),
        .I1(new_sboxw[23]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[14]),
        .I5(round_key[23]),
        .O(\block_w3_reg[23]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[23]_i_4__0 
       (.I0(enc_new_block[78]),
        .I1(enc_new_block[31]),
        .I2(enc_new_block[79]),
        .I3(enc_new_block[39]),
        .I4(enc_new_block[118]),
        .O(mixcolumns_return025_out[7]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[24]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[24]_i_2_n_0 ),
        .I3(enc_new_block[24]),
        .I4(round_key[24]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[24]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[24]_i_2 
       (.I0(mixcolumns_return028_out[0]),
        .I1(new_sboxw[24]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[15]),
        .I5(round_key[24]),
        .O(\block_w3_reg[24]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[24]_i_4__0 
       (.I0(enc_new_block[119]),
        .I1(enc_new_block[112]),
        .I2(enc_new_block[72]),
        .I3(enc_new_block[32]),
        .I4(enc_new_block[31]),
        .O(mixcolumns_return028_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[25]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[25]_i_2_n_0 ),
        .I3(enc_new_block[25]),
        .I4(round_key[25]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[25]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w3_reg[25]_i_2 
       (.I0(\block_w3_reg[25]_i_4__0_n_0 ),
        .I1(\block_w3_reg[25]_i_5_n_0 ),
        .I2(new_sboxw[25]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(p_0_out[0]),
        .O(\block_w3_reg[25]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[25]_i_4__0 
       (.I0(enc_new_block[119]),
        .I1(enc_new_block[31]),
        .O(\block_w3_reg[25]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[25]_i_5 
       (.I0(enc_new_block[33]),
        .I1(enc_new_block[112]),
        .I2(enc_new_block[113]),
        .I3(round_key[25]),
        .I4(enc_new_block[73]),
        .I5(enc_new_block[24]),
        .O(\block_w3_reg[25]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w3_reg[25]_i_8 
       (.I0(enc_round_nr[3]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [3]),
        .O(muxed_round_nr[3]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[26]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[26]_i_2_n_0 ),
        .I3(enc_new_block[26]),
        .I4(round_key[26]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[26]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[26]_i_2 
       (.I0(mixcolumns_return028_out[2]),
        .I1(new_sboxw[26]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[16]),
        .I5(round_key[26]),
        .O(\block_w3_reg[26]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[26]_i_4__0 
       (.I0(enc_new_block[113]),
        .I1(enc_new_block[114]),
        .I2(enc_new_block[74]),
        .I3(enc_new_block[34]),
        .I4(enc_new_block[25]),
        .O(mixcolumns_return028_out[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[27]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[27]_i_2_n_0 ),
        .I3(enc_new_block[27]),
        .I4(round_key[27]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[27]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w3_reg[27]_i_2 
       (.I0(addroundkey0_return__514[27]),
        .I1(new_sboxw[27]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[1]),
        .O(\block_w3_reg[27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[27]_i_4 
       (.I0(enc_new_block[35]),
        .I1(enc_new_block[75]),
        .I2(\block_w3_reg[25]_i_4__0_n_0 ),
        .I3(enc_new_block[115]),
        .I4(round_key[27]),
        .I5(\block_w3_reg[27]_i_9__0_n_0 ),
        .O(addroundkey0_return__514[27]));
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[27]_i_9__0 
       (.I0(enc_new_block[114]),
        .I1(enc_new_block[26]),
        .O(\block_w3_reg[27]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[28]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[28]_i_2_n_0 ),
        .I3(enc_new_block[28]),
        .I4(round_key[28]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[28]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w3_reg[28]_i_2 
       (.I0(addroundkey0_return__514[28]),
        .I1(new_sboxw[28]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(p_0_out[2]),
        .O(\block_w3_reg[28]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[28]_i_4 
       (.I0(\block_w3_reg[28]_i_9__0_n_0 ),
        .I1(\block_w3_reg[25]_i_4__0_n_0 ),
        .I2(enc_new_block[116]),
        .I3(round_key[28]),
        .I4(enc_new_block[36]),
        .I5(enc_new_block[76]),
        .O(addroundkey0_return__514[28]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[28]_i_9__0 
       (.I0(enc_new_block[115]),
        .I1(enc_new_block[27]),
        .O(\block_w3_reg[28]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[29]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[29]_i_2_n_0 ),
        .I3(enc_new_block[29]),
        .I4(round_key[29]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[29]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[29]_i_2 
       (.I0(mixcolumns_return028_out[5]),
        .I1(new_sboxw[29]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[17]),
        .I5(round_key[29]),
        .O(\block_w3_reg[29]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[29]_i_4__0 
       (.I0(enc_new_block[116]),
        .I1(enc_new_block[117]),
        .I2(enc_new_block[77]),
        .I3(enc_new_block[37]),
        .I4(enc_new_block[28]),
        .O(mixcolumns_return028_out[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[2]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[2]_i_2_n_0 ),
        .I3(enc_new_block[34]),
        .I4(round_key[2]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[2]_i_2 
       (.I0(mixcolumns_return0[2]),
        .I1(new_sboxw[2]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[1]),
        .I5(round_key[2]),
        .O(\block_w3_reg[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[2]_i_4__0 
       (.I0(enc_new_block[33]),
        .I1(enc_new_block[74]),
        .I2(enc_new_block[114]),
        .I3(enc_new_block[26]),
        .I4(enc_new_block[25]),
        .O(mixcolumns_return0[2]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[30]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[30]_i_2_n_0 ),
        .I3(enc_new_block[30]),
        .I4(round_key[30]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[30]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[30]_i_2 
       (.I0(mixcolumns_return028_out[6]),
        .I1(new_sboxw[30]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[18]),
        .I5(round_key[30]),
        .O(\block_w3_reg[30]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[30]_i_4__0 
       (.I0(enc_new_block[117]),
        .I1(enc_new_block[118]),
        .I2(enc_new_block[78]),
        .I3(enc_new_block[38]),
        .I4(enc_new_block[29]),
        .O(mixcolumns_return028_out[6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w3_reg[31]_i_10 
       (.I0(enc_round_nr[1]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [1]),
        .O(\round_ctr_reg_reg[1]_4 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \block_w3_reg[31]_i_11 
       (.I0(enc_round_nr[0]),
        .I1(p_1_in[2]),
        .I2(\block_w2_reg[28]_i_3 [0]),
        .O(\round_ctr_reg_reg[0]_3 ));
  LUT5 #(
    .INIT(32'h54446666)) 
    \block_w3_reg[31]_i_1__0 
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(p_0_in[1]),
        .I3(p_0_in[0]),
        .I4(update_type__0[1]),
        .O(block_w3_we));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[31]_i_2 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[31]_i_3_n_0 ),
        .I3(enc_new_block[31]),
        .I4(round_key[31]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[31]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[31]_i_3 
       (.I0(mixcolumns_return028_out[7]),
        .I1(new_sboxw[31]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[19]),
        .I5(round_key[31]),
        .O(\block_w3_reg[31]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[31]_i_5__0 
       (.I0(enc_new_block[118]),
        .I1(enc_new_block[119]),
        .I2(enc_new_block[79]),
        .I3(enc_new_block[39]),
        .I4(enc_new_block[30]),
        .O(mixcolumns_return028_out[7]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[3]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[3]_i_2_n_0 ),
        .I3(enc_new_block[35]),
        .I4(round_key[3]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[3]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \block_w3_reg[3]_i_2 
       (.I0(addroundkey0_return__514[3]),
        .I1(new_sboxw[3]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(addroundkey_return[1]),
        .O(\block_w3_reg[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[3]_i_4 
       (.I0(\block_w3_reg[28]_i_9__0_n_0 ),
        .I1(\block_w3_reg[4]_i_4__0_n_0 ),
        .I2(enc_new_block[26]),
        .I3(round_key[3]),
        .I4(enc_new_block[75]),
        .I5(enc_new_block[34]),
        .O(addroundkey0_return__514[3]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[4]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[4]_i_2_n_0 ),
        .I3(enc_new_block[36]),
        .I4(round_key[4]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w3_reg[4]_i_2 
       (.I0(\block_w3_reg[4]_i_4__0_n_0 ),
        .I1(\block_w3_reg[4]_i_5_n_0 ),
        .I2(new_sboxw[4]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(addroundkey_return[2]),
        .O(\block_w3_reg[4]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[4]_i_4__0 
       (.I0(enc_new_block[39]),
        .I1(enc_new_block[31]),
        .O(\block_w3_reg[4]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[4]_i_5 
       (.I0(enc_new_block[35]),
        .I1(enc_new_block[76]),
        .I2(enc_new_block[27]),
        .I3(round_key[4]),
        .I4(enc_new_block[116]),
        .I5(enc_new_block[28]),
        .O(\block_w3_reg[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[5]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[5]_i_2_n_0 ),
        .I3(enc_new_block[37]),
        .I4(round_key[5]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[5]_i_2 
       (.I0(mixcolumns_return0[5]),
        .I1(new_sboxw[5]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[2]),
        .I5(round_key[5]),
        .O(\block_w3_reg[5]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[5]_i_4__0 
       (.I0(enc_new_block[36]),
        .I1(enc_new_block[77]),
        .I2(enc_new_block[117]),
        .I3(enc_new_block[29]),
        .I4(enc_new_block[28]),
        .O(mixcolumns_return0[5]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[6]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[6]_i_2_n_0 ),
        .I3(enc_new_block[38]),
        .I4(round_key[6]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[6]_i_2 
       (.I0(mixcolumns_return0[6]),
        .I1(new_sboxw[6]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[3]),
        .I5(round_key[6]),
        .O(\block_w3_reg[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[6]_i_4__0 
       (.I0(enc_new_block[37]),
        .I1(enc_new_block[78]),
        .I2(enc_new_block[118]),
        .I3(enc_new_block[30]),
        .I4(enc_new_block[29]),
        .O(mixcolumns_return0[6]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[7]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[7]_i_2_n_0 ),
        .I3(enc_new_block[39]),
        .I4(round_key[7]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[7]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[7]_i_2 
       (.I0(mixcolumns_return0[7]),
        .I1(new_sboxw[7]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[4]),
        .I5(round_key[7]),
        .O(\block_w3_reg[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[7]_i_4__0 
       (.I0(enc_new_block[38]),
        .I1(enc_new_block[79]),
        .I2(enc_new_block[119]),
        .I3(enc_new_block[31]),
        .I4(enc_new_block[30]),
        .O(mixcolumns_return0[7]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[8]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[8]_i_2_n_0 ),
        .I3(enc_new_block[72]),
        .I4(round_key[8]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[8]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h50C05FC0AFC0A0C0)) 
    \block_w3_reg[8]_i_2 
       (.I0(mixcolumns_return022_out[0]),
        .I1(new_sboxw[8]),
        .I2(update_type__0[1]),
        .I3(update_type__0[0]),
        .I4(core_block[5]),
        .I5(round_key[8]),
        .O(\block_w3_reg[8]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[8]_i_4__0 
       (.I0(enc_new_block[79]),
        .I1(enc_new_block[32]),
        .I2(enc_new_block[112]),
        .I3(enc_new_block[24]),
        .I4(enc_new_block[39]),
        .O(mixcolumns_return022_out[0]));
  LUT6 #(
    .INIT(64'hB0B0B0B000444400)) 
    \block_w3_reg[9]_i_1 
       (.I0(update_type__0[1]),
        .I1(ready_new),
        .I2(\block_w3_reg[9]_i_2_n_0 ),
        .I3(enc_new_block[73]),
        .I4(round_key[9]),
        .I5(\block_w2_reg[31]_i_8_n_0 ),
        .O(\block_w3_reg[9]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h66FFF0006600F000)) 
    \block_w3_reg[9]_i_2 
       (.I0(\block_w3_reg[9]_i_4__0_n_0 ),
        .I1(\block_w3_reg[9]_i_5_n_0 ),
        .I2(new_sboxw[9]),
        .I3(update_type__0[1]),
        .I4(update_type__0[0]),
        .I5(addroundkey_return[3]),
        .O(\block_w3_reg[9]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[9]_i_4__0 
       (.I0(enc_new_block[79]),
        .I1(enc_new_block[39]),
        .O(\block_w3_reg[9]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[9]_i_5 
       (.I0(enc_new_block[72]),
        .I1(enc_new_block[33]),
        .I2(enc_new_block[25]),
        .I3(round_key[9]),
        .I4(enc_new_block[32]),
        .I5(enc_new_block[113]),
        .O(\block_w3_reg[9]_i_5_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[0] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[0]_i_1__0_n_0 ),
        .Q(enc_new_block[0]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[10] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[10]_i_1_n_0 ),
        .Q(enc_new_block[10]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[11] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[11]_i_1_n_0 ),
        .Q(enc_new_block[11]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[12] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[12]_i_1_n_0 ),
        .Q(enc_new_block[12]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[13] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[13]_i_1_n_0 ),
        .Q(enc_new_block[13]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[14] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[14]_i_1_n_0 ),
        .Q(enc_new_block[14]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[15] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[15]_i_1_n_0 ),
        .Q(enc_new_block[15]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[16] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[16]_i_1__0_n_0 ),
        .Q(enc_new_block[16]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[17] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[17]_i_1_n_0 ),
        .Q(enc_new_block[17]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[18] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[18]_i_1_n_0 ),
        .Q(enc_new_block[18]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[19] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[19]_i_1_n_0 ),
        .Q(enc_new_block[19]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[1] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[1]_i_1_n_0 ),
        .Q(enc_new_block[1]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[20] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[20]_i_1_n_0 ),
        .Q(enc_new_block[20]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[21] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[21]_i_1_n_0 ),
        .Q(enc_new_block[21]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[22] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[22]_i_1_n_0 ),
        .Q(enc_new_block[22]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[23] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[23]_i_1_n_0 ),
        .Q(enc_new_block[23]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[24] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[24]_i_1_n_0 ),
        .Q(enc_new_block[24]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[25] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[25]_i_1_n_0 ),
        .Q(enc_new_block[25]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[26] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[26]_i_1_n_0 ),
        .Q(enc_new_block[26]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[27] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[27]_i_1_n_0 ),
        .Q(enc_new_block[27]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[28] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[28]_i_1_n_0 ),
        .Q(enc_new_block[28]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[29] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[29]_i_1_n_0 ),
        .Q(enc_new_block[29]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[2] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[2]_i_1_n_0 ),
        .Q(enc_new_block[2]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[30] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[30]_i_1_n_0 ),
        .Q(enc_new_block[30]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[31] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[31]_i_2_n_0 ),
        .Q(enc_new_block[31]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[3] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[3]_i_1_n_0 ),
        .Q(enc_new_block[3]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[4] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[4]_i_1_n_0 ),
        .Q(enc_new_block[4]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[5] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[5]_i_1_n_0 ),
        .Q(enc_new_block[5]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[6] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[6]_i_1_n_0 ),
        .Q(enc_new_block[6]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[7] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[7]_i_1_n_0 ),
        .Q(enc_new_block[7]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[8] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[8]_i_1_n_0 ),
        .Q(enc_new_block[8]));
  FDCE #(
    .INIT(1'b0)) 
    \block_w3_reg_reg[9] 
       (.C(clk_i),
        .CE(block_w3_we),
        .CLR(rst_i),
        .D(\block_w3_reg[9]_i_1_n_0 ),
        .Q(enc_new_block[9]));
  LUT6 #(
    .INIT(64'hB14EDE67096C6EED)) 
    g0_b0__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0] ));
  LUT6 #(
    .INIT(64'hB14EDE67096C6EED)) 
    g0_b0__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8] ));
  LUT6 #(
    .INIT(64'hB14EDE67096C6EED)) 
    g0_b0__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16] ));
  LUT6 #(
    .INIT(64'hB14EDE67096C6EED)) 
    g0_b0__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24] ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_10__3
       (.I0(enc_new_block[66]),
        .I1(enc_new_block[98]),
        .I2(enc_new_block[2]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[34]),
        .O(muxed_sboxw__0[2]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_10__4
       (.I0(enc_new_block[75]),
        .I1(enc_new_block[107]),
        .I2(enc_new_block[11]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[43]),
        .O(muxed_sboxw__0[11]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_10__5
       (.I0(enc_new_block[83]),
        .I1(enc_new_block[115]),
        .I2(enc_new_block[19]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[51]),
        .O(muxed_sboxw__0[19]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_10__6
       (.I0(enc_new_block[91]),
        .I1(enc_new_block[123]),
        .I2(enc_new_block[27]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[59]),
        .O(muxed_sboxw__0[27]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_11__3
       (.I0(enc_new_block[67]),
        .I1(enc_new_block[99]),
        .I2(enc_new_block[3]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[35]),
        .O(muxed_sboxw__0[3]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_11__4
       (.I0(enc_new_block[76]),
        .I1(enc_new_block[108]),
        .I2(enc_new_block[12]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[44]),
        .O(muxed_sboxw__0[12]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_11__5
       (.I0(enc_new_block[84]),
        .I1(enc_new_block[116]),
        .I2(enc_new_block[20]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[52]),
        .O(muxed_sboxw__0[20]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_11__6
       (.I0(enc_new_block[92]),
        .I1(enc_new_block[124]),
        .I2(enc_new_block[28]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[60]),
        .O(muxed_sboxw__0[28]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_12__3
       (.I0(enc_new_block[68]),
        .I1(enc_new_block[100]),
        .I2(enc_new_block[4]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[36]),
        .O(muxed_sboxw__0[4]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_12__4
       (.I0(enc_new_block[77]),
        .I1(enc_new_block[109]),
        .I2(enc_new_block[13]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[45]),
        .O(muxed_sboxw__0[13]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_12__5
       (.I0(enc_new_block[85]),
        .I1(enc_new_block[117]),
        .I2(enc_new_block[21]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[53]),
        .O(muxed_sboxw__0[21]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_12__6
       (.I0(enc_new_block[93]),
        .I1(enc_new_block[125]),
        .I2(enc_new_block[29]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[61]),
        .O(muxed_sboxw__0[29]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_13__0
       (.I0(enc_new_block[69]),
        .I1(enc_new_block[101]),
        .I2(enc_new_block[5]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[37]),
        .O(muxed_sboxw__0[5]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_1__3
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[24]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[24]),
        .I5(init_state),
        .O(muxed_sboxw[24]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_1__4
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[16]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[16]),
        .I5(init_state),
        .O(muxed_sboxw[16]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_1__5
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[8]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[8]),
        .I5(init_state),
        .O(muxed_sboxw[8]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_1__6
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[0]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[0]),
        .I5(init_state),
        .O(muxed_sboxw[0]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_2__3
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[25]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[25]),
        .I5(init_state),
        .O(muxed_sboxw[25]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_2__4
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[17]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[17]),
        .I5(init_state),
        .O(muxed_sboxw[17]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_2__5
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[9]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[9]),
        .I5(init_state),
        .O(muxed_sboxw[9]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_2__6
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[1]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[1]),
        .I5(init_state),
        .O(muxed_sboxw[1]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_3__3
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[26]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[26]),
        .I5(init_state),
        .O(muxed_sboxw[26]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_3__4
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[18]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[18]),
        .I5(init_state),
        .O(muxed_sboxw[18]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_3__5
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[10]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[10]),
        .I5(init_state),
        .O(muxed_sboxw[10]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_3__6
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[2]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[2]),
        .I5(init_state),
        .O(muxed_sboxw[2]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_4__3
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[27]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[27]),
        .I5(init_state),
        .O(muxed_sboxw[27]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_4__4
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[19]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[19]),
        .I5(init_state),
        .O(muxed_sboxw[19]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_4__5
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[11]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[11]),
        .I5(init_state),
        .O(muxed_sboxw[11]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_4__6
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[3]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[3]),
        .I5(init_state),
        .O(muxed_sboxw[3]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_5__3
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[28]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[28]),
        .I5(init_state),
        .O(muxed_sboxw[28]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_5__4
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[20]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[20]),
        .I5(init_state),
        .O(muxed_sboxw[20]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_5__5
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[12]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[12]),
        .I5(init_state),
        .O(muxed_sboxw[12]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_5__6
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[4]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[4]),
        .I5(init_state),
        .O(muxed_sboxw[4]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_6__3
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[29]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[29]),
        .I5(init_state),
        .O(muxed_sboxw[29]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_6__4
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[21]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[21]),
        .I5(init_state),
        .O(muxed_sboxw[21]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_6__5
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[13]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[13]),
        .I5(init_state),
        .O(muxed_sboxw[13]));
  LUT6 #(
    .INIT(64'hF0F0F0F011000000)) 
    g0_b0_i_6__6
       (.I0(ready_new),
        .I1(update_type__0[0]),
        .I2(Q[5]),
        .I3(update_type__0[1]),
        .I4(muxed_sboxw__0[5]),
        .I5(init_state),
        .O(muxed_sboxw[5]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_7__3
       (.I0(enc_new_block[64]),
        .I1(enc_new_block[96]),
        .I2(enc_new_block[0]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[32]),
        .O(muxed_sboxw__0[0]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_7__4
       (.I0(enc_new_block[72]),
        .I1(enc_new_block[104]),
        .I2(enc_new_block[8]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[40]),
        .O(muxed_sboxw__0[8]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_7__5
       (.I0(enc_new_block[80]),
        .I1(enc_new_block[112]),
        .I2(enc_new_block[16]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[48]),
        .O(muxed_sboxw__0[16]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_7__6
       (.I0(enc_new_block[88]),
        .I1(enc_new_block[120]),
        .I2(enc_new_block[24]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[56]),
        .O(muxed_sboxw__0[24]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_8__3
       (.I0(enc_new_block[73]),
        .I1(enc_new_block[105]),
        .I2(enc_new_block[9]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[41]),
        .O(muxed_sboxw__0[9]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_8__4
       (.I0(enc_new_block[81]),
        .I1(enc_new_block[113]),
        .I2(enc_new_block[17]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[49]),
        .O(muxed_sboxw__0[17]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_8__5
       (.I0(enc_new_block[89]),
        .I1(enc_new_block[121]),
        .I2(enc_new_block[25]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[57]),
        .O(muxed_sboxw__0[25]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_9__3
       (.I0(enc_new_block[65]),
        .I1(enc_new_block[97]),
        .I2(enc_new_block[1]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[33]),
        .O(muxed_sboxw__0[1]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_9__4
       (.I0(enc_new_block[74]),
        .I1(enc_new_block[106]),
        .I2(enc_new_block[10]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[42]),
        .O(muxed_sboxw__0[10]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_9__5
       (.I0(enc_new_block[82]),
        .I1(enc_new_block[114]),
        .I2(enc_new_block[18]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[50]),
        .O(muxed_sboxw__0[18]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    g0_b0_i_9__6
       (.I0(enc_new_block[90]),
        .I1(enc_new_block[122]),
        .I2(enc_new_block[26]),
        .I3(p_0_in[1]),
        .I4(p_0_in[0]),
        .I5(enc_new_block[58]),
        .O(muxed_sboxw__0[26]));
  LUT6 #(
    .INIT(64'h7BAE007D4C53FC7D)) 
    g0_b1__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h7BAE007D4C53FC7D)) 
    g0_b1__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h7BAE007D4C53FC7D)) 
    g0_b1__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_0 ));
  LUT6 #(
    .INIT(64'h7BAE007D4C53FC7D)) 
    g0_b1__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_0 ));
  LUT6 #(
    .INIT(64'hA16387FB3B48B4C6)) 
    g0_b2__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_1 ));
  LUT6 #(
    .INIT(64'hA16387FB3B48B4C6)) 
    g0_b2__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_1 ));
  LUT6 #(
    .INIT(64'hA16387FB3B48B4C6)) 
    g0_b2__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_1 ));
  LUT6 #(
    .INIT(64'hA16387FB3B48B4C6)) 
    g0_b2__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_1 ));
  LUT6 #(
    .INIT(64'h109020A2193D586A)) 
    g0_b3__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_2 ));
  LUT6 #(
    .INIT(64'h109020A2193D586A)) 
    g0_b3__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_2 ));
  LUT6 #(
    .INIT(64'h109020A2193D586A)) 
    g0_b3__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_2 ));
  LUT6 #(
    .INIT(64'h109020A2193D586A)) 
    g0_b3__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_2 ));
  LUT6 #(
    .INIT(64'hC2B0F97752B8B11E)) 
    g0_b4__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_3 ));
  LUT6 #(
    .INIT(64'hC2B0F97752B8B11E)) 
    g0_b4__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_3 ));
  LUT6 #(
    .INIT(64'hC2B0F97752B8B11E)) 
    g0_b4__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_3 ));
  LUT6 #(
    .INIT(64'hC2B0F97752B8B11E)) 
    g0_b4__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_3 ));
  LUT6 #(
    .INIT(64'hF8045F7B6D98DD7F)) 
    g0_b5__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_4 ));
  LUT6 #(
    .INIT(64'hF8045F7B6D98DD7F)) 
    g0_b5__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_4 ));
  LUT6 #(
    .INIT(64'hF8045F7B6D98DD7F)) 
    g0_b5__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_4 ));
  LUT6 #(
    .INIT(64'hF8045F7B6D98DD7F)) 
    g0_b5__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_4 ));
  LUT6 #(
    .INIT(64'h980A3CC2C2FDB4FF)) 
    g0_b6__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_5 ));
  LUT6 #(
    .INIT(64'h980A3CC2C2FDB4FF)) 
    g0_b6__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_5 ));
  LUT6 #(
    .INIT(64'h980A3CC2C2FDB4FF)) 
    g0_b6__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_5 ));
  LUT6 #(
    .INIT(64'h980A3CC2C2FDB4FF)) 
    g0_b6__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_5 ));
  LUT6 #(
    .INIT(64'h5CAA2EC7BF977090)) 
    g0_b7__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_6 ));
  LUT6 #(
    .INIT(64'h5CAA2EC7BF977090)) 
    g0_b7__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_6 ));
  LUT6 #(
    .INIT(64'h5CAA2EC7BF977090)) 
    g0_b7__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_6 ));
  LUT6 #(
    .INIT(64'h5CAA2EC7BF977090)) 
    g0_b7__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_6 ));
  LUT6 #(
    .INIT(64'h68AB4BFA8ACB7A13)) 
    g1_b0__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_7 ));
  LUT6 #(
    .INIT(64'h68AB4BFA8ACB7A13)) 
    g1_b0__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_7 ));
  LUT6 #(
    .INIT(64'h68AB4BFA8ACB7A13)) 
    g1_b0__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_7 ));
  LUT6 #(
    .INIT(64'h68AB4BFA8ACB7A13)) 
    g1_b0__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_7 ));
  LUT6 #(
    .INIT(64'hE61A4C5E97816F7A)) 
    g1_b1__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_8 ));
  LUT6 #(
    .INIT(64'hE61A4C5E97816F7A)) 
    g1_b1__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_8 ));
  LUT6 #(
    .INIT(64'hE61A4C5E97816F7A)) 
    g1_b1__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_8 ));
  LUT6 #(
    .INIT(64'hE61A4C5E97816F7A)) 
    g1_b1__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_8 ));
  LUT6 #(
    .INIT(64'h23A869A2A428C424)) 
    g1_b2__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_9 ));
  LUT6 #(
    .INIT(64'h23A869A2A428C424)) 
    g1_b2__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_9 ));
  LUT6 #(
    .INIT(64'h23A869A2A428C424)) 
    g1_b2__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_9 ));
  LUT6 #(
    .INIT(64'h23A869A2A428C424)) 
    g1_b2__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_9 ));
  LUT6 #(
    .INIT(64'h2568EA2EFFA8527D)) 
    g1_b3__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_10 ));
  LUT6 #(
    .INIT(64'h2568EA2EFFA8527D)) 
    g1_b3__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_10 ));
  LUT6 #(
    .INIT(64'h2568EA2EFFA8527D)) 
    g1_b3__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_10 ));
  LUT6 #(
    .INIT(64'h2568EA2EFFA8527D)) 
    g1_b3__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_10 ));
  LUT6 #(
    .INIT(64'hF7F17A494CE30F58)) 
    g1_b4__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_11 ));
  LUT6 #(
    .INIT(64'hF7F17A494CE30F58)) 
    g1_b4__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_11 ));
  LUT6 #(
    .INIT(64'hF7F17A494CE30F58)) 
    g1_b4__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_11 ));
  LUT6 #(
    .INIT(64'hF7F17A494CE30F58)) 
    g1_b4__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_11 ));
  LUT6 #(
    .INIT(64'h6BC2AA4E0D787AA4)) 
    g1_b5__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_12 ));
  LUT6 #(
    .INIT(64'h6BC2AA4E0D787AA4)) 
    g1_b5__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_12 ));
  LUT6 #(
    .INIT(64'h6BC2AA4E0D787AA4)) 
    g1_b5__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_12 ));
  LUT6 #(
    .INIT(64'h6BC2AA4E0D787AA4)) 
    g1_b5__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_12 ));
  LUT6 #(
    .INIT(64'hE4851B3BF3AB2560)) 
    g1_b6__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_13 ));
  LUT6 #(
    .INIT(64'hE4851B3BF3AB2560)) 
    g1_b6__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_13 ));
  LUT6 #(
    .INIT(64'hE4851B3BF3AB2560)) 
    g1_b6__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_13 ));
  LUT6 #(
    .INIT(64'hE4851B3BF3AB2560)) 
    g1_b6__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_13 ));
  LUT6 #(
    .INIT(64'hE7BAC28F866AAC82)) 
    g1_b7__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_14 ));
  LUT6 #(
    .INIT(64'hE7BAC28F866AAC82)) 
    g1_b7__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_14 ));
  LUT6 #(
    .INIT(64'hE7BAC28F866AAC82)) 
    g1_b7__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_14 ));
  LUT6 #(
    .INIT(64'hE7BAC28F866AAC82)) 
    g1_b7__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_14 ));
  LUT6 #(
    .INIT(64'h10BDB210C006EAB5)) 
    g2_b0__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_15 ));
  LUT6 #(
    .INIT(64'h10BDB210C006EAB5)) 
    g2_b0__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_15 ));
  LUT6 #(
    .INIT(64'h10BDB210C006EAB5)) 
    g2_b0__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_15 ));
  LUT6 #(
    .INIT(64'h10BDB210C006EAB5)) 
    g2_b0__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_15 ));
  LUT6 #(
    .INIT(64'h6A450B2EF33486B4)) 
    g2_b1__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_16 ));
  LUT6 #(
    .INIT(64'h6A450B2EF33486B4)) 
    g2_b1__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_16 ));
  LUT6 #(
    .INIT(64'h6A450B2EF33486B4)) 
    g2_b1__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_16 ));
  LUT6 #(
    .INIT(64'h6A450B2EF33486B4)) 
    g2_b1__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_16 ));
  LUT6 #(
    .INIT(64'h577D64E03B0C3FFB)) 
    g2_b2__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_17 ));
  LUT6 #(
    .INIT(64'h577D64E03B0C3FFB)) 
    g2_b2__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_17 ));
  LUT6 #(
    .INIT(64'h577D64E03B0C3FFB)) 
    g2_b2__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_17 ));
  LUT6 #(
    .INIT(64'h577D64E03B0C3FFB)) 
    g2_b2__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_17 ));
  LUT6 #(
    .INIT(64'hE9DA849CF6AC6C1B)) 
    g2_b3__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_18 ));
  LUT6 #(
    .INIT(64'hE9DA849CF6AC6C1B)) 
    g2_b3__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_18 ));
  LUT6 #(
    .INIT(64'hE9DA849CF6AC6C1B)) 
    g2_b3__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_18 ));
  LUT6 #(
    .INIT(64'hE9DA849CF6AC6C1B)) 
    g2_b3__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_18 ));
  LUT6 #(
    .INIT(64'h2624B286BC48ECB4)) 
    g2_b4__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_19 ));
  LUT6 #(
    .INIT(64'h2624B286BC48ECB4)) 
    g2_b4__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_19 ));
  LUT6 #(
    .INIT(64'h2624B286BC48ECB4)) 
    g2_b4__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_19 ));
  LUT6 #(
    .INIT(64'h2624B286BC48ECB4)) 
    g2_b4__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_19 ));
  LUT6 #(
    .INIT(64'h7D8DCC4706319E08)) 
    g2_b5__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_20 ));
  LUT6 #(
    .INIT(64'h7D8DCC4706319E08)) 
    g2_b5__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_20 ));
  LUT6 #(
    .INIT(64'h7D8DCC4706319E08)) 
    g2_b5__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_20 ));
  LUT6 #(
    .INIT(64'h7D8DCC4706319E08)) 
    g2_b5__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_20 ));
  LUT6 #(
    .INIT(64'h3F6BCB91B30DB559)) 
    g2_b6__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_21 ));
  LUT6 #(
    .INIT(64'h3F6BCB91B30DB559)) 
    g2_b6__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_21 ));
  LUT6 #(
    .INIT(64'h3F6BCB91B30DB559)) 
    g2_b6__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_21 ));
  LUT6 #(
    .INIT(64'h3F6BCB91B30DB559)) 
    g2_b6__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_21 ));
  LUT6 #(
    .INIT(64'h4CB3770196CA0329)) 
    g2_b7__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_22 ));
  LUT6 #(
    .INIT(64'h4CB3770196CA0329)) 
    g2_b7__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_22 ));
  LUT6 #(
    .INIT(64'h4CB3770196CA0329)) 
    g2_b7__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_22 ));
  LUT6 #(
    .INIT(64'h4CB3770196CA0329)) 
    g2_b7__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_22 ));
  LUT6 #(
    .INIT(64'h4F1EAD396F247A04)) 
    g3_b0__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_23 ));
  LUT6 #(
    .INIT(64'h4F1EAD396F247A04)) 
    g3_b0__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_23 ));
  LUT6 #(
    .INIT(64'h4F1EAD396F247A04)) 
    g3_b0__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_23 ));
  LUT6 #(
    .INIT(64'h4F1EAD396F247A04)) 
    g3_b0__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_23 ));
  LUT6 #(
    .INIT(64'hC870974094EAD8A9)) 
    g3_b1__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_24 ));
  LUT6 #(
    .INIT(64'hC870974094EAD8A9)) 
    g3_b1__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_24 ));
  LUT6 #(
    .INIT(64'hC870974094EAD8A9)) 
    g3_b1__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_24 ));
  LUT6 #(
    .INIT(64'hC870974094EAD8A9)) 
    g3_b1__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_24 ));
  LUT6 #(
    .INIT(64'hAC39B6C0D6CE2EFC)) 
    g3_b2__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_25 ));
  LUT6 #(
    .INIT(64'hAC39B6C0D6CE2EFC)) 
    g3_b2__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_25 ));
  LUT6 #(
    .INIT(64'hAC39B6C0D6CE2EFC)) 
    g3_b2__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_25 ));
  LUT6 #(
    .INIT(64'hAC39B6C0D6CE2EFC)) 
    g3_b2__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_25 ));
  LUT6 #(
    .INIT(64'h4E9DDB76C892FB1B)) 
    g3_b3__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_26 ));
  LUT6 #(
    .INIT(64'h4E9DDB76C892FB1B)) 
    g3_b3__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_26 ));
  LUT6 #(
    .INIT(64'h4E9DDB76C892FB1B)) 
    g3_b3__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_26 ));
  LUT6 #(
    .INIT(64'h4E9DDB76C892FB1B)) 
    g3_b3__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_26 ));
  LUT6 #(
    .INIT(64'hF210A3AECE472E53)) 
    g3_b4__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_27 ));
  LUT6 #(
    .INIT(64'hF210A3AECE472E53)) 
    g3_b4__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_27 ));
  LUT6 #(
    .INIT(64'hF210A3AECE472E53)) 
    g3_b4__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_27 ));
  LUT6 #(
    .INIT(64'hF210A3AECE472E53)) 
    g3_b4__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_27 ));
  LUT6 #(
    .INIT(64'h54B248130B4F256F)) 
    g3_b5__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_28 ));
  LUT6 #(
    .INIT(64'h54B248130B4F256F)) 
    g3_b5__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_28 ));
  LUT6 #(
    .INIT(64'h54B248130B4F256F)) 
    g3_b5__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_28 ));
  LUT6 #(
    .INIT(64'h54B248130B4F256F)) 
    g3_b5__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_28 ));
  LUT6 #(
    .INIT(64'h21E0B83325591782)) 
    g3_b6__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_29 ));
  LUT6 #(
    .INIT(64'h21E0B83325591782)) 
    g3_b6__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_29 ));
  LUT6 #(
    .INIT(64'h21E0B83325591782)) 
    g3_b6__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_29 ));
  LUT6 #(
    .INIT(64'h21E0B83325591782)) 
    g3_b6__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_29 ));
  LUT6 #(
    .INIT(64'h52379DE7B844E3E1)) 
    g3_b7__3
       (.I0(muxed_sboxw[0]),
        .I1(muxed_sboxw[1]),
        .I2(muxed_sboxw[2]),
        .I3(muxed_sboxw[3]),
        .I4(muxed_sboxw[4]),
        .I5(muxed_sboxw[5]),
        .O(\prev_key1_reg_reg[0]_30 ));
  LUT6 #(
    .INIT(64'h52379DE7B844E3E1)) 
    g3_b7__4
       (.I0(muxed_sboxw[8]),
        .I1(muxed_sboxw[9]),
        .I2(muxed_sboxw[10]),
        .I3(muxed_sboxw[11]),
        .I4(muxed_sboxw[12]),
        .I5(muxed_sboxw[13]),
        .O(\prev_key1_reg_reg[8]_30 ));
  LUT6 #(
    .INIT(64'h52379DE7B844E3E1)) 
    g3_b7__5
       (.I0(muxed_sboxw[16]),
        .I1(muxed_sboxw[17]),
        .I2(muxed_sboxw[18]),
        .I3(muxed_sboxw[19]),
        .I4(muxed_sboxw[20]),
        .I5(muxed_sboxw[21]),
        .O(\prev_key1_reg_reg[16]_30 ));
  LUT6 #(
    .INIT(64'h52379DE7B844E3E1)) 
    g3_b7__6
       (.I0(muxed_sboxw[24]),
        .I1(muxed_sboxw[25]),
        .I2(muxed_sboxw[26]),
        .I3(muxed_sboxw[27]),
        .I4(muxed_sboxw[28]),
        .I5(muxed_sboxw[29]),
        .O(\prev_key1_reg_reg[24]_30 ));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[120]_i_4 
       (.I0(new_sboxw[16]),
        .I1(\prev_key1_reg[127]_i_5 [0]),
        .O(p_19_in[0]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[121]_i_4 
       (.I0(new_sboxw[17]),
        .I1(\prev_key1_reg[127]_i_5 [1]),
        .O(p_19_in[1]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[122]_i_4 
       (.I0(new_sboxw[18]),
        .I1(\prev_key1_reg[127]_i_5 [2]),
        .O(p_19_in[2]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[123]_i_4 
       (.I0(new_sboxw[19]),
        .I1(\prev_key1_reg[127]_i_5 [3]),
        .O(p_19_in[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[124]_i_4 
       (.I0(new_sboxw[20]),
        .I1(\prev_key1_reg[127]_i_5 [4]),
        .O(p_19_in[4]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[125]_i_4 
       (.I0(new_sboxw[21]),
        .I1(\prev_key1_reg[127]_i_5 [5]),
        .O(p_19_in[5]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[126]_i_4 
       (.I0(new_sboxw[22]),
        .I1(\prev_key1_reg[127]_i_5 [6]),
        .O(p_19_in[6]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[127]_i_6 
       (.I0(new_sboxw[23]),
        .I1(\prev_key1_reg[127]_i_5 [7]),
        .O(p_19_in[7]));
  LUT6 #(
    .INIT(64'hFFFFCFFF44440000)) 
    ready_reg_i_1
       (.I0(ready_reg_i_2__0_n_0),
        .I1(round_ctr_inc),
        .I2(p_1_in[1]),
        .I3(p_1_in[2]),
        .I4(enc_ctrl_reg),
        .I5(enc_ready),
        .O(ready_reg_i_1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT4 #(
    .INIT(16'h71FF)) 
    ready_reg_i_2__0
       (.I0(enc_round_nr[1]),
        .I1(enc_round_nr[2]),
        .I2(p_1_in[3]),
        .I3(enc_round_nr[3]),
        .O(ready_reg_i_2__0_n_0));
  FDPE #(
    .INIT(1'b1)) 
    ready_reg_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(ready_reg_i_1_n_0),
        .PRE(rst_i),
        .Q(enc_ready));
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[0]_i_1 
       (.I0(enc_new_block[0]),
        .I1(dec_new_block[0]),
        .I2(p_1_in[2]),
        .O(D[0]));
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[100]_i_1 
       (.I0(enc_new_block[100]),
        .I1(dec_new_block[100]),
        .I2(p_1_in[2]),
        .O(D[100]));
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[101]_i_1 
       (.I0(enc_new_block[101]),
        .I1(dec_new_block[101]),
        .I2(p_1_in[2]),
        .O(D[101]));
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[102]_i_1 
       (.I0(enc_new_block[102]),
        .I1(dec_new_block[102]),
        .I2(p_1_in[2]),
        .O(D[102]));
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[103]_i_1 
       (.I0(enc_new_block[103]),
        .I1(dec_new_block[103]),
        .I2(p_1_in[2]),
        .O(D[103]));
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[104]_i_1 
       (.I0(enc_new_block[104]),
        .I1(dec_new_block[104]),
        .I2(p_1_in[2]),
        .O(D[104]));
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[105]_i_1 
       (.I0(enc_new_block[105]),
        .I1(dec_new_block[105]),
        .I2(p_1_in[2]),
        .O(D[105]));
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[106]_i_1 
       (.I0(enc_new_block[106]),
        .I1(dec_new_block[106]),
        .I2(p_1_in[2]),
        .O(D[106]));
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[107]_i_1 
       (.I0(enc_new_block[107]),
        .I1(dec_new_block[107]),
        .I2(p_1_in[2]),
        .O(D[107]));
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[108]_i_1 
       (.I0(enc_new_block[108]),
        .I1(dec_new_block[108]),
        .I2(p_1_in[2]),
        .O(D[108]));
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[109]_i_1 
       (.I0(enc_new_block[109]),
        .I1(dec_new_block[109]),
        .I2(p_1_in[2]),
        .O(D[109]));
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[10]_i_1 
       (.I0(enc_new_block[10]),
        .I1(dec_new_block[10]),
        .I2(p_1_in[2]),
        .O(D[10]));
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[110]_i_1 
       (.I0(enc_new_block[110]),
        .I1(dec_new_block[110]),
        .I2(p_1_in[2]),
        .O(D[110]));
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[111]_i_1 
       (.I0(enc_new_block[111]),
        .I1(dec_new_block[111]),
        .I2(p_1_in[2]),
        .O(D[111]));
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[112]_i_1 
       (.I0(enc_new_block[112]),
        .I1(dec_new_block[112]),
        .I2(p_1_in[2]),
        .O(D[112]));
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[113]_i_1 
       (.I0(enc_new_block[113]),
        .I1(dec_new_block[113]),
        .I2(p_1_in[2]),
        .O(D[113]));
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[114]_i_1 
       (.I0(enc_new_block[114]),
        .I1(dec_new_block[114]),
        .I2(p_1_in[2]),
        .O(D[114]));
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[115]_i_1 
       (.I0(enc_new_block[115]),
        .I1(dec_new_block[115]),
        .I2(p_1_in[2]),
        .O(D[115]));
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[116]_i_1 
       (.I0(enc_new_block[116]),
        .I1(dec_new_block[116]),
        .I2(p_1_in[2]),
        .O(D[116]));
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[117]_i_1 
       (.I0(enc_new_block[117]),
        .I1(dec_new_block[117]),
        .I2(p_1_in[2]),
        .O(D[117]));
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[118]_i_1 
       (.I0(enc_new_block[118]),
        .I1(dec_new_block[118]),
        .I2(p_1_in[2]),
        .O(D[118]));
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[119]_i_1 
       (.I0(enc_new_block[119]),
        .I1(dec_new_block[119]),
        .I2(p_1_in[2]),
        .O(D[119]));
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[11]_i_1 
       (.I0(enc_new_block[11]),
        .I1(dec_new_block[11]),
        .I2(p_1_in[2]),
        .O(D[11]));
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[120]_i_1 
       (.I0(enc_new_block[120]),
        .I1(dec_new_block[120]),
        .I2(p_1_in[2]),
        .O(D[120]));
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[121]_i_1 
       (.I0(enc_new_block[121]),
        .I1(dec_new_block[121]),
        .I2(p_1_in[2]),
        .O(D[121]));
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[122]_i_1 
       (.I0(enc_new_block[122]),
        .I1(dec_new_block[122]),
        .I2(p_1_in[2]),
        .O(D[122]));
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[123]_i_1 
       (.I0(enc_new_block[123]),
        .I1(dec_new_block[123]),
        .I2(p_1_in[2]),
        .O(D[123]));
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[124]_i_1 
       (.I0(enc_new_block[124]),
        .I1(dec_new_block[124]),
        .I2(p_1_in[2]),
        .O(D[124]));
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[125]_i_1 
       (.I0(enc_new_block[125]),
        .I1(dec_new_block[125]),
        .I2(p_1_in[2]),
        .O(D[125]));
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[126]_i_1 
       (.I0(enc_new_block[126]),
        .I1(dec_new_block[126]),
        .I2(p_1_in[2]),
        .O(D[126]));
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[127]_i_1 
       (.I0(enc_new_block[127]),
        .I1(dec_new_block[127]),
        .I2(p_1_in[2]),
        .O(D[127]));
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[12]_i_1 
       (.I0(enc_new_block[12]),
        .I1(dec_new_block[12]),
        .I2(p_1_in[2]),
        .O(D[12]));
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[13]_i_1 
       (.I0(enc_new_block[13]),
        .I1(dec_new_block[13]),
        .I2(p_1_in[2]),
        .O(D[13]));
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[14]_i_1 
       (.I0(enc_new_block[14]),
        .I1(dec_new_block[14]),
        .I2(p_1_in[2]),
        .O(D[14]));
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[15]_i_1 
       (.I0(enc_new_block[15]),
        .I1(dec_new_block[15]),
        .I2(p_1_in[2]),
        .O(D[15]));
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[16]_i_1 
       (.I0(enc_new_block[16]),
        .I1(dec_new_block[16]),
        .I2(p_1_in[2]),
        .O(D[16]));
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[17]_i_1 
       (.I0(enc_new_block[17]),
        .I1(dec_new_block[17]),
        .I2(p_1_in[2]),
        .O(D[17]));
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[18]_i_1 
       (.I0(enc_new_block[18]),
        .I1(dec_new_block[18]),
        .I2(p_1_in[2]),
        .O(D[18]));
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[19]_i_1 
       (.I0(enc_new_block[19]),
        .I1(dec_new_block[19]),
        .I2(p_1_in[2]),
        .O(D[19]));
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[1]_i_1 
       (.I0(enc_new_block[1]),
        .I1(dec_new_block[1]),
        .I2(p_1_in[2]),
        .O(D[1]));
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[20]_i_1 
       (.I0(enc_new_block[20]),
        .I1(dec_new_block[20]),
        .I2(p_1_in[2]),
        .O(D[20]));
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[21]_i_1 
       (.I0(enc_new_block[21]),
        .I1(dec_new_block[21]),
        .I2(p_1_in[2]),
        .O(D[21]));
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[22]_i_1 
       (.I0(enc_new_block[22]),
        .I1(dec_new_block[22]),
        .I2(p_1_in[2]),
        .O(D[22]));
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[23]_i_1 
       (.I0(enc_new_block[23]),
        .I1(dec_new_block[23]),
        .I2(p_1_in[2]),
        .O(D[23]));
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[24]_i_1 
       (.I0(enc_new_block[24]),
        .I1(dec_new_block[24]),
        .I2(p_1_in[2]),
        .O(D[24]));
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[25]_i_1 
       (.I0(enc_new_block[25]),
        .I1(dec_new_block[25]),
        .I2(p_1_in[2]),
        .O(D[25]));
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[26]_i_1 
       (.I0(enc_new_block[26]),
        .I1(dec_new_block[26]),
        .I2(p_1_in[2]),
        .O(D[26]));
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[27]_i_1 
       (.I0(enc_new_block[27]),
        .I1(dec_new_block[27]),
        .I2(p_1_in[2]),
        .O(D[27]));
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[28]_i_1 
       (.I0(enc_new_block[28]),
        .I1(dec_new_block[28]),
        .I2(p_1_in[2]),
        .O(D[28]));
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[29]_i_1 
       (.I0(enc_new_block[29]),
        .I1(dec_new_block[29]),
        .I2(p_1_in[2]),
        .O(D[29]));
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[2]_i_1 
       (.I0(enc_new_block[2]),
        .I1(dec_new_block[2]),
        .I2(p_1_in[2]),
        .O(D[2]));
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[30]_i_1 
       (.I0(enc_new_block[30]),
        .I1(dec_new_block[30]),
        .I2(p_1_in[2]),
        .O(D[30]));
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[31]_i_1 
       (.I0(enc_new_block[31]),
        .I1(dec_new_block[31]),
        .I2(p_1_in[2]),
        .O(D[31]));
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[32]_i_1 
       (.I0(enc_new_block[32]),
        .I1(dec_new_block[32]),
        .I2(p_1_in[2]),
        .O(D[32]));
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[33]_i_1 
       (.I0(enc_new_block[33]),
        .I1(dec_new_block[33]),
        .I2(p_1_in[2]),
        .O(D[33]));
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[34]_i_1 
       (.I0(enc_new_block[34]),
        .I1(dec_new_block[34]),
        .I2(p_1_in[2]),
        .O(D[34]));
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[35]_i_1 
       (.I0(enc_new_block[35]),
        .I1(dec_new_block[35]),
        .I2(p_1_in[2]),
        .O(D[35]));
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[36]_i_1 
       (.I0(enc_new_block[36]),
        .I1(dec_new_block[36]),
        .I2(p_1_in[2]),
        .O(D[36]));
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[37]_i_1 
       (.I0(enc_new_block[37]),
        .I1(dec_new_block[37]),
        .I2(p_1_in[2]),
        .O(D[37]));
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[38]_i_1 
       (.I0(enc_new_block[38]),
        .I1(dec_new_block[38]),
        .I2(p_1_in[2]),
        .O(D[38]));
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[39]_i_1 
       (.I0(enc_new_block[39]),
        .I1(dec_new_block[39]),
        .I2(p_1_in[2]),
        .O(D[39]));
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[3]_i_1 
       (.I0(enc_new_block[3]),
        .I1(dec_new_block[3]),
        .I2(p_1_in[2]),
        .O(D[3]));
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[40]_i_1 
       (.I0(enc_new_block[40]),
        .I1(dec_new_block[40]),
        .I2(p_1_in[2]),
        .O(D[40]));
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[41]_i_1 
       (.I0(enc_new_block[41]),
        .I1(dec_new_block[41]),
        .I2(p_1_in[2]),
        .O(D[41]));
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[42]_i_1 
       (.I0(enc_new_block[42]),
        .I1(dec_new_block[42]),
        .I2(p_1_in[2]),
        .O(D[42]));
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[43]_i_1 
       (.I0(enc_new_block[43]),
        .I1(dec_new_block[43]),
        .I2(p_1_in[2]),
        .O(D[43]));
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[44]_i_1 
       (.I0(enc_new_block[44]),
        .I1(dec_new_block[44]),
        .I2(p_1_in[2]),
        .O(D[44]));
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[45]_i_1 
       (.I0(enc_new_block[45]),
        .I1(dec_new_block[45]),
        .I2(p_1_in[2]),
        .O(D[45]));
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[46]_i_1 
       (.I0(enc_new_block[46]),
        .I1(dec_new_block[46]),
        .I2(p_1_in[2]),
        .O(D[46]));
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[47]_i_1 
       (.I0(enc_new_block[47]),
        .I1(dec_new_block[47]),
        .I2(p_1_in[2]),
        .O(D[47]));
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[48]_i_1 
       (.I0(enc_new_block[48]),
        .I1(dec_new_block[48]),
        .I2(p_1_in[2]),
        .O(D[48]));
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[49]_i_1 
       (.I0(enc_new_block[49]),
        .I1(dec_new_block[49]),
        .I2(p_1_in[2]),
        .O(D[49]));
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[4]_i_1 
       (.I0(enc_new_block[4]),
        .I1(dec_new_block[4]),
        .I2(p_1_in[2]),
        .O(D[4]));
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[50]_i_1 
       (.I0(enc_new_block[50]),
        .I1(dec_new_block[50]),
        .I2(p_1_in[2]),
        .O(D[50]));
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[51]_i_1 
       (.I0(enc_new_block[51]),
        .I1(dec_new_block[51]),
        .I2(p_1_in[2]),
        .O(D[51]));
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[52]_i_1 
       (.I0(enc_new_block[52]),
        .I1(dec_new_block[52]),
        .I2(p_1_in[2]),
        .O(D[52]));
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[53]_i_1 
       (.I0(enc_new_block[53]),
        .I1(dec_new_block[53]),
        .I2(p_1_in[2]),
        .O(D[53]));
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[54]_i_1 
       (.I0(enc_new_block[54]),
        .I1(dec_new_block[54]),
        .I2(p_1_in[2]),
        .O(D[54]));
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[55]_i_1 
       (.I0(enc_new_block[55]),
        .I1(dec_new_block[55]),
        .I2(p_1_in[2]),
        .O(D[55]));
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[56]_i_1 
       (.I0(enc_new_block[56]),
        .I1(dec_new_block[56]),
        .I2(p_1_in[2]),
        .O(D[56]));
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[57]_i_1 
       (.I0(enc_new_block[57]),
        .I1(dec_new_block[57]),
        .I2(p_1_in[2]),
        .O(D[57]));
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[58]_i_1 
       (.I0(enc_new_block[58]),
        .I1(dec_new_block[58]),
        .I2(p_1_in[2]),
        .O(D[58]));
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[59]_i_1 
       (.I0(enc_new_block[59]),
        .I1(dec_new_block[59]),
        .I2(p_1_in[2]),
        .O(D[59]));
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[5]_i_1 
       (.I0(enc_new_block[5]),
        .I1(dec_new_block[5]),
        .I2(p_1_in[2]),
        .O(D[5]));
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[60]_i_1 
       (.I0(enc_new_block[60]),
        .I1(dec_new_block[60]),
        .I2(p_1_in[2]),
        .O(D[60]));
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[61]_i_1 
       (.I0(enc_new_block[61]),
        .I1(dec_new_block[61]),
        .I2(p_1_in[2]),
        .O(D[61]));
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[62]_i_1 
       (.I0(enc_new_block[62]),
        .I1(dec_new_block[62]),
        .I2(p_1_in[2]),
        .O(D[62]));
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[63]_i_1 
       (.I0(enc_new_block[63]),
        .I1(dec_new_block[63]),
        .I2(p_1_in[2]),
        .O(D[63]));
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[64]_i_1 
       (.I0(enc_new_block[64]),
        .I1(dec_new_block[64]),
        .I2(p_1_in[2]),
        .O(D[64]));
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[65]_i_1 
       (.I0(enc_new_block[65]),
        .I1(dec_new_block[65]),
        .I2(p_1_in[2]),
        .O(D[65]));
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[66]_i_1 
       (.I0(enc_new_block[66]),
        .I1(dec_new_block[66]),
        .I2(p_1_in[2]),
        .O(D[66]));
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[67]_i_1 
       (.I0(enc_new_block[67]),
        .I1(dec_new_block[67]),
        .I2(p_1_in[2]),
        .O(D[67]));
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[68]_i_1 
       (.I0(enc_new_block[68]),
        .I1(dec_new_block[68]),
        .I2(p_1_in[2]),
        .O(D[68]));
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[69]_i_1 
       (.I0(enc_new_block[69]),
        .I1(dec_new_block[69]),
        .I2(p_1_in[2]),
        .O(D[69]));
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[6]_i_1 
       (.I0(enc_new_block[6]),
        .I1(dec_new_block[6]),
        .I2(p_1_in[2]),
        .O(D[6]));
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[70]_i_1 
       (.I0(enc_new_block[70]),
        .I1(dec_new_block[70]),
        .I2(p_1_in[2]),
        .O(D[70]));
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[71]_i_1 
       (.I0(enc_new_block[71]),
        .I1(dec_new_block[71]),
        .I2(p_1_in[2]),
        .O(D[71]));
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[72]_i_1 
       (.I0(enc_new_block[72]),
        .I1(dec_new_block[72]),
        .I2(p_1_in[2]),
        .O(D[72]));
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[73]_i_1 
       (.I0(enc_new_block[73]),
        .I1(dec_new_block[73]),
        .I2(p_1_in[2]),
        .O(D[73]));
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[74]_i_1 
       (.I0(enc_new_block[74]),
        .I1(dec_new_block[74]),
        .I2(p_1_in[2]),
        .O(D[74]));
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[75]_i_1 
       (.I0(enc_new_block[75]),
        .I1(dec_new_block[75]),
        .I2(p_1_in[2]),
        .O(D[75]));
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[76]_i_1 
       (.I0(enc_new_block[76]),
        .I1(dec_new_block[76]),
        .I2(p_1_in[2]),
        .O(D[76]));
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[77]_i_1 
       (.I0(enc_new_block[77]),
        .I1(dec_new_block[77]),
        .I2(p_1_in[2]),
        .O(D[77]));
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[78]_i_1 
       (.I0(enc_new_block[78]),
        .I1(dec_new_block[78]),
        .I2(p_1_in[2]),
        .O(D[78]));
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[79]_i_1 
       (.I0(enc_new_block[79]),
        .I1(dec_new_block[79]),
        .I2(p_1_in[2]),
        .O(D[79]));
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[7]_i_1 
       (.I0(enc_new_block[7]),
        .I1(dec_new_block[7]),
        .I2(p_1_in[2]),
        .O(D[7]));
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[80]_i_1 
       (.I0(enc_new_block[80]),
        .I1(dec_new_block[80]),
        .I2(p_1_in[2]),
        .O(D[80]));
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[81]_i_1 
       (.I0(enc_new_block[81]),
        .I1(dec_new_block[81]),
        .I2(p_1_in[2]),
        .O(D[81]));
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[82]_i_1 
       (.I0(enc_new_block[82]),
        .I1(dec_new_block[82]),
        .I2(p_1_in[2]),
        .O(D[82]));
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[83]_i_1 
       (.I0(enc_new_block[83]),
        .I1(dec_new_block[83]),
        .I2(p_1_in[2]),
        .O(D[83]));
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[84]_i_1 
       (.I0(enc_new_block[84]),
        .I1(dec_new_block[84]),
        .I2(p_1_in[2]),
        .O(D[84]));
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[85]_i_1 
       (.I0(enc_new_block[85]),
        .I1(dec_new_block[85]),
        .I2(p_1_in[2]),
        .O(D[85]));
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[86]_i_1 
       (.I0(enc_new_block[86]),
        .I1(dec_new_block[86]),
        .I2(p_1_in[2]),
        .O(D[86]));
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[87]_i_1 
       (.I0(enc_new_block[87]),
        .I1(dec_new_block[87]),
        .I2(p_1_in[2]),
        .O(D[87]));
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[88]_i_1 
       (.I0(enc_new_block[88]),
        .I1(dec_new_block[88]),
        .I2(p_1_in[2]),
        .O(D[88]));
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[89]_i_1 
       (.I0(enc_new_block[89]),
        .I1(dec_new_block[89]),
        .I2(p_1_in[2]),
        .O(D[89]));
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[8]_i_1 
       (.I0(enc_new_block[8]),
        .I1(dec_new_block[8]),
        .I2(p_1_in[2]),
        .O(D[8]));
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[90]_i_1 
       (.I0(enc_new_block[90]),
        .I1(dec_new_block[90]),
        .I2(p_1_in[2]),
        .O(D[90]));
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[91]_i_1 
       (.I0(enc_new_block[91]),
        .I1(dec_new_block[91]),
        .I2(p_1_in[2]),
        .O(D[91]));
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[92]_i_1 
       (.I0(enc_new_block[92]),
        .I1(dec_new_block[92]),
        .I2(p_1_in[2]),
        .O(D[92]));
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[93]_i_1 
       (.I0(enc_new_block[93]),
        .I1(dec_new_block[93]),
        .I2(p_1_in[2]),
        .O(D[93]));
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[94]_i_1 
       (.I0(enc_new_block[94]),
        .I1(dec_new_block[94]),
        .I2(p_1_in[2]),
        .O(D[94]));
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[95]_i_1 
       (.I0(enc_new_block[95]),
        .I1(dec_new_block[95]),
        .I2(p_1_in[2]),
        .O(D[95]));
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[96]_i_1 
       (.I0(enc_new_block[96]),
        .I1(dec_new_block[96]),
        .I2(p_1_in[2]),
        .O(D[96]));
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[97]_i_1 
       (.I0(enc_new_block[97]),
        .I1(dec_new_block[97]),
        .I2(p_1_in[2]),
        .O(D[97]));
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[98]_i_1 
       (.I0(enc_new_block[98]),
        .I1(dec_new_block[98]),
        .I2(p_1_in[2]),
        .O(D[98]));
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[99]_i_1 
       (.I0(enc_new_block[99]),
        .I1(dec_new_block[99]),
        .I2(p_1_in[2]),
        .O(D[99]));
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \result_reg[9]_i_1 
       (.I0(enc_new_block[9]),
        .I1(dec_new_block[9]),
        .I2(p_1_in[2]),
        .O(D[9]));
  LUT6 #(
    .INIT(64'hFFFFF1F10000F000)) 
    result_valid_reg_i_1
       (.I0(p_1_in[1]),
        .I1(p_1_in[0]),
        .I2(result_valid_reg_reg[1]),
        .I3(muxed_ready),
        .I4(result_valid_reg_reg[0]),
        .I5(core_valid),
        .O(next_reg_reg));
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \round_ctr_reg[0]_i_1__0 
       (.I0(enc_round_nr[0]),
        .I1(round_ctr_inc),
        .O(round_ctr_new[0]));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT3 #(
    .INIT(8'h60)) 
    \round_ctr_reg[1]_i_1__0 
       (.I0(enc_round_nr[0]),
        .I1(enc_round_nr[1]),
        .I2(round_ctr_inc),
        .O(round_ctr_new[1]));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT5 #(
    .INIT(32'h00007800)) 
    \round_ctr_reg[2]_i_1__0 
       (.I0(enc_round_nr[0]),
        .I1(enc_round_nr[1]),
        .I2(enc_round_nr[2]),
        .I3(round_ctr_inc),
        .I4(round_ctr_rst__1),
        .O(round_ctr_new[2]));
  LUT4 #(
    .INIT(16'hFF40)) 
    \round_ctr_reg[3]_i_1__0 
       (.I0(enc_ctrl_reg),
        .I1(p_1_in[2]),
        .I2(p_1_in[1]),
        .I3(round_ctr_inc),
        .O(round_ctr_we));
  LUT6 #(
    .INIT(64'h000000007F800000)) 
    \round_ctr_reg[3]_i_2__0 
       (.I0(enc_round_nr[1]),
        .I1(enc_round_nr[0]),
        .I2(enc_round_nr[2]),
        .I3(enc_round_nr[3]),
        .I4(round_ctr_inc),
        .I5(round_ctr_rst__1),
        .O(round_ctr_new[3]));
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \round_ctr_reg[3]_i_3 
       (.I0(p_1_in[1]),
        .I1(p_1_in[2]),
        .I2(round_ctr_inc),
        .I3(enc_ctrl_reg),
        .O(round_ctr_rst__1));
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[0] 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(round_ctr_new[0]),
        .Q(enc_round_nr[0]));
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[1] 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(round_ctr_new[1]),
        .Q(enc_round_nr[1]));
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[2] 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(round_ctr_new[2]),
        .Q(enc_round_nr[2]));
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[3] 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(round_ctr_new[3]),
        .Q(enc_round_nr[3]));
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \sword_ctr_reg[0]_i_1 
       (.I0(p_0_in[0]),
        .I1(enc_ctrl_reg),
        .I2(round_ctr_inc),
        .O(sword_ctr_new[0]));
  LUT2 #(
    .INIT(4'hE)) 
    \sword_ctr_reg[1]_i_1 
       (.I0(round_ctr_inc),
        .I1(enc_ctrl_reg),
        .O(sword_ctr_we));
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT4 #(
    .INIT(16'h0060)) 
    \sword_ctr_reg[1]_i_2 
       (.I0(p_0_in[0]),
        .I1(p_0_in[1]),
        .I2(enc_ctrl_reg),
        .I3(round_ctr_inc),
        .O(sword_ctr_new[1]));
  FDCE #(
    .INIT(1'b0)) 
    \sword_ctr_reg_reg[0] 
       (.C(clk_i),
        .CE(sword_ctr_we),
        .CLR(rst_i),
        .D(sword_ctr_new[0]),
        .Q(p_0_in[0]));
  FDCE #(
    .INIT(1'b0)) 
    \sword_ctr_reg_reg[1] 
       (.C(clk_i),
        .CE(sword_ctr_we),
        .CLR(rst_i),
        .D(sword_ctr_new[1]),
        .Q(p_0_in[1]));
endmodule

(* ORIG_REF_NAME = "aes_inv_sbox" *) 
module switch_elements_aes_inv_sbox
   (\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11_0 ,
    new_sboxw,
    tmp_sboxw_0,
    \block_w3_reg_reg[0]_i_8_0 ,
    \block_w3_reg_reg[0]_i_8_1 ,
    \block_w3_reg_reg[0]_i_8_2 ,
    \block_w3_reg_reg[0]_i_8_3 ,
    \block_w3_reg_reg[1]_i_5_0 ,
    \block_w3_reg_reg[1]_i_5_1 ,
    \block_w3_reg_reg[1]_i_5_2 ,
    \block_w3_reg_reg[1]_i_5_3 ,
    \block_w3_reg_reg[2]_i_6_0 ,
    \block_w3_reg_reg[2]_i_6_1 ,
    \block_w3_reg_reg[2]_i_6_2 ,
    \block_w3_reg_reg[2]_i_6_3 ,
    \block_w3_reg_reg[3]_i_5_0 ,
    \block_w3_reg_reg[3]_i_5_1 ,
    \block_w3_reg_reg[3]_i_5_2 ,
    \block_w3_reg_reg[3]_i_5_3 ,
    \block_w3_reg_reg[4]_i_5_0 ,
    \block_w3_reg_reg[4]_i_5_1 ,
    \block_w3_reg_reg[4]_i_5_2 ,
    \block_w3_reg_reg[4]_i_5_3 ,
    \block_w3_reg_reg[5]_i_6_0 ,
    \block_w3_reg_reg[5]_i_6_1 ,
    \block_w3_reg_reg[5]_i_6_2 ,
    \block_w3_reg_reg[5]_i_6_3 ,
    \block_w3_reg_reg[6]_i_6_0 ,
    \block_w3_reg_reg[6]_i_6_1 ,
    \block_w3_reg_reg[6]_i_6_2 ,
    \block_w3_reg_reg[6]_i_6_3 ,
    \block_w3_reg_reg[7]_i_6_0 ,
    \block_w3_reg_reg[7]_i_6_1 ,
    \block_w3_reg_reg[7]_i_6_2 ,
    \block_w3_reg_reg[7]_i_6_3 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_0 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_1 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_2 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_3 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_0 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_1 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_2 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_3 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_0 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_1 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_2 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_3 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_0 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_1 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_2 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_3 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_0 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_1 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_2 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_3 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_0 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_1 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_2 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_3 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_0 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_1 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_2 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_3 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_0 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_1 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_2 ,
    \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_3 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_0 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_1 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_2 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_3 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_0 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_1 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_2 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_3 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_0 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_1 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_2 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_3 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_0 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_1 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_2 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_3 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_0 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_1 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_2 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_3 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_0 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_1 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_2 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_3 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_0 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_1 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_2 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_3 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_0 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_1 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_2 ,
    \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_3 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_0 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_1 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_2 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_3 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_0 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_1 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_2 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_3 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_0 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_1 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_2 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_3 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_0 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_1 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_2 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_3 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_0 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_1 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_2 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_3 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_0 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_1 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_2 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_3 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_0 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_1 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_2 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_3 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_0 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_1 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_2 ,
    \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_3 );
  output [2:0]\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11_0 ;
  output [28:0]new_sboxw;
  input [7:0]tmp_sboxw_0;
  input \block_w3_reg_reg[0]_i_8_0 ;
  input \block_w3_reg_reg[0]_i_8_1 ;
  input \block_w3_reg_reg[0]_i_8_2 ;
  input \block_w3_reg_reg[0]_i_8_3 ;
  input \block_w3_reg_reg[1]_i_5_0 ;
  input \block_w3_reg_reg[1]_i_5_1 ;
  input \block_w3_reg_reg[1]_i_5_2 ;
  input \block_w3_reg_reg[1]_i_5_3 ;
  input \block_w3_reg_reg[2]_i_6_0 ;
  input \block_w3_reg_reg[2]_i_6_1 ;
  input \block_w3_reg_reg[2]_i_6_2 ;
  input \block_w3_reg_reg[2]_i_6_3 ;
  input \block_w3_reg_reg[3]_i_5_0 ;
  input \block_w3_reg_reg[3]_i_5_1 ;
  input \block_w3_reg_reg[3]_i_5_2 ;
  input \block_w3_reg_reg[3]_i_5_3 ;
  input \block_w3_reg_reg[4]_i_5_0 ;
  input \block_w3_reg_reg[4]_i_5_1 ;
  input \block_w3_reg_reg[4]_i_5_2 ;
  input \block_w3_reg_reg[4]_i_5_3 ;
  input \block_w3_reg_reg[5]_i_6_0 ;
  input \block_w3_reg_reg[5]_i_6_1 ;
  input \block_w3_reg_reg[5]_i_6_2 ;
  input \block_w3_reg_reg[5]_i_6_3 ;
  input \block_w3_reg_reg[6]_i_6_0 ;
  input \block_w3_reg_reg[6]_i_6_1 ;
  input \block_w3_reg_reg[6]_i_6_2 ;
  input \block_w3_reg_reg[6]_i_6_3 ;
  input \block_w3_reg_reg[7]_i_6_0 ;
  input \block_w3_reg_reg[7]_i_6_1 ;
  input \block_w3_reg_reg[7]_i_6_2 ;
  input \block_w3_reg_reg[7]_i_6_3 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_0 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_1 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_2 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_3 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_0 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_1 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_2 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_3 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_0 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_1 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_2 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_3 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_0 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_1 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_2 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_3 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_0 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_1 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_2 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_3 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_0 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_1 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_2 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_3 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_0 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_1 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_2 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_3 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_0 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_1 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_2 ;
  input \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_3 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_0 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_1 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_2 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_3 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_0 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_1 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_2 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_3 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_0 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_1 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_2 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_3 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_0 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_1 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_2 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_3 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_0 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_1 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_2 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_3 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_0 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_1 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_2 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_3 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_0 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_1 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_2 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_3 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_0 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_1 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_2 ;
  input \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_3 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_0 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_1 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_2 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_3 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_0 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_1 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_2 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_3 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_0 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_1 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_2 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_3 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_0 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_1 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_2 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_3 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_0 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_1 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_2 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_3 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_0 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_1 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_2 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_3 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_0 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_1 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_2 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_3 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_0 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_1 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_2 ;
  input \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_3 ;

  wire \block_w3_reg_reg[0]_i_10_n_0 ;
  wire \block_w3_reg_reg[0]_i_8_0 ;
  wire \block_w3_reg_reg[0]_i_8_1 ;
  wire \block_w3_reg_reg[0]_i_8_2 ;
  wire \block_w3_reg_reg[0]_i_8_3 ;
  wire \block_w3_reg_reg[0]_i_9_n_0 ;
  wire \block_w3_reg_reg[1]_i_5_0 ;
  wire \block_w3_reg_reg[1]_i_5_1 ;
  wire \block_w3_reg_reg[1]_i_5_2 ;
  wire \block_w3_reg_reg[1]_i_5_3 ;
  wire \block_w3_reg_reg[1]_i_7_n_0 ;
  wire \block_w3_reg_reg[1]_i_8_n_0 ;
  wire \block_w3_reg_reg[2]_i_6_0 ;
  wire \block_w3_reg_reg[2]_i_6_1 ;
  wire \block_w3_reg_reg[2]_i_6_2 ;
  wire \block_w3_reg_reg[2]_i_6_3 ;
  wire \block_w3_reg_reg[2]_i_8_n_0 ;
  wire \block_w3_reg_reg[2]_i_9_n_0 ;
  wire \block_w3_reg_reg[3]_i_5_0 ;
  wire \block_w3_reg_reg[3]_i_5_1 ;
  wire \block_w3_reg_reg[3]_i_5_2 ;
  wire \block_w3_reg_reg[3]_i_5_3 ;
  wire \block_w3_reg_reg[3]_i_7_n_0 ;
  wire \block_w3_reg_reg[3]_i_8_n_0 ;
  wire \block_w3_reg_reg[4]_i_5_0 ;
  wire \block_w3_reg_reg[4]_i_5_1 ;
  wire \block_w3_reg_reg[4]_i_5_2 ;
  wire \block_w3_reg_reg[4]_i_5_3 ;
  wire \block_w3_reg_reg[4]_i_7_n_0 ;
  wire \block_w3_reg_reg[4]_i_8_n_0 ;
  wire \block_w3_reg_reg[5]_i_6_0 ;
  wire \block_w3_reg_reg[5]_i_6_1 ;
  wire \block_w3_reg_reg[5]_i_6_2 ;
  wire \block_w3_reg_reg[5]_i_6_3 ;
  wire \block_w3_reg_reg[5]_i_8_n_0 ;
  wire \block_w3_reg_reg[5]_i_9_n_0 ;
  wire \block_w3_reg_reg[6]_i_6_0 ;
  wire \block_w3_reg_reg[6]_i_6_1 ;
  wire \block_w3_reg_reg[6]_i_6_2 ;
  wire \block_w3_reg_reg[6]_i_6_3 ;
  wire \block_w3_reg_reg[6]_i_8_n_0 ;
  wire \block_w3_reg_reg[6]_i_9_n_0 ;
  wire \block_w3_reg_reg[7]_i_10_n_0 ;
  wire \block_w3_reg_reg[7]_i_6_0 ;
  wire \block_w3_reg_reg[7]_i_6_1 ;
  wire \block_w3_reg_reg[7]_i_6_2 ;
  wire \block_w3_reg_reg[7]_i_6_3 ;
  wire \block_w3_reg_reg[7]_i_9_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_1 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_2 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_3 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_8_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_9_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_1 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_2 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_3 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_6_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_7_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_1 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_2 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_3 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_7_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_8_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_1 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_2 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_3 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_8_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_9_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_1 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_2 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_3 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_8_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_9_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_10_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_1 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_2 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_3 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_9_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_1 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_2 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_3 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_8_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_9_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_1 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_2 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_3 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_7_n_0 ;
  wire \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_8_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_10_n_0 ;
  wire [2:0]\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_1 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_2 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_3 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_1 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_2 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_3 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_7_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_8_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_1 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_2 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_3 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_7_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_8_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_1 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_2 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_3 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_7_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_8_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_1 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_2 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_3 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_7_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_8_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_1 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_2 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_3 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_8_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_9_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_1 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_2 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_3 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_8_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_9_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_10_n_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_0 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_1 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_2 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_3 ;
  wire \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_9_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_1 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_2 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_3 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_8_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_9_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_1 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_2 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_3 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_7_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_8_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_1 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_2 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_3 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_7_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_8_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_1 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_2 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_3 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_6_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_7_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_1 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_2 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_3 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_7_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_8_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_1 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_2 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_3 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_8_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_9_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_1 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_2 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_3 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_8_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_9_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_11_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_12_n_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_0 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_1 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_2 ;
  wire \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_3 ;
  wire [28:0]new_sboxw;
  wire [7:0]tmp_sboxw_0;

  MUXF7 \block_w3_reg_reg[0]_i_10 
       (.I0(\block_w3_reg_reg[0]_i_8_2 ),
        .I1(\block_w3_reg_reg[0]_i_8_3 ),
        .O(\block_w3_reg_reg[0]_i_10_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF8 \block_w3_reg_reg[0]_i_8 
       (.I0(\block_w3_reg_reg[0]_i_9_n_0 ),
        .I1(\block_w3_reg_reg[0]_i_10_n_0 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11_0 [0]),
        .S(tmp_sboxw_0[1]));
  MUXF7 \block_w3_reg_reg[0]_i_9 
       (.I0(\block_w3_reg_reg[0]_i_8_0 ),
        .I1(\block_w3_reg_reg[0]_i_8_1 ),
        .O(\block_w3_reg_reg[0]_i_9_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF8 \block_w3_reg_reg[1]_i_5 
       (.I0(\block_w3_reg_reg[1]_i_7_n_0 ),
        .I1(\block_w3_reg_reg[1]_i_8_n_0 ),
        .O(new_sboxw[0]),
        .S(tmp_sboxw_0[1]));
  MUXF7 \block_w3_reg_reg[1]_i_7 
       (.I0(\block_w3_reg_reg[1]_i_5_0 ),
        .I1(\block_w3_reg_reg[1]_i_5_1 ),
        .O(\block_w3_reg_reg[1]_i_7_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF7 \block_w3_reg_reg[1]_i_8 
       (.I0(\block_w3_reg_reg[1]_i_5_2 ),
        .I1(\block_w3_reg_reg[1]_i_5_3 ),
        .O(\block_w3_reg_reg[1]_i_8_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF8 \block_w3_reg_reg[2]_i_6 
       (.I0(\block_w3_reg_reg[2]_i_8_n_0 ),
        .I1(\block_w3_reg_reg[2]_i_9_n_0 ),
        .O(new_sboxw[1]),
        .S(tmp_sboxw_0[1]));
  MUXF7 \block_w3_reg_reg[2]_i_8 
       (.I0(\block_w3_reg_reg[2]_i_6_0 ),
        .I1(\block_w3_reg_reg[2]_i_6_1 ),
        .O(\block_w3_reg_reg[2]_i_8_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF7 \block_w3_reg_reg[2]_i_9 
       (.I0(\block_w3_reg_reg[2]_i_6_2 ),
        .I1(\block_w3_reg_reg[2]_i_6_3 ),
        .O(\block_w3_reg_reg[2]_i_9_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF8 \block_w3_reg_reg[3]_i_5 
       (.I0(\block_w3_reg_reg[3]_i_7_n_0 ),
        .I1(\block_w3_reg_reg[3]_i_8_n_0 ),
        .O(new_sboxw[2]),
        .S(tmp_sboxw_0[1]));
  MUXF7 \block_w3_reg_reg[3]_i_7 
       (.I0(\block_w3_reg_reg[3]_i_5_0 ),
        .I1(\block_w3_reg_reg[3]_i_5_1 ),
        .O(\block_w3_reg_reg[3]_i_7_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF7 \block_w3_reg_reg[3]_i_8 
       (.I0(\block_w3_reg_reg[3]_i_5_2 ),
        .I1(\block_w3_reg_reg[3]_i_5_3 ),
        .O(\block_w3_reg_reg[3]_i_8_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF8 \block_w3_reg_reg[4]_i_5 
       (.I0(\block_w3_reg_reg[4]_i_7_n_0 ),
        .I1(\block_w3_reg_reg[4]_i_8_n_0 ),
        .O(new_sboxw[3]),
        .S(tmp_sboxw_0[1]));
  MUXF7 \block_w3_reg_reg[4]_i_7 
       (.I0(\block_w3_reg_reg[4]_i_5_0 ),
        .I1(\block_w3_reg_reg[4]_i_5_1 ),
        .O(\block_w3_reg_reg[4]_i_7_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF7 \block_w3_reg_reg[4]_i_8 
       (.I0(\block_w3_reg_reg[4]_i_5_2 ),
        .I1(\block_w3_reg_reg[4]_i_5_3 ),
        .O(\block_w3_reg_reg[4]_i_8_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF8 \block_w3_reg_reg[5]_i_6 
       (.I0(\block_w3_reg_reg[5]_i_8_n_0 ),
        .I1(\block_w3_reg_reg[5]_i_9_n_0 ),
        .O(new_sboxw[4]),
        .S(tmp_sboxw_0[1]));
  MUXF7 \block_w3_reg_reg[5]_i_8 
       (.I0(\block_w3_reg_reg[5]_i_6_0 ),
        .I1(\block_w3_reg_reg[5]_i_6_1 ),
        .O(\block_w3_reg_reg[5]_i_8_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF7 \block_w3_reg_reg[5]_i_9 
       (.I0(\block_w3_reg_reg[5]_i_6_2 ),
        .I1(\block_w3_reg_reg[5]_i_6_3 ),
        .O(\block_w3_reg_reg[5]_i_9_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF8 \block_w3_reg_reg[6]_i_6 
       (.I0(\block_w3_reg_reg[6]_i_8_n_0 ),
        .I1(\block_w3_reg_reg[6]_i_9_n_0 ),
        .O(new_sboxw[5]),
        .S(tmp_sboxw_0[1]));
  MUXF7 \block_w3_reg_reg[6]_i_8 
       (.I0(\block_w3_reg_reg[6]_i_6_0 ),
        .I1(\block_w3_reg_reg[6]_i_6_1 ),
        .O(\block_w3_reg_reg[6]_i_8_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF7 \block_w3_reg_reg[6]_i_9 
       (.I0(\block_w3_reg_reg[6]_i_6_2 ),
        .I1(\block_w3_reg_reg[6]_i_6_3 ),
        .O(\block_w3_reg_reg[6]_i_9_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF7 \block_w3_reg_reg[7]_i_10 
       (.I0(\block_w3_reg_reg[7]_i_6_2 ),
        .I1(\block_w3_reg_reg[7]_i_6_3 ),
        .O(\block_w3_reg_reg[7]_i_10_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF8 \block_w3_reg_reg[7]_i_6 
       (.I0(\block_w3_reg_reg[7]_i_9_n_0 ),
        .I1(\block_w3_reg_reg[7]_i_10_n_0 ),
        .O(new_sboxw[6]),
        .S(tmp_sboxw_0[1]));
  MUXF7 \block_w3_reg_reg[7]_i_9 
       (.I0(\block_w3_reg_reg[7]_i_6_0 ),
        .I1(\block_w3_reg_reg[7]_i_6_1 ),
        .O(\block_w3_reg_reg[7]_i_9_n_0 ),
        .S(tmp_sboxw_0[0]));
  MUXF8 \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[10]_i_8_n_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[10]_i_9_n_0 ),
        .O(new_sboxw[8]),
        .S(tmp_sboxw_0[3]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_8 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_1 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[10]_i_8_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[10]_i_9 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_2 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[10]_i_6_3 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[10]_i_9_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF8 \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[11]_i_6_n_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[11]_i_7_n_0 ),
        .O(new_sboxw[9]),
        .S(tmp_sboxw_0[3]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_6 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_1 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[11]_i_6_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[11]_i_7 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_2 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[11]_i_4_3 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[11]_i_7_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF8 \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[12]_i_7_n_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[12]_i_8_n_0 ),
        .O(new_sboxw[10]),
        .S(tmp_sboxw_0[3]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_7 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_1 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[12]_i_7_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[12]_i_8 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_2 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[12]_i_5_3 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[12]_i_8_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF8 \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[13]_i_8_n_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[13]_i_9_n_0 ),
        .O(new_sboxw[11]),
        .S(tmp_sboxw_0[3]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_8 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_1 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[13]_i_8_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[13]_i_9 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_2 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[13]_i_6_3 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[13]_i_9_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF8 \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[14]_i_8_n_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[14]_i_9_n_0 ),
        .O(new_sboxw[12]),
        .S(tmp_sboxw_0[3]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_8 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_1 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[14]_i_8_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[14]_i_9 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_2 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[14]_i_6_3 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[14]_i_9_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_10 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_2 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_3 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[15]_i_10_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF8 \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[15]_i_9_n_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[15]_i_10_n_0 ),
        .O(new_sboxw[13]),
        .S(tmp_sboxw_0[3]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[15]_i_9 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[15]_i_6_1 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[15]_i_9_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF8 \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[8]_i_8_n_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[8]_i_9_n_0 ),
        .O(new_sboxw[7]),
        .S(tmp_sboxw_0[3]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_8 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_1 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[8]_i_8_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[8]_i_9 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_2 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[8]_i_6_3 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[8]_i_9_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF8 \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[9]_i_7_n_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[9]_i_8_n_0 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11_0 [1]),
        .S(tmp_sboxw_0[3]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_7 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_0 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_1 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[9]_i_7_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF7 \inv_sbox_inferred__0/block_w3_reg_reg[9]_i_8 
       (.I0(\inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_2 ),
        .I1(\inv_sbox_inferred__0/block_w3_reg_reg[9]_i_5_3 ),
        .O(\inv_sbox_inferred__0/block_w3_reg_reg[9]_i_8_n_0 ),
        .S(tmp_sboxw_0[2]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_10 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_1 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_10_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_2 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9_3 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF8 \inv_sbox_inferred__1/block_w3_reg_reg[16]_i_9 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_10_n_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11_n_0 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[16]_i_11_0 [2]),
        .S(tmp_sboxw_0[5]));
  MUXF8 \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[17]_i_7_n_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[17]_i_8_n_0 ),
        .O(new_sboxw[14]),
        .S(tmp_sboxw_0[5]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_7 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_1 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[17]_i_7_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[17]_i_8 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_2 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[17]_i_5_3 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[17]_i_8_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF8 \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[18]_i_7_n_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[18]_i_8_n_0 ),
        .O(new_sboxw[15]),
        .S(tmp_sboxw_0[5]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_7 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_1 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[18]_i_7_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[18]_i_8 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_2 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[18]_i_5_3 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[18]_i_8_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF8 \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[19]_i_7_n_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[19]_i_8_n_0 ),
        .O(new_sboxw[16]),
        .S(tmp_sboxw_0[5]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_7 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_1 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[19]_i_7_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[19]_i_8 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_2 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[19]_i_5_3 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[19]_i_8_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF8 \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[20]_i_7_n_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[20]_i_8_n_0 ),
        .O(new_sboxw[17]),
        .S(tmp_sboxw_0[5]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_7 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_1 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[20]_i_7_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[20]_i_8 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_2 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[20]_i_5_3 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[20]_i_8_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF8 \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[21]_i_8_n_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[21]_i_9_n_0 ),
        .O(new_sboxw[18]),
        .S(tmp_sboxw_0[5]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_8 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_1 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[21]_i_8_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[21]_i_9 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_2 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[21]_i_6_3 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[21]_i_9_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF8 \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[22]_i_8_n_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[22]_i_9_n_0 ),
        .O(new_sboxw[19]),
        .S(tmp_sboxw_0[5]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_8 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_1 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[22]_i_8_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[22]_i_9 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_2 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[22]_i_6_3 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[22]_i_9_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_10 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_2 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_3 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[23]_i_10_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF8 \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[23]_i_9_n_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[23]_i_10_n_0 ),
        .O(new_sboxw[20]),
        .S(tmp_sboxw_0[5]));
  MUXF7 \inv_sbox_inferred__1/block_w3_reg_reg[23]_i_9 
       (.I0(\inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_0 ),
        .I1(\inv_sbox_inferred__1/block_w3_reg_reg[23]_i_6_1 ),
        .O(\inv_sbox_inferred__1/block_w3_reg_reg[23]_i_9_n_0 ),
        .S(tmp_sboxw_0[4]));
  MUXF8 \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[24]_i_8_n_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[24]_i_9_n_0 ),
        .O(new_sboxw[21]),
        .S(tmp_sboxw_0[7]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_8 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_1 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[24]_i_8_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[24]_i_9 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_2 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[24]_i_6_3 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[24]_i_9_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF8 \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[25]_i_7_n_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[25]_i_8_n_0 ),
        .O(new_sboxw[22]),
        .S(tmp_sboxw_0[7]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_7 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_1 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[25]_i_7_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[25]_i_8 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_2 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[25]_i_5_3 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[25]_i_8_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF8 \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[26]_i_7_n_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[26]_i_8_n_0 ),
        .O(new_sboxw[23]),
        .S(tmp_sboxw_0[7]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_7 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_1 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[26]_i_7_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[26]_i_8 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_2 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[26]_i_5_3 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[26]_i_8_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF8 \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[27]_i_6_n_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[27]_i_7_n_0 ),
        .O(new_sboxw[24]),
        .S(tmp_sboxw_0[7]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_6 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_1 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[27]_i_6_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[27]_i_7 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_2 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[27]_i_4_3 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[27]_i_7_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF8 \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[28]_i_7_n_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[28]_i_8_n_0 ),
        .O(new_sboxw[25]),
        .S(tmp_sboxw_0[7]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_7 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_1 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[28]_i_7_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[28]_i_8 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_2 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[28]_i_5_3 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[28]_i_8_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF8 \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[29]_i_8_n_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[29]_i_9_n_0 ),
        .O(new_sboxw[26]),
        .S(tmp_sboxw_0[7]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_8 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_1 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[29]_i_8_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[29]_i_9 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_2 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[29]_i_6_3 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[29]_i_9_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF8 \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[30]_i_8_n_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[30]_i_9_n_0 ),
        .O(new_sboxw[27]),
        .S(tmp_sboxw_0[7]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_8 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_1 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[30]_i_8_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[30]_i_9 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_2 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[30]_i_6_3 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[30]_i_9_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_11 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_1 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[31]_i_11_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF7 \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_12 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_2 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8_3 ),
        .O(\inv_sbox_inferred__2/block_w3_reg_reg[31]_i_12_n_0 ),
        .S(tmp_sboxw_0[6]));
  MUXF8 \inv_sbox_inferred__2/block_w3_reg_reg[31]_i_8 
       (.I0(\inv_sbox_inferred__2/block_w3_reg_reg[31]_i_11_n_0 ),
        .I1(\inv_sbox_inferred__2/block_w3_reg_reg[31]_i_12_n_0 ),
        .O(new_sboxw[28]),
        .S(tmp_sboxw_0[7]));
endmodule

(* ORIG_REF_NAME = "aes_key_mem" *) 
module switch_elements_aes_key_mem
   (\block_w0_reg_reg[31] ,
    \block_w0_reg_reg[30] ,
    \block_w0_reg_reg[29] ,
    \block_w0_reg_reg[28] ,
    \block_w0_reg_reg[25] ,
    \block_w0_reg_reg[24] ,
    \block_w0_reg_reg[23] ,
    \block_w0_reg_reg[16] ,
    \block_w0_reg_reg[22] ,
    \block_w0_reg_reg[21] ,
    \block_w0_reg_reg[20] ,
    \block_w0_reg_reg[19] ,
    \block_w0_reg_reg[17] ,
    \block_w0_reg_reg[15] ,
    \block_w0_reg_reg[14] ,
    \block_w0_reg_reg[13] ,
    \block_w0_reg_reg[12] ,
    \block_w0_reg_reg[10] ,
    \block_w0_reg_reg[9] ,
    \block_w0_reg_reg[8] ,
    \block_w0_reg_reg[7] ,
    \block_w0_reg_reg[6] ,
    \block_w0_reg_reg[0] ,
    \block_w0_reg_reg[5] ,
    \block_w0_reg_reg[4] ,
    \block_w0_reg_reg[3] ,
    \block_w0_reg_reg[2] ,
    \block_w0_reg_reg[1] ,
    \block_w1_reg_reg[31] ,
    \block_w1_reg_reg[30] ,
    \block_w1_reg_reg[29] ,
    \block_w1_reg_reg[28] ,
    \block_w1_reg_reg[25] ,
    \block_w1_reg_reg[24] ,
    \block_w1_reg_reg[23] ,
    \block_w1_reg_reg[16] ,
    \block_w1_reg_reg[22] ,
    \block_w1_reg_reg[21] ,
    \block_w1_reg_reg[20] ,
    \block_w1_reg_reg[19] ,
    \block_w1_reg_reg[17] ,
    \block_w1_reg_reg[15] ,
    \block_w1_reg_reg[9] ,
    \block_w1_reg_reg[14] ,
    \block_w1_reg_reg[13] ,
    \block_w1_reg_reg[12] ,
    \block_w1_reg_reg[10] ,
    \block_w1_reg_reg[8] ,
    \block_w1_reg_reg[7] ,
    \block_w1_reg_reg[6] ,
    \block_w1_reg_reg[0] ,
    \block_w1_reg_reg[5] ,
    \block_w1_reg_reg[4] ,
    \block_w1_reg_reg[3] ,
    \block_w1_reg_reg[2] ,
    \block_w1_reg_reg[1] ,
    \block_w2_reg_reg[31] ,
    \block_w2_reg_reg[30] ,
    \block_w2_reg_reg[29] ,
    \block_w2_reg_reg[28] ,
    \block_w2_reg_reg[25] ,
    \block_w2_reg_reg[24] ,
    \block_w2_reg_reg[23] ,
    \block_w2_reg_reg[16] ,
    \block_w2_reg_reg[22] ,
    \block_w2_reg_reg[21] ,
    \block_w2_reg_reg[20] ,
    \block_w2_reg_reg[19] ,
    \block_w2_reg_reg[17] ,
    \block_w2_reg_reg[15] ,
    \block_w2_reg_reg[9] ,
    \block_w2_reg_reg[14] ,
    \block_w2_reg_reg[13] ,
    \block_w2_reg_reg[12] ,
    \block_w2_reg_reg[10] ,
    \block_w2_reg_reg[8] ,
    \block_w2_reg_reg[7] ,
    \block_w2_reg_reg[6] ,
    \block_w2_reg_reg[0] ,
    \block_w2_reg_reg[5] ,
    \block_w2_reg_reg[4] ,
    \block_w2_reg_reg[3] ,
    \block_w2_reg_reg[2] ,
    \block_w2_reg_reg[1] ,
    \block_w3_reg_reg[31] ,
    \block_w3_reg_reg[30] ,
    \block_w3_reg_reg[29] ,
    \block_w3_reg_reg[28] ,
    \block_w3_reg_reg[25] ,
    \block_w3_reg_reg[24] ,
    \block_w3_reg_reg[23] ,
    \block_w3_reg_reg[16] ,
    \block_w3_reg_reg[22] ,
    \block_w3_reg_reg[21] ,
    \block_w3_reg_reg[20] ,
    \block_w3_reg_reg[19] ,
    \block_w3_reg_reg[17] ,
    \block_w3_reg_reg[15] ,
    \block_w3_reg_reg[14] ,
    \block_w3_reg_reg[13] ,
    \block_w3_reg_reg[12] ,
    \block_w3_reg_reg[10] ,
    \block_w3_reg_reg[9] ,
    \block_w3_reg_reg[8] ,
    \block_w3_reg_reg[7] ,
    \block_w3_reg_reg[6] ,
    \block_w3_reg_reg[0] ,
    \block_w3_reg_reg[5] ,
    \block_w3_reg_reg[4] ,
    \block_w3_reg_reg[3] ,
    \block_w3_reg_reg[2] ,
    \block_w3_reg_reg[1] ,
    \block_reg_reg[3][0] ,
    round_key,
    \block_reg_reg[0][16] ,
    \block_reg_reg[0][0] ,
    \block_reg_reg[1][16] ,
    \block_reg_reg[1][0] ,
    \block_reg_reg[2][16] ,
    \block_reg_reg[2][0] ,
    \block_reg_reg[3][16] ,
    Q,
    \rcon_reg_reg[7]_0 ,
    \block_w1_reg_reg[31]_0 ,
    \block_w2_reg_reg[31]_0 ,
    \block_w3_reg_reg[31]_0 ,
    \block_w0_reg_reg[31]_0 ,
    \block_w3_reg_reg[8]_0 ,
    \block_w0_reg_reg[8]_0 ,
    \block_w3_reg_reg[0]_0 ,
    \block_w0_reg_reg[0]_0 ,
    \block_w1_reg_reg[0]_0 ,
    \block_w2_reg_reg[0]_0 ,
    inv_mixcolumns_return0__55,
    inv_mixcolumns_return0124_out__47,
    inv_mixcolumns_return0110_out__47,
    inv_mixcolumns_return0117_out__50,
    p_0_out,
    inv_mixcolumns_return0198_out__63,
    inv_mixcolumns_return0213_out__55,
    inv_mixcolumns_return0206_out__55,
    inv_mixcolumns_return0220_out__63,
    inv_mixcolumns_return0174_out__63,
    inv_mixcolumns_return0166_out__55,
    inv_mixcolumns_return0181_out__58,
    inv_mixcolumns_return0188_out__55,
    addroundkey_return,
    inv_mixcolumns_return0134_out__63,
    inv_mixcolumns_return0149_out__55,
    inv_mixcolumns_return0142_out__55,
    inv_mixcolumns_return0156_out__63,
    ready_new,
    key_ready,
    init_state,
    \block_w0_reg_reg[31]_1 ,
    p_1_in,
    core_block,
    \block_w0_reg_reg[0]_1 ,
    core_key,
    \key_mem_reg[14][36]_0 ,
    \key_mem_reg[14][127]_0 ,
    new_sboxw,
    p_19_in,
    \block_w0_reg_reg[16]_0 ,
    muxed_round_nr,
    \block_w0_reg_reg[31]_2 ,
    dec_new_block,
    \block_w3_reg_reg[26] ,
    ready_reg_reg_0,
    enc_ready,
    dec_ready,
    clk_i,
    rst_i,
    \block_w3_reg[30]_i_4_0 ,
    \block_w3_reg[30]_i_4_1 ,
    \block_w3_reg[1]_i_4__0_0 ,
    \block_w0_reg[31]_i_6__0_0 ,
    \block_w0_reg[31]_i_6__0_1 ,
    \block_w2_reg[29]_i_4_0 ,
    \block_w2_reg[29]_i_4_1 ,
    \block_w1_reg[29]_i_4_0 ,
    \block_w1_reg[29]_i_4_1 );
  output \block_w0_reg_reg[31] ;
  output \block_w0_reg_reg[30] ;
  output \block_w0_reg_reg[29] ;
  output \block_w0_reg_reg[28] ;
  output \block_w0_reg_reg[25] ;
  output \block_w0_reg_reg[24] ;
  output \block_w0_reg_reg[23] ;
  output [0:0]\block_w0_reg_reg[16] ;
  output \block_w0_reg_reg[22] ;
  output \block_w0_reg_reg[21] ;
  output \block_w0_reg_reg[20] ;
  output \block_w0_reg_reg[19] ;
  output \block_w0_reg_reg[17] ;
  output \block_w0_reg_reg[15] ;
  output \block_w0_reg_reg[14] ;
  output \block_w0_reg_reg[13] ;
  output \block_w0_reg_reg[12] ;
  output \block_w0_reg_reg[10] ;
  output \block_w0_reg_reg[9] ;
  output \block_w0_reg_reg[8] ;
  output \block_w0_reg_reg[7] ;
  output \block_w0_reg_reg[6] ;
  output [0:0]\block_w0_reg_reg[0] ;
  output \block_w0_reg_reg[5] ;
  output \block_w0_reg_reg[4] ;
  output \block_w0_reg_reg[3] ;
  output \block_w0_reg_reg[2] ;
  output \block_w0_reg_reg[1] ;
  output \block_w1_reg_reg[31] ;
  output \block_w1_reg_reg[30] ;
  output \block_w1_reg_reg[29] ;
  output \block_w1_reg_reg[28] ;
  output \block_w1_reg_reg[25] ;
  output \block_w1_reg_reg[24] ;
  output \block_w1_reg_reg[23] ;
  output [0:0]\block_w1_reg_reg[16] ;
  output \block_w1_reg_reg[22] ;
  output \block_w1_reg_reg[21] ;
  output \block_w1_reg_reg[20] ;
  output \block_w1_reg_reg[19] ;
  output \block_w1_reg_reg[17] ;
  output \block_w1_reg_reg[15] ;
  output [0:0]\block_w1_reg_reg[9] ;
  output \block_w1_reg_reg[14] ;
  output \block_w1_reg_reg[13] ;
  output \block_w1_reg_reg[12] ;
  output \block_w1_reg_reg[10] ;
  output \block_w1_reg_reg[8] ;
  output \block_w1_reg_reg[7] ;
  output \block_w1_reg_reg[6] ;
  output [0:0]\block_w1_reg_reg[0] ;
  output \block_w1_reg_reg[5] ;
  output \block_w1_reg_reg[4] ;
  output \block_w1_reg_reg[3] ;
  output \block_w1_reg_reg[2] ;
  output \block_w1_reg_reg[1] ;
  output \block_w2_reg_reg[31] ;
  output \block_w2_reg_reg[30] ;
  output \block_w2_reg_reg[29] ;
  output \block_w2_reg_reg[28] ;
  output \block_w2_reg_reg[25] ;
  output \block_w2_reg_reg[24] ;
  output \block_w2_reg_reg[23] ;
  output [0:0]\block_w2_reg_reg[16] ;
  output \block_w2_reg_reg[22] ;
  output \block_w2_reg_reg[21] ;
  output \block_w2_reg_reg[20] ;
  output \block_w2_reg_reg[19] ;
  output \block_w2_reg_reg[17] ;
  output \block_w2_reg_reg[15] ;
  output [0:0]\block_w2_reg_reg[9] ;
  output \block_w2_reg_reg[14] ;
  output \block_w2_reg_reg[13] ;
  output \block_w2_reg_reg[12] ;
  output \block_w2_reg_reg[10] ;
  output \block_w2_reg_reg[8] ;
  output \block_w2_reg_reg[7] ;
  output \block_w2_reg_reg[6] ;
  output [0:0]\block_w2_reg_reg[0] ;
  output \block_w2_reg_reg[5] ;
  output \block_w2_reg_reg[4] ;
  output \block_w2_reg_reg[3] ;
  output \block_w2_reg_reg[2] ;
  output \block_w2_reg_reg[1] ;
  output \block_w3_reg_reg[31] ;
  output \block_w3_reg_reg[30] ;
  output \block_w3_reg_reg[29] ;
  output \block_w3_reg_reg[28] ;
  output \block_w3_reg_reg[25] ;
  output \block_w3_reg_reg[24] ;
  output \block_w3_reg_reg[23] ;
  output [0:0]\block_w3_reg_reg[16] ;
  output \block_w3_reg_reg[22] ;
  output \block_w3_reg_reg[21] ;
  output \block_w3_reg_reg[20] ;
  output \block_w3_reg_reg[19] ;
  output \block_w3_reg_reg[17] ;
  output \block_w3_reg_reg[15] ;
  output \block_w3_reg_reg[14] ;
  output \block_w3_reg_reg[13] ;
  output \block_w3_reg_reg[12] ;
  output \block_w3_reg_reg[10] ;
  output \block_w3_reg_reg[9] ;
  output \block_w3_reg_reg[8] ;
  output \block_w3_reg_reg[7] ;
  output \block_w3_reg_reg[6] ;
  output [0:0]\block_w3_reg_reg[0] ;
  output \block_w3_reg_reg[5] ;
  output \block_w3_reg_reg[4] ;
  output \block_w3_reg_reg[3] ;
  output \block_w3_reg_reg[2] ;
  output \block_w3_reg_reg[1] ;
  output \block_reg_reg[3][0] ;
  output [127:0]round_key;
  output \block_reg_reg[0][16] ;
  output \block_reg_reg[0][0] ;
  output \block_reg_reg[1][16] ;
  output \block_reg_reg[1][0] ;
  output \block_reg_reg[2][16] ;
  output \block_reg_reg[2][0] ;
  output \block_reg_reg[3][16] ;
  output [31:0]Q;
  output [7:0]\rcon_reg_reg[7]_0 ;
  output \block_w1_reg_reg[31]_0 ;
  output \block_w2_reg_reg[31]_0 ;
  output \block_w3_reg_reg[31]_0 ;
  output \block_w0_reg_reg[31]_0 ;
  output \block_w3_reg_reg[8]_0 ;
  output \block_w0_reg_reg[8]_0 ;
  output \block_w3_reg_reg[0]_0 ;
  output \block_w0_reg_reg[0]_0 ;
  output \block_w1_reg_reg[0]_0 ;
  output \block_w2_reg_reg[0]_0 ;
  output [6:0]inv_mixcolumns_return0__55;
  output [7:0]inv_mixcolumns_return0124_out__47;
  output [6:0]inv_mixcolumns_return0110_out__47;
  output [6:0]inv_mixcolumns_return0117_out__50;
  output [75:0]p_0_out;
  output [6:0]inv_mixcolumns_return0198_out__63;
  output [6:0]inv_mixcolumns_return0213_out__55;
  output [6:0]inv_mixcolumns_return0206_out__55;
  output [7:0]inv_mixcolumns_return0220_out__63;
  output [7:0]inv_mixcolumns_return0174_out__63;
  output [6:0]inv_mixcolumns_return0166_out__55;
  output [6:0]inv_mixcolumns_return0181_out__58;
  output [7:0]inv_mixcolumns_return0188_out__55;
  output [43:0]addroundkey_return;
  output [6:0]inv_mixcolumns_return0134_out__63;
  output [6:0]inv_mixcolumns_return0149_out__55;
  output [7:0]inv_mixcolumns_return0142_out__55;
  output [7:0]inv_mixcolumns_return0156_out__63;
  output ready_new;
  output key_ready;
  output init_state;
  input \block_w0_reg_reg[31]_1 ;
  input [2:0]p_1_in;
  input [127:0]core_block;
  input [0:0]\block_w0_reg_reg[0]_1 ;
  input [255:0]core_key;
  input \key_mem_reg[14][36]_0 ;
  input \key_mem_reg[14][127]_0 ;
  input [31:0]new_sboxw;
  input [7:0]p_19_in;
  input [2:0]\block_w0_reg_reg[16]_0 ;
  input [3:0]muxed_round_nr;
  input \block_w0_reg_reg[31]_2 ;
  input [127:0]dec_new_block;
  input \block_w3_reg_reg[26] ;
  input [1:0]ready_reg_reg_0;
  input enc_ready;
  input dec_ready;
  input clk_i;
  input rst_i;
  input \block_w3_reg[30]_i_4_0 ;
  input \block_w3_reg[30]_i_4_1 ;
  input \block_w3_reg[1]_i_4__0_0 ;
  input \block_w0_reg[31]_i_6__0_0 ;
  input \block_w0_reg[31]_i_6__0_1 ;
  input \block_w2_reg[29]_i_4_0 ;
  input \block_w2_reg[29]_i_4_1 ;
  input \block_w1_reg[29]_i_4_0 ;
  input \block_w1_reg[29]_i_4_1 ;

  wire \FSM_sequential_key_mem_ctrl_reg[1]_i_1_n_0 ;
  wire [31:0]Q;
  wire [43:0]addroundkey_return;
  wire \block_reg_reg[0][0] ;
  wire \block_reg_reg[0][16] ;
  wire \block_reg_reg[1][0] ;
  wire \block_reg_reg[1][16] ;
  wire \block_reg_reg[2][0] ;
  wire \block_reg_reg[2][16] ;
  wire \block_reg_reg[3][0] ;
  wire \block_reg_reg[3][16] ;
  wire \block_w0_reg[0]_i_5__0_n_0 ;
  wire \block_w0_reg[0]_i_5_n_0 ;
  wire \block_w0_reg[0]_i_6_n_0 ;
  wire \block_w0_reg[0]_i_7_n_0 ;
  wire \block_w0_reg[0]_i_8_n_0 ;
  wire \block_w0_reg[10]_i_5__0_n_0 ;
  wire \block_w0_reg[10]_i_6__0_n_0 ;
  wire \block_w0_reg[10]_i_7_n_0 ;
  wire \block_w0_reg[10]_i_8_n_0 ;
  wire \block_w0_reg[11]_i_5__0_n_0 ;
  wire \block_w0_reg[11]_i_6_n_0 ;
  wire \block_w0_reg[11]_i_7_n_0 ;
  wire \block_w0_reg[11]_i_8_n_0 ;
  wire \block_w0_reg[11]_i_9_n_0 ;
  wire \block_w0_reg[12]_i_6__0_n_0 ;
  wire \block_w0_reg[12]_i_6_n_0 ;
  wire \block_w0_reg[12]_i_7_n_0 ;
  wire \block_w0_reg[12]_i_8_n_0 ;
  wire \block_w0_reg[12]_i_9_n_0 ;
  wire \block_w0_reg[13]_i_5__0_n_0 ;
  wire \block_w0_reg[13]_i_6__0_n_0 ;
  wire \block_w0_reg[13]_i_7__0_n_0 ;
  wire \block_w0_reg[13]_i_7_n_0 ;
  wire \block_w0_reg[13]_i_8_n_0 ;
  wire \block_w0_reg[14]_i_5__0_n_0 ;
  wire \block_w0_reg[14]_i_6__0_n_0 ;
  wire \block_w0_reg[14]_i_7__0_n_0 ;
  wire \block_w0_reg[14]_i_7_n_0 ;
  wire \block_w0_reg[14]_i_8_n_0 ;
  wire \block_w0_reg[15]_i_5__0_n_0 ;
  wire \block_w0_reg[15]_i_6__0_n_0 ;
  wire \block_w0_reg[15]_i_7_n_0 ;
  wire \block_w0_reg[15]_i_8_n_0 ;
  wire \block_w0_reg[16]_i_5__0_n_0 ;
  wire \block_w0_reg[16]_i_5_n_0 ;
  wire \block_w0_reg[16]_i_6__0_n_0 ;
  wire \block_w0_reg[16]_i_6_n_0 ;
  wire \block_w0_reg[16]_i_7_n_0 ;
  wire \block_w0_reg[16]_i_8_n_0 ;
  wire \block_w0_reg[17]_i_6_n_0 ;
  wire \block_w0_reg[17]_i_7_n_0 ;
  wire \block_w0_reg[17]_i_8_n_0 ;
  wire \block_w0_reg[17]_i_9_n_0 ;
  wire \block_w0_reg[18]_i_5__0_n_0 ;
  wire \block_w0_reg[18]_i_6__0_n_0 ;
  wire \block_w0_reg[18]_i_6_n_0 ;
  wire \block_w0_reg[18]_i_7_n_0 ;
  wire \block_w0_reg[18]_i_8_n_0 ;
  wire \block_w0_reg[19]_i_6__0_n_0 ;
  wire \block_w0_reg[19]_i_6_n_0 ;
  wire \block_w0_reg[19]_i_7__0_n_0 ;
  wire \block_w0_reg[19]_i_8__0_n_0 ;
  wire \block_w0_reg[19]_i_9_n_0 ;
  wire \block_w0_reg[1]_i_6_n_0 ;
  wire \block_w0_reg[1]_i_7_n_0 ;
  wire \block_w0_reg[1]_i_8_n_0 ;
  wire \block_w0_reg[1]_i_9_n_0 ;
  wire \block_w0_reg[20]_i_10_n_0 ;
  wire \block_w0_reg[20]_i_7_n_0 ;
  wire \block_w0_reg[20]_i_8_n_0 ;
  wire \block_w0_reg[20]_i_9_n_0 ;
  wire \block_w0_reg[21]_i_5__0_n_0 ;
  wire \block_w0_reg[21]_i_6__0_n_0 ;
  wire \block_w0_reg[21]_i_7__0_n_0 ;
  wire \block_w0_reg[21]_i_7_n_0 ;
  wire \block_w0_reg[21]_i_8_n_0 ;
  wire \block_w0_reg[22]_i_5__0_n_0 ;
  wire \block_w0_reg[22]_i_6__0_n_0 ;
  wire \block_w0_reg[22]_i_7__0_n_0 ;
  wire \block_w0_reg[22]_i_7_n_0 ;
  wire \block_w0_reg[22]_i_8_n_0 ;
  wire \block_w0_reg[23]_i_5__0_n_0 ;
  wire \block_w0_reg[23]_i_6__0_n_0 ;
  wire \block_w0_reg[23]_i_7_n_0 ;
  wire \block_w0_reg[23]_i_8_n_0 ;
  wire \block_w0_reg[24]_i_5__0_n_0 ;
  wire \block_w0_reg[24]_i_6__0_n_0 ;
  wire \block_w0_reg[24]_i_7_n_0 ;
  wire \block_w0_reg[24]_i_8_n_0 ;
  wire \block_w0_reg[25]_i_10_n_0 ;
  wire \block_w0_reg[25]_i_6_n_0 ;
  wire \block_w0_reg[25]_i_7_n_0 ;
  wire \block_w0_reg[25]_i_8_n_0 ;
  wire \block_w0_reg[25]_i_9_n_0 ;
  wire \block_w0_reg[26]_i_5__0_n_0 ;
  wire \block_w0_reg[26]_i_6__0_n_0 ;
  wire \block_w0_reg[26]_i_6_n_0 ;
  wire \block_w0_reg[26]_i_7_n_0 ;
  wire \block_w0_reg[26]_i_8_n_0 ;
  wire \block_w0_reg[27]_i_10_n_0 ;
  wire \block_w0_reg[27]_i_6_n_0 ;
  wire \block_w0_reg[27]_i_7_n_0 ;
  wire \block_w0_reg[27]_i_8_n_0 ;
  wire \block_w0_reg[28]_i_10_n_0 ;
  wire \block_w0_reg[28]_i_6__0_n_0 ;
  wire \block_w0_reg[28]_i_6_n_0 ;
  wire \block_w0_reg[28]_i_7_n_0 ;
  wire \block_w0_reg[28]_i_8_n_0 ;
  wire \block_w0_reg[29]_i_5__0_n_0 ;
  wire \block_w0_reg[29]_i_6__0_n_0 ;
  wire \block_w0_reg[29]_i_7__0_n_0 ;
  wire \block_w0_reg[29]_i_7_n_0 ;
  wire \block_w0_reg[29]_i_8_n_0 ;
  wire \block_w0_reg[2]_i_5__0_n_0 ;
  wire \block_w0_reg[2]_i_6__0_n_0 ;
  wire \block_w0_reg[2]_i_7_n_0 ;
  wire \block_w0_reg[2]_i_8_n_0 ;
  wire \block_w0_reg[30]_i_5__0_n_0 ;
  wire \block_w0_reg[30]_i_6__0_n_0 ;
  wire \block_w0_reg[30]_i_7__0_n_0 ;
  wire \block_w0_reg[30]_i_7_n_0 ;
  wire \block_w0_reg[30]_i_8_n_0 ;
  wire \block_w0_reg[31]_i_6__0_0 ;
  wire \block_w0_reg[31]_i_6__0_1 ;
  wire \block_w0_reg[31]_i_6__0_n_0 ;
  wire \block_w0_reg[31]_i_7_n_0 ;
  wire \block_w0_reg[31]_i_8_n_0 ;
  wire \block_w0_reg[31]_i_9_n_0 ;
  wire \block_w0_reg[3]_i_6__0_n_0 ;
  wire \block_w0_reg[3]_i_6_n_0 ;
  wire \block_w0_reg[3]_i_7__0_n_0 ;
  wire \block_w0_reg[3]_i_7_n_0 ;
  wire \block_w0_reg[3]_i_8_n_0 ;
  wire \block_w0_reg[3]_i_9_n_0 ;
  wire \block_w0_reg[4]_i_10_n_0 ;
  wire \block_w0_reg[4]_i_7_n_0 ;
  wire \block_w0_reg[4]_i_8_n_0 ;
  wire \block_w0_reg[4]_i_9_n_0 ;
  wire \block_w0_reg[5]_i_5__0_n_0 ;
  wire \block_w0_reg[5]_i_6__0_n_0 ;
  wire \block_w0_reg[5]_i_7__0_n_0 ;
  wire \block_w0_reg[5]_i_7_n_0 ;
  wire \block_w0_reg[5]_i_8_n_0 ;
  wire \block_w0_reg[6]_i_5__0_n_0 ;
  wire \block_w0_reg[6]_i_6__0_n_0 ;
  wire \block_w0_reg[6]_i_7__0_n_0 ;
  wire \block_w0_reg[6]_i_7_n_0 ;
  wire \block_w0_reg[6]_i_8_n_0 ;
  wire \block_w0_reg[7]_i_4_n_0 ;
  wire \block_w0_reg[7]_i_5__0_n_0 ;
  wire \block_w0_reg[7]_i_6__0_n_0 ;
  wire \block_w0_reg[7]_i_7_n_0 ;
  wire \block_w0_reg[7]_i_8_n_0 ;
  wire \block_w0_reg[8]_i_5__0_n_0 ;
  wire \block_w0_reg[8]_i_6_n_0 ;
  wire \block_w0_reg[8]_i_7_n_0 ;
  wire \block_w0_reg[8]_i_8_n_0 ;
  wire \block_w0_reg[9]_i_10_n_0 ;
  wire \block_w0_reg[9]_i_6__0_n_0 ;
  wire \block_w0_reg[9]_i_7__0_n_0 ;
  wire \block_w0_reg[9]_i_7_n_0 ;
  wire \block_w0_reg[9]_i_8_n_0 ;
  wire \block_w0_reg[9]_i_9_n_0 ;
  wire [0:0]\block_w0_reg_reg[0] ;
  wire \block_w0_reg_reg[0]_0 ;
  wire [0:0]\block_w0_reg_reg[0]_1 ;
  wire \block_w0_reg_reg[10] ;
  wire \block_w0_reg_reg[12] ;
  wire \block_w0_reg_reg[13] ;
  wire \block_w0_reg_reg[14] ;
  wire \block_w0_reg_reg[15] ;
  wire [0:0]\block_w0_reg_reg[16] ;
  wire [2:0]\block_w0_reg_reg[16]_0 ;
  wire \block_w0_reg_reg[17] ;
  wire \block_w0_reg_reg[19] ;
  wire \block_w0_reg_reg[1] ;
  wire \block_w0_reg_reg[20] ;
  wire \block_w0_reg_reg[21] ;
  wire \block_w0_reg_reg[22] ;
  wire \block_w0_reg_reg[23] ;
  wire \block_w0_reg_reg[24] ;
  wire \block_w0_reg_reg[25] ;
  wire \block_w0_reg_reg[28] ;
  wire \block_w0_reg_reg[29] ;
  wire \block_w0_reg_reg[2] ;
  wire \block_w0_reg_reg[30] ;
  wire \block_w0_reg_reg[31] ;
  wire \block_w0_reg_reg[31]_0 ;
  wire \block_w0_reg_reg[31]_1 ;
  wire \block_w0_reg_reg[31]_2 ;
  wire \block_w0_reg_reg[3] ;
  wire \block_w0_reg_reg[4] ;
  wire \block_w0_reg_reg[5] ;
  wire \block_w0_reg_reg[6] ;
  wire \block_w0_reg_reg[7] ;
  wire \block_w0_reg_reg[8] ;
  wire \block_w0_reg_reg[8]_0 ;
  wire \block_w0_reg_reg[9] ;
  wire \block_w1_reg[0]_i_5__0_n_0 ;
  wire \block_w1_reg[0]_i_5_n_0 ;
  wire \block_w1_reg[0]_i_6_n_0 ;
  wire \block_w1_reg[0]_i_7_n_0 ;
  wire \block_w1_reg[0]_i_8_n_0 ;
  wire \block_w1_reg[10]_i_5__0_n_0 ;
  wire \block_w1_reg[10]_i_6__0_n_0 ;
  wire \block_w1_reg[10]_i_7_n_0 ;
  wire \block_w1_reg[10]_i_8_n_0 ;
  wire \block_w1_reg[11]_i_5__0_n_0 ;
  wire \block_w1_reg[11]_i_6_n_0 ;
  wire \block_w1_reg[11]_i_7_n_0 ;
  wire \block_w1_reg[11]_i_8_n_0 ;
  wire \block_w1_reg[11]_i_9_n_0 ;
  wire \block_w1_reg[12]_i_6__0_n_0 ;
  wire \block_w1_reg[12]_i_6_n_0 ;
  wire \block_w1_reg[12]_i_7__0_n_0 ;
  wire \block_w1_reg[12]_i_7_n_0 ;
  wire \block_w1_reg[12]_i_8_n_0 ;
  wire \block_w1_reg[12]_i_9_n_0 ;
  wire \block_w1_reg[13]_i_5__0_n_0 ;
  wire \block_w1_reg[13]_i_6__0_n_0 ;
  wire \block_w1_reg[13]_i_7__0_n_0 ;
  wire \block_w1_reg[13]_i_7_n_0 ;
  wire \block_w1_reg[13]_i_8_n_0 ;
  wire \block_w1_reg[14]_i_5__0_n_0 ;
  wire \block_w1_reg[14]_i_6__0_n_0 ;
  wire \block_w1_reg[14]_i_7__0_n_0 ;
  wire \block_w1_reg[14]_i_7_n_0 ;
  wire \block_w1_reg[14]_i_8_n_0 ;
  wire \block_w1_reg[15]_i_5__0_n_0 ;
  wire \block_w1_reg[15]_i_6__0_n_0 ;
  wire \block_w1_reg[15]_i_7_n_0 ;
  wire \block_w1_reg[15]_i_8_n_0 ;
  wire \block_w1_reg[16]_i_5__0_n_0 ;
  wire \block_w1_reg[16]_i_5_n_0 ;
  wire \block_w1_reg[16]_i_6__0_n_0 ;
  wire \block_w1_reg[16]_i_6_n_0 ;
  wire \block_w1_reg[16]_i_7_n_0 ;
  wire \block_w1_reg[16]_i_8_n_0 ;
  wire \block_w1_reg[17]_i_6_n_0 ;
  wire \block_w1_reg[17]_i_7_n_0 ;
  wire \block_w1_reg[17]_i_8_n_0 ;
  wire \block_w1_reg[17]_i_9_n_0 ;
  wire \block_w1_reg[18]_i_5__0_n_0 ;
  wire \block_w1_reg[18]_i_6__0_n_0 ;
  wire \block_w1_reg[18]_i_6_n_0 ;
  wire \block_w1_reg[18]_i_7_n_0 ;
  wire \block_w1_reg[18]_i_8_n_0 ;
  wire \block_w1_reg[19]_i_6__0_n_0 ;
  wire \block_w1_reg[19]_i_6_n_0 ;
  wire \block_w1_reg[19]_i_7__0_n_0 ;
  wire \block_w1_reg[19]_i_8__0_n_0 ;
  wire \block_w1_reg[19]_i_9_n_0 ;
  wire \block_w1_reg[1]_i_6_n_0 ;
  wire \block_w1_reg[1]_i_7_n_0 ;
  wire \block_w1_reg[1]_i_8_n_0 ;
  wire \block_w1_reg[1]_i_9_n_0 ;
  wire \block_w1_reg[20]_i_10_n_0 ;
  wire \block_w1_reg[20]_i_7_n_0 ;
  wire \block_w1_reg[20]_i_8_n_0 ;
  wire \block_w1_reg[20]_i_9_n_0 ;
  wire \block_w1_reg[21]_i_5__0_n_0 ;
  wire \block_w1_reg[21]_i_6__0_n_0 ;
  wire \block_w1_reg[21]_i_7__0_n_0 ;
  wire \block_w1_reg[21]_i_7_n_0 ;
  wire \block_w1_reg[21]_i_8_n_0 ;
  wire \block_w1_reg[22]_i_5__0_n_0 ;
  wire \block_w1_reg[22]_i_6__0_n_0 ;
  wire \block_w1_reg[22]_i_7__0_n_0 ;
  wire \block_w1_reg[22]_i_7_n_0 ;
  wire \block_w1_reg[22]_i_8_n_0 ;
  wire \block_w1_reg[23]_i_5__0_n_0 ;
  wire \block_w1_reg[23]_i_6__0_n_0 ;
  wire \block_w1_reg[23]_i_7__0_n_0 ;
  wire \block_w1_reg[23]_i_7_n_0 ;
  wire \block_w1_reg[23]_i_8_n_0 ;
  wire \block_w1_reg[24]_i_5__0_n_0 ;
  wire \block_w1_reg[24]_i_6__0_n_0 ;
  wire \block_w1_reg[24]_i_7__0_n_0 ;
  wire \block_w1_reg[24]_i_7_n_0 ;
  wire \block_w1_reg[24]_i_8_n_0 ;
  wire \block_w1_reg[25]_i_10_n_0 ;
  wire \block_w1_reg[25]_i_7_n_0 ;
  wire \block_w1_reg[25]_i_8_n_0 ;
  wire \block_w1_reg[25]_i_9_n_0 ;
  wire \block_w1_reg[26]_i_5__0_n_0 ;
  wire \block_w1_reg[26]_i_6__0_n_0 ;
  wire \block_w1_reg[26]_i_6_n_0 ;
  wire \block_w1_reg[26]_i_7_n_0 ;
  wire \block_w1_reg[26]_i_8_n_0 ;
  wire \block_w1_reg[27]_i_10_n_0 ;
  wire \block_w1_reg[27]_i_6__0_n_0 ;
  wire \block_w1_reg[27]_i_6_n_0 ;
  wire \block_w1_reg[27]_i_7_n_0 ;
  wire \block_w1_reg[27]_i_8_n_0 ;
  wire \block_w1_reg[28]_i_10_n_0 ;
  wire \block_w1_reg[28]_i_6__0_n_0 ;
  wire \block_w1_reg[28]_i_6_n_0 ;
  wire \block_w1_reg[28]_i_7__0_n_0 ;
  wire \block_w1_reg[28]_i_7_n_0 ;
  wire \block_w1_reg[28]_i_8_n_0 ;
  wire \block_w1_reg[29]_i_4_0 ;
  wire \block_w1_reg[29]_i_4_1 ;
  wire \block_w1_reg[29]_i_5__0_n_0 ;
  wire \block_w1_reg[29]_i_6__0_n_0 ;
  wire \block_w1_reg[29]_i_7__0_n_0 ;
  wire \block_w1_reg[29]_i_7_n_0 ;
  wire \block_w1_reg[29]_i_8_n_0 ;
  wire \block_w1_reg[2]_i_5__0_n_0 ;
  wire \block_w1_reg[2]_i_6__0_n_0 ;
  wire \block_w1_reg[2]_i_7_n_0 ;
  wire \block_w1_reg[2]_i_8_n_0 ;
  wire \block_w1_reg[30]_i_5__0_n_0 ;
  wire \block_w1_reg[30]_i_6__0_n_0 ;
  wire \block_w1_reg[30]_i_7__0_n_0 ;
  wire \block_w1_reg[30]_i_7_n_0 ;
  wire \block_w1_reg[30]_i_8_n_0 ;
  wire \block_w1_reg[31]_i_6__0_n_0 ;
  wire \block_w1_reg[31]_i_7__0_n_0 ;
  wire \block_w1_reg[31]_i_8_n_0 ;
  wire \block_w1_reg[31]_i_9_n_0 ;
  wire \block_w1_reg[3]_i_6__0_n_0 ;
  wire \block_w1_reg[3]_i_6_n_0 ;
  wire \block_w1_reg[3]_i_7__0_n_0 ;
  wire \block_w1_reg[3]_i_7_n_0 ;
  wire \block_w1_reg[3]_i_8__0_n_0 ;
  wire \block_w1_reg[3]_i_8_n_0 ;
  wire \block_w1_reg[3]_i_9_n_0 ;
  wire \block_w1_reg[4]_i_10_n_0 ;
  wire \block_w1_reg[4]_i_7_n_0 ;
  wire \block_w1_reg[4]_i_8_n_0 ;
  wire \block_w1_reg[4]_i_9_n_0 ;
  wire \block_w1_reg[5]_i_5__0_n_0 ;
  wire \block_w1_reg[5]_i_6__0_n_0 ;
  wire \block_w1_reg[5]_i_7__0_n_0 ;
  wire \block_w1_reg[5]_i_7_n_0 ;
  wire \block_w1_reg[5]_i_8_n_0 ;
  wire \block_w1_reg[6]_i_5__0_n_0 ;
  wire \block_w1_reg[6]_i_6__0_n_0 ;
  wire \block_w1_reg[6]_i_7__0_n_0 ;
  wire \block_w1_reg[6]_i_7_n_0 ;
  wire \block_w1_reg[6]_i_8_n_0 ;
  wire \block_w1_reg[7]_i_4_n_0 ;
  wire \block_w1_reg[7]_i_5__0_n_0 ;
  wire \block_w1_reg[7]_i_6__0_n_0 ;
  wire \block_w1_reg[7]_i_7__0_n_0 ;
  wire \block_w1_reg[7]_i_7_n_0 ;
  wire \block_w1_reg[7]_i_8_n_0 ;
  wire \block_w1_reg[8]_i_5__0_n_0 ;
  wire \block_w1_reg[8]_i_6__0_n_0 ;
  wire \block_w1_reg[8]_i_7__0_n_0 ;
  wire \block_w1_reg[8]_i_7_n_0 ;
  wire \block_w1_reg[8]_i_8_n_0 ;
  wire \block_w1_reg[9]_i_10_n_0 ;
  wire \block_w1_reg[9]_i_5_n_0 ;
  wire \block_w1_reg[9]_i_6__0_n_0 ;
  wire \block_w1_reg[9]_i_7_n_0 ;
  wire \block_w1_reg[9]_i_8_n_0 ;
  wire \block_w1_reg[9]_i_9_n_0 ;
  wire [0:0]\block_w1_reg_reg[0] ;
  wire \block_w1_reg_reg[0]_0 ;
  wire \block_w1_reg_reg[10] ;
  wire \block_w1_reg_reg[12] ;
  wire \block_w1_reg_reg[13] ;
  wire \block_w1_reg_reg[14] ;
  wire \block_w1_reg_reg[15] ;
  wire [0:0]\block_w1_reg_reg[16] ;
  wire \block_w1_reg_reg[17] ;
  wire \block_w1_reg_reg[19] ;
  wire \block_w1_reg_reg[1] ;
  wire \block_w1_reg_reg[20] ;
  wire \block_w1_reg_reg[21] ;
  wire \block_w1_reg_reg[22] ;
  wire \block_w1_reg_reg[23] ;
  wire \block_w1_reg_reg[24] ;
  wire \block_w1_reg_reg[25] ;
  wire \block_w1_reg_reg[28] ;
  wire \block_w1_reg_reg[29] ;
  wire \block_w1_reg_reg[2] ;
  wire \block_w1_reg_reg[30] ;
  wire \block_w1_reg_reg[31] ;
  wire \block_w1_reg_reg[31]_0 ;
  wire \block_w1_reg_reg[3] ;
  wire \block_w1_reg_reg[4] ;
  wire \block_w1_reg_reg[5] ;
  wire \block_w1_reg_reg[6] ;
  wire \block_w1_reg_reg[7] ;
  wire \block_w1_reg_reg[8] ;
  wire [0:0]\block_w1_reg_reg[9] ;
  wire \block_w2_reg[0]_i_11_n_0 ;
  wire \block_w2_reg[0]_i_5_n_0 ;
  wire \block_w2_reg[0]_i_6__0_n_0 ;
  wire \block_w2_reg[0]_i_6_n_0 ;
  wire \block_w2_reg[0]_i_7_n_0 ;
  wire \block_w2_reg[0]_i_8_n_0 ;
  wire \block_w2_reg[10]_i_11_n_0 ;
  wire \block_w2_reg[10]_i_6__0_n_0 ;
  wire \block_w2_reg[10]_i_7_n_0 ;
  wire \block_w2_reg[10]_i_8_n_0 ;
  wire \block_w2_reg[11]_i_12_n_0 ;
  wire \block_w2_reg[11]_i_5_n_0 ;
  wire \block_w2_reg[11]_i_7_n_0 ;
  wire \block_w2_reg[11]_i_8_n_0 ;
  wire \block_w2_reg[11]_i_9_n_0 ;
  wire \block_w2_reg[12]_i_12_n_0 ;
  wire \block_w2_reg[12]_i_6_n_0 ;
  wire \block_w2_reg[12]_i_7__0_n_0 ;
  wire \block_w2_reg[12]_i_7_n_0 ;
  wire \block_w2_reg[12]_i_8_n_0 ;
  wire \block_w2_reg[12]_i_9_n_0 ;
  wire \block_w2_reg[13]_i_11_n_0 ;
  wire \block_w2_reg[13]_i_6__0_n_0 ;
  wire \block_w2_reg[13]_i_7__0_n_0 ;
  wire \block_w2_reg[13]_i_7_n_0 ;
  wire \block_w2_reg[13]_i_8__0_n_0 ;
  wire \block_w2_reg[13]_i_8_n_0 ;
  wire \block_w2_reg[14]_i_11_n_0 ;
  wire \block_w2_reg[14]_i_6__0_n_0 ;
  wire \block_w2_reg[14]_i_7__0_n_0 ;
  wire \block_w2_reg[14]_i_7_n_0 ;
  wire \block_w2_reg[14]_i_8__0_n_0 ;
  wire \block_w2_reg[14]_i_8_n_0 ;
  wire \block_w2_reg[15]_i_12_n_0 ;
  wire \block_w2_reg[15]_i_6__0_n_0 ;
  wire \block_w2_reg[15]_i_7_n_0 ;
  wire \block_w2_reg[15]_i_8_n_0 ;
  wire \block_w2_reg[16]_i_11_n_0 ;
  wire \block_w2_reg[16]_i_5_n_0 ;
  wire \block_w2_reg[16]_i_6__0_n_0 ;
  wire \block_w2_reg[16]_i_6_n_0 ;
  wire \block_w2_reg[16]_i_7__0_n_0 ;
  wire \block_w2_reg[16]_i_7_n_0 ;
  wire \block_w2_reg[16]_i_8_n_0 ;
  wire \block_w2_reg[17]_i_12_n_0 ;
  wire \block_w2_reg[17]_i_7_n_0 ;
  wire \block_w2_reg[17]_i_8_n_0 ;
  wire \block_w2_reg[17]_i_9_n_0 ;
  wire \block_w2_reg[18]_i_11_n_0 ;
  wire \block_w2_reg[18]_i_6__0_n_0 ;
  wire \block_w2_reg[18]_i_6_n_0 ;
  wire \block_w2_reg[18]_i_7__0_n_0 ;
  wire \block_w2_reg[18]_i_7_n_0 ;
  wire \block_w2_reg[18]_i_8_n_0 ;
  wire \block_w2_reg[19]_i_12_n_0 ;
  wire \block_w2_reg[19]_i_6_n_0 ;
  wire \block_w2_reg[19]_i_7__0_n_0 ;
  wire \block_w2_reg[19]_i_8__0_n_0 ;
  wire \block_w2_reg[19]_i_9_n_0 ;
  wire \block_w2_reg[1]_i_12_n_0 ;
  wire \block_w2_reg[1]_i_7_n_0 ;
  wire \block_w2_reg[1]_i_8_n_0 ;
  wire \block_w2_reg[1]_i_9_n_0 ;
  wire \block_w2_reg[20]_i_10_n_0 ;
  wire \block_w2_reg[20]_i_13_n_0 ;
  wire \block_w2_reg[20]_i_8_n_0 ;
  wire \block_w2_reg[20]_i_9_n_0 ;
  wire \block_w2_reg[21]_i_11_n_0 ;
  wire \block_w2_reg[21]_i_6__0_n_0 ;
  wire \block_w2_reg[21]_i_7__0_n_0 ;
  wire \block_w2_reg[21]_i_7_n_0 ;
  wire \block_w2_reg[21]_i_8__0_n_0 ;
  wire \block_w2_reg[21]_i_8_n_0 ;
  wire \block_w2_reg[22]_i_11_n_0 ;
  wire \block_w2_reg[22]_i_6__0_n_0 ;
  wire \block_w2_reg[22]_i_7__0_n_0 ;
  wire \block_w2_reg[22]_i_7_n_0 ;
  wire \block_w2_reg[22]_i_8_n_0 ;
  wire \block_w2_reg[23]_i_12_n_0 ;
  wire \block_w2_reg[23]_i_6__0_n_0 ;
  wire \block_w2_reg[23]_i_7__0_n_0 ;
  wire \block_w2_reg[23]_i_7_n_0 ;
  wire \block_w2_reg[23]_i_8_n_0 ;
  wire \block_w2_reg[24]_i_11_n_0 ;
  wire \block_w2_reg[24]_i_6__0_n_0 ;
  wire \block_w2_reg[24]_i_7__0_n_0 ;
  wire \block_w2_reg[24]_i_7_n_0 ;
  wire \block_w2_reg[24]_i_8__0_n_0 ;
  wire \block_w2_reg[24]_i_8_n_0 ;
  wire \block_w2_reg[24]_i_9_n_0 ;
  wire \block_w2_reg[25]_i_10_n_0 ;
  wire \block_w2_reg[25]_i_13_n_0 ;
  wire \block_w2_reg[25]_i_8_n_0 ;
  wire \block_w2_reg[25]_i_9_n_0 ;
  wire \block_w2_reg[26]_i_11_n_0 ;
  wire \block_w2_reg[26]_i_6__0_n_0 ;
  wire \block_w2_reg[26]_i_6_n_0 ;
  wire \block_w2_reg[26]_i_7_n_0 ;
  wire \block_w2_reg[26]_i_8_n_0 ;
  wire \block_w2_reg[27]_i_10_n_0 ;
  wire \block_w2_reg[27]_i_14_n_0 ;
  wire \block_w2_reg[27]_i_6_n_0 ;
  wire \block_w2_reg[27]_i_7_n_0 ;
  wire \block_w2_reg[27]_i_9_n_0 ;
  wire \block_w2_reg[28]_i_13_n_0 ;
  wire \block_w2_reg[28]_i_6__0_n_0 ;
  wire \block_w2_reg[28]_i_7__0_n_0 ;
  wire \block_w2_reg[28]_i_7_n_0 ;
  wire \block_w2_reg[28]_i_8_n_0 ;
  wire \block_w2_reg[28]_i_9_n_0 ;
  wire \block_w2_reg[29]_i_11_n_0 ;
  wire \block_w2_reg[29]_i_4_0 ;
  wire \block_w2_reg[29]_i_4_1 ;
  wire \block_w2_reg[29]_i_6__0_n_0 ;
  wire \block_w2_reg[29]_i_7__0_n_0 ;
  wire \block_w2_reg[29]_i_7_n_0 ;
  wire \block_w2_reg[29]_i_8__0_n_0 ;
  wire \block_w2_reg[29]_i_8_n_0 ;
  wire \block_w2_reg[2]_i_11_n_0 ;
  wire \block_w2_reg[2]_i_6__0_n_0 ;
  wire \block_w2_reg[2]_i_7__0_n_0 ;
  wire \block_w2_reg[2]_i_7_n_0 ;
  wire \block_w2_reg[2]_i_8_n_0 ;
  wire \block_w2_reg[30]_i_11_n_0 ;
  wire \block_w2_reg[30]_i_6__0_n_0 ;
  wire \block_w2_reg[30]_i_7__0_n_0 ;
  wire \block_w2_reg[30]_i_7_n_0 ;
  wire \block_w2_reg[30]_i_8__0_n_0 ;
  wire \block_w2_reg[30]_i_8_n_0 ;
  wire \block_w2_reg[31]_i_11_n_0 ;
  wire \block_w2_reg[31]_i_13_n_0 ;
  wire \block_w2_reg[31]_i_15_n_0 ;
  wire \block_w2_reg[31]_i_19_n_0 ;
  wire \block_w2_reg[31]_i_21_n_0 ;
  wire \block_w2_reg[3]_i_12_n_0 ;
  wire \block_w2_reg[3]_i_6__0_n_0 ;
  wire \block_w2_reg[3]_i_7__0_n_0 ;
  wire \block_w2_reg[3]_i_7_n_0 ;
  wire \block_w2_reg[3]_i_8__0_n_0 ;
  wire \block_w2_reg[3]_i_8_n_0 ;
  wire \block_w2_reg[3]_i_9_n_0 ;
  wire \block_w2_reg[4]_i_10_n_0 ;
  wire \block_w2_reg[4]_i_13_n_0 ;
  wire \block_w2_reg[4]_i_8_n_0 ;
  wire \block_w2_reg[4]_i_9_n_0 ;
  wire \block_w2_reg[5]_i_11_n_0 ;
  wire \block_w2_reg[5]_i_6__0_n_0 ;
  wire \block_w2_reg[5]_i_7__0_n_0 ;
  wire \block_w2_reg[5]_i_7_n_0 ;
  wire \block_w2_reg[5]_i_8__0_n_0 ;
  wire \block_w2_reg[5]_i_8_n_0 ;
  wire \block_w2_reg[6]_i_11_n_0 ;
  wire \block_w2_reg[6]_i_6__0_n_0 ;
  wire \block_w2_reg[6]_i_7__0_n_0 ;
  wire \block_w2_reg[6]_i_7_n_0 ;
  wire \block_w2_reg[6]_i_8_n_0 ;
  wire \block_w2_reg[7]_i_12_n_0 ;
  wire \block_w2_reg[7]_i_4_n_0 ;
  wire \block_w2_reg[7]_i_6__0_n_0 ;
  wire \block_w2_reg[7]_i_7__0_n_0 ;
  wire \block_w2_reg[7]_i_7_n_0 ;
  wire \block_w2_reg[7]_i_8_n_0 ;
  wire \block_w2_reg[8]_i_11_n_0 ;
  wire \block_w2_reg[8]_i_6__0_n_0 ;
  wire \block_w2_reg[8]_i_7__0_n_0 ;
  wire \block_w2_reg[8]_i_7_n_0 ;
  wire \block_w2_reg[8]_i_8__0_n_0 ;
  wire \block_w2_reg[8]_i_8_n_0 ;
  wire \block_w2_reg[9]_i_10_n_0 ;
  wire \block_w2_reg[9]_i_13_n_0 ;
  wire \block_w2_reg[9]_i_5_n_0 ;
  wire \block_w2_reg[9]_i_6_n_0 ;
  wire \block_w2_reg[9]_i_8_n_0 ;
  wire \block_w2_reg[9]_i_9_n_0 ;
  wire [0:0]\block_w2_reg_reg[0] ;
  wire \block_w2_reg_reg[0]_0 ;
  wire \block_w2_reg_reg[10] ;
  wire \block_w2_reg_reg[12] ;
  wire \block_w2_reg_reg[13] ;
  wire \block_w2_reg_reg[14] ;
  wire \block_w2_reg_reg[15] ;
  wire [0:0]\block_w2_reg_reg[16] ;
  wire \block_w2_reg_reg[17] ;
  wire \block_w2_reg_reg[19] ;
  wire \block_w2_reg_reg[1] ;
  wire \block_w2_reg_reg[20] ;
  wire \block_w2_reg_reg[21] ;
  wire \block_w2_reg_reg[22] ;
  wire \block_w2_reg_reg[23] ;
  wire \block_w2_reg_reg[24] ;
  wire \block_w2_reg_reg[25] ;
  wire \block_w2_reg_reg[28] ;
  wire \block_w2_reg_reg[29] ;
  wire \block_w2_reg_reg[2] ;
  wire \block_w2_reg_reg[30] ;
  wire \block_w2_reg_reg[31] ;
  wire \block_w2_reg_reg[31]_0 ;
  wire \block_w2_reg_reg[3] ;
  wire \block_w2_reg_reg[4] ;
  wire \block_w2_reg_reg[5] ;
  wire \block_w2_reg_reg[6] ;
  wire \block_w2_reg_reg[7] ;
  wire \block_w2_reg_reg[8] ;
  wire [0:0]\block_w2_reg_reg[9] ;
  wire \block_w3_reg[0]_i_5__0_n_0 ;
  wire \block_w3_reg[0]_i_6__0_n_0 ;
  wire \block_w3_reg[0]_i_6_n_0 ;
  wire \block_w3_reg[0]_i_7__0_n_0 ;
  wire \block_w3_reg[0]_i_7_n_0 ;
  wire \block_w3_reg[0]_i_8_n_0 ;
  wire \block_w3_reg[10]_i_10_n_0 ;
  wire \block_w3_reg[10]_i_5__0_n_0 ;
  wire \block_w3_reg[10]_i_6_n_0 ;
  wire \block_w3_reg[10]_i_7__0_n_0 ;
  wire \block_w3_reg[10]_i_8_n_0 ;
  wire \block_w3_reg[11]_i_10_n_0 ;
  wire \block_w3_reg[11]_i_6_n_0 ;
  wire \block_w3_reg[11]_i_7_n_0 ;
  wire \block_w3_reg[11]_i_8__0_n_0 ;
  wire \block_w3_reg[11]_i_8_n_0 ;
  wire \block_w3_reg[11]_i_9__0_n_0 ;
  wire \block_w3_reg[11]_i_9_n_0 ;
  wire \block_w3_reg[12]_i_10_n_0 ;
  wire \block_w3_reg[12]_i_11_n_0 ;
  wire \block_w3_reg[12]_i_12_n_0 ;
  wire \block_w3_reg[12]_i_13_n_0 ;
  wire \block_w3_reg[12]_i_6__0_n_0 ;
  wire \block_w3_reg[12]_i_7_n_0 ;
  wire \block_w3_reg[12]_i_8_n_0 ;
  wire \block_w3_reg[12]_i_9__0_n_0 ;
  wire \block_w3_reg[12]_i_9_n_0 ;
  wire \block_w3_reg[13]_i_10_n_0 ;
  wire \block_w3_reg[13]_i_11_n_0 ;
  wire \block_w3_reg[13]_i_12_n_0 ;
  wire \block_w3_reg[13]_i_13_n_0 ;
  wire \block_w3_reg[13]_i_14_n_0 ;
  wire \block_w3_reg[13]_i_5__0_n_0 ;
  wire \block_w3_reg[13]_i_6_n_0 ;
  wire \block_w3_reg[13]_i_7__0_n_0 ;
  wire \block_w3_reg[13]_i_8_n_0 ;
  wire \block_w3_reg[14]_i_10_n_0 ;
  wire \block_w3_reg[14]_i_11_n_0 ;
  wire \block_w3_reg[14]_i_12_n_0 ;
  wire \block_w3_reg[14]_i_13_n_0 ;
  wire \block_w3_reg[14]_i_14_n_0 ;
  wire \block_w3_reg[14]_i_5__0_n_0 ;
  wire \block_w3_reg[14]_i_6_n_0 ;
  wire \block_w3_reg[14]_i_7__0_n_0 ;
  wire \block_w3_reg[14]_i_8_n_0 ;
  wire \block_w3_reg[15]_i_11_n_0 ;
  wire \block_w3_reg[15]_i_12_n_0 ;
  wire \block_w3_reg[15]_i_5__0_n_0 ;
  wire \block_w3_reg[15]_i_6_n_0 ;
  wire \block_w3_reg[15]_i_7__0_n_0 ;
  wire \block_w3_reg[15]_i_8_n_0 ;
  wire \block_w3_reg[16]_i_5_n_0 ;
  wire \block_w3_reg[16]_i_6__0_n_0 ;
  wire \block_w3_reg[16]_i_6_n_0 ;
  wire \block_w3_reg[16]_i_7__0_n_0 ;
  wire \block_w3_reg[16]_i_7_n_0 ;
  wire \block_w3_reg[16]_i_8__0_n_0 ;
  wire \block_w3_reg[16]_i_8_n_0 ;
  wire \block_w3_reg[17]_i_6__0_n_0 ;
  wire \block_w3_reg[17]_i_7_n_0 ;
  wire \block_w3_reg[17]_i_8_n_0 ;
  wire \block_w3_reg[17]_i_9__0_n_0 ;
  wire \block_w3_reg[17]_i_9_n_0 ;
  wire \block_w3_reg[18]_i_10_n_0 ;
  wire \block_w3_reg[18]_i_5_n_0 ;
  wire \block_w3_reg[18]_i_6__0_n_0 ;
  wire \block_w3_reg[18]_i_7_n_0 ;
  wire \block_w3_reg[18]_i_8_n_0 ;
  wire \block_w3_reg[18]_i_9_n_0 ;
  wire \block_w3_reg[19]_i_10__0_n_0 ;
  wire \block_w3_reg[19]_i_10_n_0 ;
  wire \block_w3_reg[19]_i_11_n_0 ;
  wire \block_w3_reg[19]_i_6__0_n_0 ;
  wire \block_w3_reg[19]_i_7_n_0 ;
  wire \block_w3_reg[19]_i_8_n_0 ;
  wire \block_w3_reg[19]_i_9_n_0 ;
  wire \block_w3_reg[1]_i_4__0_0 ;
  wire \block_w3_reg[1]_i_6__0_n_0 ;
  wire \block_w3_reg[1]_i_7_n_0 ;
  wire \block_w3_reg[1]_i_8_n_0 ;
  wire \block_w3_reg[1]_i_9__0_n_0 ;
  wire \block_w3_reg[1]_i_9_n_0 ;
  wire \block_w3_reg[20]_i_10__0_n_0 ;
  wire \block_w3_reg[20]_i_10_n_0 ;
  wire \block_w3_reg[20]_i_11_n_0 ;
  wire \block_w3_reg[20]_i_7_n_0 ;
  wire \block_w3_reg[20]_i_8_n_0 ;
  wire \block_w3_reg[20]_i_9__0_n_0 ;
  wire \block_w3_reg[20]_i_9_n_0 ;
  wire \block_w3_reg[21]_i_10_n_0 ;
  wire \block_w3_reg[21]_i_11_n_0 ;
  wire \block_w3_reg[21]_i_12_n_0 ;
  wire \block_w3_reg[21]_i_13_n_0 ;
  wire \block_w3_reg[21]_i_14_n_0 ;
  wire \block_w3_reg[21]_i_5__0_n_0 ;
  wire \block_w3_reg[21]_i_6_n_0 ;
  wire \block_w3_reg[21]_i_7__0_n_0 ;
  wire \block_w3_reg[21]_i_8_n_0 ;
  wire \block_w3_reg[22]_i_10_n_0 ;
  wire \block_w3_reg[22]_i_11_n_0 ;
  wire \block_w3_reg[22]_i_12_n_0 ;
  wire \block_w3_reg[22]_i_13_n_0 ;
  wire \block_w3_reg[22]_i_14_n_0 ;
  wire \block_w3_reg[22]_i_5__0_n_0 ;
  wire \block_w3_reg[22]_i_6_n_0 ;
  wire \block_w3_reg[22]_i_7__0_n_0 ;
  wire \block_w3_reg[22]_i_8_n_0 ;
  wire \block_w3_reg[23]_i_11_n_0 ;
  wire \block_w3_reg[23]_i_12_n_0 ;
  wire \block_w3_reg[23]_i_5__0_n_0 ;
  wire \block_w3_reg[23]_i_6_n_0 ;
  wire \block_w3_reg[23]_i_7__0_n_0 ;
  wire \block_w3_reg[23]_i_8_n_0 ;
  wire \block_w3_reg[24]_i_10_n_0 ;
  wire \block_w3_reg[24]_i_11_n_0 ;
  wire \block_w3_reg[24]_i_12_n_0 ;
  wire \block_w3_reg[24]_i_13_n_0 ;
  wire \block_w3_reg[24]_i_5__0_n_0 ;
  wire \block_w3_reg[24]_i_6_n_0 ;
  wire \block_w3_reg[24]_i_7__0_n_0 ;
  wire \block_w3_reg[24]_i_8_n_0 ;
  wire \block_w3_reg[25]_i_10_n_0 ;
  wire \block_w3_reg[25]_i_11_n_0 ;
  wire \block_w3_reg[25]_i_7_n_0 ;
  wire \block_w3_reg[25]_i_9__0_n_0 ;
  wire \block_w3_reg[25]_i_9_n_0 ;
  wire \block_w3_reg[26]_i_5_n_0 ;
  wire \block_w3_reg[26]_i_6__0_n_0 ;
  wire \block_w3_reg[26]_i_7_n_0 ;
  wire \block_w3_reg[26]_i_8_n_0 ;
  wire \block_w3_reg[26]_i_9_n_0 ;
  wire \block_w3_reg[27]_i_10__0_n_0 ;
  wire \block_w3_reg[27]_i_10_n_0 ;
  wire \block_w3_reg[27]_i_6_n_0 ;
  wire \block_w3_reg[27]_i_7_n_0 ;
  wire \block_w3_reg[27]_i_8__0_n_0 ;
  wire \block_w3_reg[27]_i_8_n_0 ;
  wire \block_w3_reg[28]_i_10__0_n_0 ;
  wire \block_w3_reg[28]_i_10_n_0 ;
  wire \block_w3_reg[28]_i_11_n_0 ;
  wire \block_w3_reg[28]_i_12_n_0 ;
  wire \block_w3_reg[28]_i_6__0_n_0 ;
  wire \block_w3_reg[28]_i_7_n_0 ;
  wire \block_w3_reg[28]_i_8_n_0 ;
  wire \block_w3_reg[28]_i_9_n_0 ;
  wire \block_w3_reg[29]_i_10_n_0 ;
  wire \block_w3_reg[29]_i_11_n_0 ;
  wire \block_w3_reg[29]_i_12_n_0 ;
  wire \block_w3_reg[29]_i_13_n_0 ;
  wire \block_w3_reg[29]_i_14_n_0 ;
  wire \block_w3_reg[29]_i_5__0_n_0 ;
  wire \block_w3_reg[29]_i_6_n_0 ;
  wire \block_w3_reg[29]_i_7__0_n_0 ;
  wire \block_w3_reg[29]_i_8_n_0 ;
  wire \block_w3_reg[2]_i_10_n_0 ;
  wire \block_w3_reg[2]_i_11_n_0 ;
  wire \block_w3_reg[2]_i_12_n_0 ;
  wire \block_w3_reg[2]_i_5__0_n_0 ;
  wire \block_w3_reg[2]_i_6_n_0 ;
  wire \block_w3_reg[2]_i_7__0_n_0 ;
  wire \block_w3_reg[2]_i_8_n_0 ;
  wire \block_w3_reg[30]_i_10_n_0 ;
  wire \block_w3_reg[30]_i_11_n_0 ;
  wire \block_w3_reg[30]_i_12_n_0 ;
  wire \block_w3_reg[30]_i_13_n_0 ;
  wire \block_w3_reg[30]_i_14_n_0 ;
  wire \block_w3_reg[30]_i_4_0 ;
  wire \block_w3_reg[30]_i_4_1 ;
  wire \block_w3_reg[30]_i_5__0_n_0 ;
  wire \block_w3_reg[30]_i_6_n_0 ;
  wire \block_w3_reg[30]_i_7__0_n_0 ;
  wire \block_w3_reg[30]_i_8_n_0 ;
  wire \block_w3_reg[31]_i_13_n_0 ;
  wire \block_w3_reg[31]_i_14_n_0 ;
  wire \block_w3_reg[31]_i_6__0_n_0 ;
  wire \block_w3_reg[31]_i_7__0_n_0 ;
  wire \block_w3_reg[31]_i_8_n_0 ;
  wire \block_w3_reg[31]_i_9__0_n_0 ;
  wire \block_w3_reg[3]_i_10_n_0 ;
  wire \block_w3_reg[3]_i_11_n_0 ;
  wire \block_w3_reg[3]_i_12_n_0 ;
  wire \block_w3_reg[3]_i_13_n_0 ;
  wire \block_w3_reg[3]_i_6__0_n_0 ;
  wire \block_w3_reg[3]_i_7_n_0 ;
  wire \block_w3_reg[3]_i_8_n_0 ;
  wire \block_w3_reg[3]_i_9__0_n_0 ;
  wire \block_w3_reg[3]_i_9_n_0 ;
  wire \block_w3_reg[4]_i_10__0_n_0 ;
  wire \block_w3_reg[4]_i_10_n_0 ;
  wire \block_w3_reg[4]_i_7_n_0 ;
  wire \block_w3_reg[4]_i_8_n_0 ;
  wire \block_w3_reg[4]_i_9__0_n_0 ;
  wire \block_w3_reg[4]_i_9_n_0 ;
  wire \block_w3_reg[5]_i_10_n_0 ;
  wire \block_w3_reg[5]_i_11_n_0 ;
  wire \block_w3_reg[5]_i_12_n_0 ;
  wire \block_w3_reg[5]_i_13_n_0 ;
  wire \block_w3_reg[5]_i_14_n_0 ;
  wire \block_w3_reg[5]_i_5__0_n_0 ;
  wire \block_w3_reg[5]_i_6_n_0 ;
  wire \block_w3_reg[5]_i_7__0_n_0 ;
  wire \block_w3_reg[5]_i_8_n_0 ;
  wire \block_w3_reg[6]_i_10_n_0 ;
  wire \block_w3_reg[6]_i_11_n_0 ;
  wire \block_w3_reg[6]_i_12_n_0 ;
  wire \block_w3_reg[6]_i_13_n_0 ;
  wire \block_w3_reg[6]_i_14_n_0 ;
  wire \block_w3_reg[6]_i_5__0_n_0 ;
  wire \block_w3_reg[6]_i_6_n_0 ;
  wire \block_w3_reg[6]_i_7__0_n_0 ;
  wire \block_w3_reg[6]_i_8_n_0 ;
  wire \block_w3_reg[7]_i_11_n_0 ;
  wire \block_w3_reg[7]_i_12_n_0 ;
  wire \block_w3_reg[7]_i_4_n_0 ;
  wire \block_w3_reg[7]_i_5__0_n_0 ;
  wire \block_w3_reg[7]_i_6_n_0 ;
  wire \block_w3_reg[7]_i_7__0_n_0 ;
  wire \block_w3_reg[7]_i_8_n_0 ;
  wire \block_w3_reg[8]_i_10_n_0 ;
  wire \block_w3_reg[8]_i_11_n_0 ;
  wire \block_w3_reg[8]_i_12_n_0 ;
  wire \block_w3_reg[8]_i_5__0_n_0 ;
  wire \block_w3_reg[8]_i_6_n_0 ;
  wire \block_w3_reg[8]_i_7__0_n_0 ;
  wire \block_w3_reg[8]_i_8_n_0 ;
  wire \block_w3_reg[9]_i_10__0_n_0 ;
  wire \block_w3_reg[9]_i_10_n_0 ;
  wire \block_w3_reg[9]_i_7_n_0 ;
  wire \block_w3_reg[9]_i_8_n_0 ;
  wire \block_w3_reg[9]_i_9__0_n_0 ;
  wire \block_w3_reg[9]_i_9_n_0 ;
  wire [0:0]\block_w3_reg_reg[0] ;
  wire \block_w3_reg_reg[0]_0 ;
  wire \block_w3_reg_reg[10] ;
  wire \block_w3_reg_reg[12] ;
  wire \block_w3_reg_reg[13] ;
  wire \block_w3_reg_reg[14] ;
  wire \block_w3_reg_reg[15] ;
  wire [0:0]\block_w3_reg_reg[16] ;
  wire \block_w3_reg_reg[17] ;
  wire \block_w3_reg_reg[19] ;
  wire \block_w3_reg_reg[1] ;
  wire \block_w3_reg_reg[20] ;
  wire \block_w3_reg_reg[21] ;
  wire \block_w3_reg_reg[22] ;
  wire \block_w3_reg_reg[23] ;
  wire \block_w3_reg_reg[24] ;
  wire \block_w3_reg_reg[25] ;
  wire \block_w3_reg_reg[26] ;
  wire \block_w3_reg_reg[28] ;
  wire \block_w3_reg_reg[29] ;
  wire \block_w3_reg_reg[2] ;
  wire \block_w3_reg_reg[30] ;
  wire \block_w3_reg_reg[31] ;
  wire \block_w3_reg_reg[31]_0 ;
  wire \block_w3_reg_reg[3] ;
  wire \block_w3_reg_reg[4] ;
  wire \block_w3_reg_reg[5] ;
  wire \block_w3_reg_reg[6] ;
  wire \block_w3_reg_reg[7] ;
  wire \block_w3_reg_reg[8] ;
  wire \block_w3_reg_reg[8]_0 ;
  wire \block_w3_reg_reg[9] ;
  wire clk_i;
  wire [127:0]core_block;
  wire [255:0]core_key;
  wire [7:0]\dec_block/op126_in ;
  wire [7:1]\dec_block/op127_in ;
  wire [7:0]\dec_block/op129_in ;
  wire [7:0]\dec_block/op158_in ;
  wire [7:1]\dec_block/op159_in ;
  wire [7:0]\dec_block/op161_in ;
  wire [7:0]\dec_block/op190_in ;
  wire [7:1]\dec_block/op191_in ;
  wire [7:0]\dec_block/op193_in ;
  wire [7:0]\dec_block/op95_in ;
  wire [7:1]\dec_block/op96_in ;
  wire [7:0]\dec_block/op98_in ;
  wire [7:2]\dec_block/p_0_in31_in ;
  wire [7:2]\dec_block/p_0_in38_in ;
  wire [7:2]\dec_block/p_0_in46_in ;
  wire [7:2]\dec_block/p_0_in54_in ;
  wire [127:0]dec_new_block;
  wire dec_ready;
  wire enc_ready;
  wire init_state;
  wire [6:0]inv_mixcolumns_return0110_out__47;
  wire [6:0]inv_mixcolumns_return0117_out__50;
  wire [7:0]inv_mixcolumns_return0124_out__47;
  wire [6:0]inv_mixcolumns_return0134_out__63;
  wire [7:0]inv_mixcolumns_return0142_out__55;
  wire [6:0]inv_mixcolumns_return0149_out__55;
  wire [7:0]inv_mixcolumns_return0156_out__63;
  wire [6:0]inv_mixcolumns_return0166_out__55;
  wire [7:0]inv_mixcolumns_return0174_out__63;
  wire [6:0]inv_mixcolumns_return0181_out__58;
  wire [7:0]inv_mixcolumns_return0188_out__55;
  wire [6:0]inv_mixcolumns_return0198_out__63;
  wire [6:0]inv_mixcolumns_return0206_out__55;
  wire [6:0]inv_mixcolumns_return0213_out__55;
  wire [7:0]inv_mixcolumns_return0220_out__63;
  wire [6:0]inv_mixcolumns_return0__55;
  wire key_mem;
  wire \key_mem[0][127]_i_3_n_0 ;
  wire \key_mem[10][127]_i_1_n_0 ;
  wire \key_mem[11][127]_i_1_n_0 ;
  wire \key_mem[12][127]_i_1_n_0 ;
  wire \key_mem[13][127]_i_1_n_0 ;
  wire \key_mem[14][127]_i_1_n_0 ;
  wire \key_mem[1][127]_i_1_n_0 ;
  wire \key_mem[2][127]_i_1_n_0 ;
  wire \key_mem[3][127]_i_1_n_0 ;
  wire \key_mem[4][127]_i_1_n_0 ;
  wire \key_mem[5][127]_i_1_n_0 ;
  wire \key_mem[6][127]_i_1_n_0 ;
  wire \key_mem[7][127]_i_1_n_0 ;
  wire \key_mem[8][127]_i_1_n_0 ;
  wire \key_mem[9][127]_i_1_n_0 ;
  wire [1:0]key_mem_ctrl_new;
  wire [1:0]key_mem_ctrl_reg;
  wire [127:0]key_mem_new;
  wire [127:0]\key_mem_reg[0]_0 ;
  wire [127:0]\key_mem_reg[10]_10 ;
  wire [127:0]\key_mem_reg[11]_11 ;
  wire [127:0]\key_mem_reg[12]_12 ;
  wire [127:0]\key_mem_reg[13]_13 ;
  wire \key_mem_reg[14][127]_0 ;
  wire \key_mem_reg[14][36]_0 ;
  wire [127:0]\key_mem_reg[14]_14 ;
  wire [127:0]\key_mem_reg[1]_1 ;
  wire [127:0]\key_mem_reg[2]_2 ;
  wire [127:0]\key_mem_reg[3]_3 ;
  wire [127:0]\key_mem_reg[4]_4 ;
  wire [127:0]\key_mem_reg[5]_5 ;
  wire [127:0]\key_mem_reg[6]_6 ;
  wire [127:0]\key_mem_reg[7]_7 ;
  wire [127:0]\key_mem_reg[8]_8 ;
  wire [127:0]\key_mem_reg[9]_9 ;
  wire key_ready;
  wire [3:0]muxed_round_nr;
  wire [31:0]new_sboxw;
  wire p_0_in;
  wire p_0_in0;
  wire [75:0]p_0_out;
  wire [31:0]p_10_in;
  wire [7:0]p_19_in;
  wire [2:0]p_1_in;
  wire [31:0]p_2_in;
  wire [31:0]p_6_in;
  wire [127:0]prev_key0_new;
  wire \prev_key0_reg[127]_i_3_n_0 ;
  wire \prev_key0_reg_reg_n_0_[0] ;
  wire \prev_key0_reg_reg_n_0_[10] ;
  wire \prev_key0_reg_reg_n_0_[11] ;
  wire \prev_key0_reg_reg_n_0_[12] ;
  wire \prev_key0_reg_reg_n_0_[13] ;
  wire \prev_key0_reg_reg_n_0_[14] ;
  wire \prev_key0_reg_reg_n_0_[15] ;
  wire \prev_key0_reg_reg_n_0_[16] ;
  wire \prev_key0_reg_reg_n_0_[17] ;
  wire \prev_key0_reg_reg_n_0_[18] ;
  wire \prev_key0_reg_reg_n_0_[19] ;
  wire \prev_key0_reg_reg_n_0_[1] ;
  wire \prev_key0_reg_reg_n_0_[20] ;
  wire \prev_key0_reg_reg_n_0_[21] ;
  wire \prev_key0_reg_reg_n_0_[22] ;
  wire \prev_key0_reg_reg_n_0_[23] ;
  wire \prev_key0_reg_reg_n_0_[24] ;
  wire \prev_key0_reg_reg_n_0_[25] ;
  wire \prev_key0_reg_reg_n_0_[26] ;
  wire \prev_key0_reg_reg_n_0_[27] ;
  wire \prev_key0_reg_reg_n_0_[28] ;
  wire \prev_key0_reg_reg_n_0_[29] ;
  wire \prev_key0_reg_reg_n_0_[2] ;
  wire \prev_key0_reg_reg_n_0_[30] ;
  wire \prev_key0_reg_reg_n_0_[31] ;
  wire \prev_key0_reg_reg_n_0_[3] ;
  wire \prev_key0_reg_reg_n_0_[4] ;
  wire \prev_key0_reg_reg_n_0_[5] ;
  wire \prev_key0_reg_reg_n_0_[6] ;
  wire \prev_key0_reg_reg_n_0_[7] ;
  wire \prev_key0_reg_reg_n_0_[8] ;
  wire \prev_key0_reg_reg_n_0_[9] ;
  wire prev_key0_we2_out;
  wire [127:0]prev_key1_new;
  wire [127:0]prev_key1_new0_in;
  wire \prev_key1_reg[0]_i_1_n_0 ;
  wire \prev_key1_reg[0]_i_4_n_0 ;
  wire \prev_key1_reg[100]_i_1_n_0 ;
  wire \prev_key1_reg[101]_i_1_n_0 ;
  wire \prev_key1_reg[102]_i_1_n_0 ;
  wire \prev_key1_reg[103]_i_1_n_0 ;
  wire \prev_key1_reg[104]_i_1_n_0 ;
  wire \prev_key1_reg[105]_i_1_n_0 ;
  wire \prev_key1_reg[106]_i_1_n_0 ;
  wire \prev_key1_reg[107]_i_1_n_0 ;
  wire \prev_key1_reg[108]_i_1_n_0 ;
  wire \prev_key1_reg[109]_i_1_n_0 ;
  wire \prev_key1_reg[10]_i_1_n_0 ;
  wire \prev_key1_reg[10]_i_4_n_0 ;
  wire \prev_key1_reg[110]_i_1_n_0 ;
  wire \prev_key1_reg[111]_i_1_n_0 ;
  wire \prev_key1_reg[112]_i_1_n_0 ;
  wire \prev_key1_reg[113]_i_1_n_0 ;
  wire \prev_key1_reg[114]_i_1_n_0 ;
  wire \prev_key1_reg[115]_i_1_n_0 ;
  wire \prev_key1_reg[116]_i_1_n_0 ;
  wire \prev_key1_reg[117]_i_1_n_0 ;
  wire \prev_key1_reg[118]_i_1_n_0 ;
  wire \prev_key1_reg[119]_i_1_n_0 ;
  wire \prev_key1_reg[11]_i_1_n_0 ;
  wire \prev_key1_reg[11]_i_4_n_0 ;
  wire \prev_key1_reg[120]_i_1_n_0 ;
  wire \prev_key1_reg[121]_i_1_n_0 ;
  wire \prev_key1_reg[122]_i_1_n_0 ;
  wire \prev_key1_reg[123]_i_1_n_0 ;
  wire \prev_key1_reg[124]_i_1_n_0 ;
  wire \prev_key1_reg[125]_i_1_n_0 ;
  wire \prev_key1_reg[126]_i_1_n_0 ;
  wire \prev_key1_reg[127]_i_2_n_0 ;
  wire \prev_key1_reg[127]_i_4_n_0 ;
  wire \prev_key1_reg[12]_i_1_n_0 ;
  wire \prev_key1_reg[12]_i_4_n_0 ;
  wire \prev_key1_reg[13]_i_1_n_0 ;
  wire \prev_key1_reg[13]_i_4_n_0 ;
  wire \prev_key1_reg[14]_i_1_n_0 ;
  wire \prev_key1_reg[14]_i_4_n_0 ;
  wire \prev_key1_reg[15]_i_1_n_0 ;
  wire \prev_key1_reg[15]_i_4_n_0 ;
  wire \prev_key1_reg[16]_i_1_n_0 ;
  wire \prev_key1_reg[16]_i_4_n_0 ;
  wire \prev_key1_reg[17]_i_1_n_0 ;
  wire \prev_key1_reg[17]_i_4_n_0 ;
  wire \prev_key1_reg[18]_i_1_n_0 ;
  wire \prev_key1_reg[18]_i_4_n_0 ;
  wire \prev_key1_reg[19]_i_1_n_0 ;
  wire \prev_key1_reg[19]_i_4_n_0 ;
  wire \prev_key1_reg[1]_i_1_n_0 ;
  wire \prev_key1_reg[1]_i_4_n_0 ;
  wire \prev_key1_reg[20]_i_1_n_0 ;
  wire \prev_key1_reg[20]_i_4_n_0 ;
  wire \prev_key1_reg[21]_i_1_n_0 ;
  wire \prev_key1_reg[21]_i_4_n_0 ;
  wire \prev_key1_reg[22]_i_1_n_0 ;
  wire \prev_key1_reg[22]_i_4_n_0 ;
  wire \prev_key1_reg[23]_i_1_n_0 ;
  wire \prev_key1_reg[23]_i_4_n_0 ;
  wire \prev_key1_reg[24]_i_1_n_0 ;
  wire \prev_key1_reg[24]_i_4_n_0 ;
  wire \prev_key1_reg[25]_i_1_n_0 ;
  wire \prev_key1_reg[25]_i_4_n_0 ;
  wire \prev_key1_reg[26]_i_1_n_0 ;
  wire \prev_key1_reg[26]_i_4_n_0 ;
  wire \prev_key1_reg[27]_i_1_n_0 ;
  wire \prev_key1_reg[27]_i_4_n_0 ;
  wire \prev_key1_reg[28]_i_1_n_0 ;
  wire \prev_key1_reg[28]_i_4_n_0 ;
  wire \prev_key1_reg[29]_i_1_n_0 ;
  wire \prev_key1_reg[29]_i_4_n_0 ;
  wire \prev_key1_reg[2]_i_1_n_0 ;
  wire \prev_key1_reg[2]_i_4_n_0 ;
  wire \prev_key1_reg[30]_i_1_n_0 ;
  wire \prev_key1_reg[30]_i_4_n_0 ;
  wire \prev_key1_reg[31]_i_1_n_0 ;
  wire \prev_key1_reg[31]_i_4_n_0 ;
  wire \prev_key1_reg[32]_i_1_n_0 ;
  wire \prev_key1_reg[33]_i_1_n_0 ;
  wire \prev_key1_reg[34]_i_1_n_0 ;
  wire \prev_key1_reg[35]_i_1_n_0 ;
  wire \prev_key1_reg[36]_i_1_n_0 ;
  wire \prev_key1_reg[37]_i_1_n_0 ;
  wire \prev_key1_reg[38]_i_1_n_0 ;
  wire \prev_key1_reg[39]_i_1_n_0 ;
  wire \prev_key1_reg[3]_i_1_n_0 ;
  wire \prev_key1_reg[3]_i_4_n_0 ;
  wire \prev_key1_reg[40]_i_1_n_0 ;
  wire \prev_key1_reg[41]_i_1_n_0 ;
  wire \prev_key1_reg[42]_i_1_n_0 ;
  wire \prev_key1_reg[43]_i_1_n_0 ;
  wire \prev_key1_reg[44]_i_1_n_0 ;
  wire \prev_key1_reg[45]_i_1_n_0 ;
  wire \prev_key1_reg[46]_i_1_n_0 ;
  wire \prev_key1_reg[47]_i_1_n_0 ;
  wire \prev_key1_reg[48]_i_1_n_0 ;
  wire \prev_key1_reg[49]_i_1_n_0 ;
  wire \prev_key1_reg[4]_i_1_n_0 ;
  wire \prev_key1_reg[4]_i_4_n_0 ;
  wire \prev_key1_reg[50]_i_1_n_0 ;
  wire \prev_key1_reg[51]_i_1_n_0 ;
  wire \prev_key1_reg[52]_i_1_n_0 ;
  wire \prev_key1_reg[53]_i_1_n_0 ;
  wire \prev_key1_reg[54]_i_1_n_0 ;
  wire \prev_key1_reg[55]_i_1_n_0 ;
  wire \prev_key1_reg[56]_i_1_n_0 ;
  wire \prev_key1_reg[57]_i_1_n_0 ;
  wire \prev_key1_reg[58]_i_1_n_0 ;
  wire \prev_key1_reg[59]_i_1_n_0 ;
  wire \prev_key1_reg[5]_i_1_n_0 ;
  wire \prev_key1_reg[5]_i_4_n_0 ;
  wire \prev_key1_reg[60]_i_1_n_0 ;
  wire \prev_key1_reg[61]_i_1_n_0 ;
  wire \prev_key1_reg[62]_i_1_n_0 ;
  wire \prev_key1_reg[63]_i_1_n_0 ;
  wire \prev_key1_reg[64]_i_1_n_0 ;
  wire \prev_key1_reg[65]_i_1_n_0 ;
  wire \prev_key1_reg[66]_i_1_n_0 ;
  wire \prev_key1_reg[67]_i_1_n_0 ;
  wire \prev_key1_reg[68]_i_1_n_0 ;
  wire \prev_key1_reg[69]_i_1_n_0 ;
  wire \prev_key1_reg[6]_i_1_n_0 ;
  wire \prev_key1_reg[6]_i_4_n_0 ;
  wire \prev_key1_reg[70]_i_1_n_0 ;
  wire \prev_key1_reg[71]_i_1_n_0 ;
  wire \prev_key1_reg[72]_i_1_n_0 ;
  wire \prev_key1_reg[73]_i_1_n_0 ;
  wire \prev_key1_reg[74]_i_1_n_0 ;
  wire \prev_key1_reg[75]_i_1_n_0 ;
  wire \prev_key1_reg[76]_i_1_n_0 ;
  wire \prev_key1_reg[77]_i_1_n_0 ;
  wire \prev_key1_reg[78]_i_1_n_0 ;
  wire \prev_key1_reg[79]_i_1_n_0 ;
  wire \prev_key1_reg[7]_i_1_n_0 ;
  wire \prev_key1_reg[7]_i_4_n_0 ;
  wire \prev_key1_reg[80]_i_1_n_0 ;
  wire \prev_key1_reg[81]_i_1_n_0 ;
  wire \prev_key1_reg[82]_i_1_n_0 ;
  wire \prev_key1_reg[83]_i_1_n_0 ;
  wire \prev_key1_reg[84]_i_1_n_0 ;
  wire \prev_key1_reg[85]_i_1_n_0 ;
  wire \prev_key1_reg[86]_i_1_n_0 ;
  wire \prev_key1_reg[87]_i_1_n_0 ;
  wire \prev_key1_reg[88]_i_1_n_0 ;
  wire \prev_key1_reg[89]_i_1_n_0 ;
  wire \prev_key1_reg[8]_i_1_n_0 ;
  wire \prev_key1_reg[8]_i_4_n_0 ;
  wire \prev_key1_reg[90]_i_1_n_0 ;
  wire \prev_key1_reg[91]_i_1_n_0 ;
  wire \prev_key1_reg[92]_i_1_n_0 ;
  wire \prev_key1_reg[93]_i_1_n_0 ;
  wire \prev_key1_reg[94]_i_1_n_0 ;
  wire \prev_key1_reg[95]_i_1_n_0 ;
  wire \prev_key1_reg[96]_i_1_n_0 ;
  wire \prev_key1_reg[97]_i_1_n_0 ;
  wire \prev_key1_reg[98]_i_1_n_0 ;
  wire \prev_key1_reg[99]_i_1_n_0 ;
  wire \prev_key1_reg[9]_i_1_n_0 ;
  wire \prev_key1_reg[9]_i_4_n_0 ;
  wire prev_key1_we1_out;
  wire [7:0]rcon_new;
  wire \rcon_reg[7]_i_1_n_0 ;
  wire [7:0]\rcon_reg_reg[7]_0 ;
  wire ready_new;
  wire ready_reg_i_1__1_n_0;
  wire [1:0]ready_reg_reg_0;
  wire [3:0]round_ctr_new;
  wire \round_ctr_reg[0]_rep_i_1__0_n_0 ;
  wire \round_ctr_reg[0]_rep_i_1__1_n_0 ;
  wire \round_ctr_reg[0]_rep_i_1_n_0 ;
  wire \round_ctr_reg[3]_i_3__1_n_0 ;
  wire \round_ctr_reg[3]_i_4__0_n_0 ;
  wire \round_ctr_reg_reg[0]_rep__0_n_0 ;
  wire \round_ctr_reg_reg[0]_rep__1_n_0 ;
  wire \round_ctr_reg_reg[0]_rep_n_0 ;
  wire \round_ctr_reg_reg_n_0_[0] ;
  wire \round_ctr_reg_reg_n_0_[2] ;
  wire \round_ctr_reg_reg_n_0_[3] ;
  wire round_ctr_we;
  wire [127:0]round_key;
  wire rst_i;
  wire [31:0]w0;
  wire [31:0]w1;
  wire [31:0]w2;
  wire [31:0]w4;
  wire [31:0]w5;
  wire [31:0]w6;

  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \FSM_sequential_key_mem_ctrl_reg[0]_i_1 
       (.I0(p_1_in[0]),
        .I1(key_mem_ctrl_reg[1]),
        .I2(p_0_in),
        .I3(key_mem_ctrl_reg[0]),
        .O(key_mem_ctrl_new[0]));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \FSM_sequential_key_mem_ctrl_reg[1]_i_1 
       (.I0(key_mem_ctrl_reg[0]),
        .I1(p_1_in[0]),
        .I2(key_mem_ctrl_reg[1]),
        .I3(p_0_in),
        .O(\FSM_sequential_key_mem_ctrl_reg[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'h62)) 
    \FSM_sequential_key_mem_ctrl_reg[1]_i_2 
       (.I0(key_mem_ctrl_reg[0]),
        .I1(key_mem_ctrl_reg[1]),
        .I2(p_0_in),
        .O(key_mem_ctrl_new[1]));
  LUT5 #(
    .INIT(32'h20000020)) 
    \FSM_sequential_key_mem_ctrl_reg[1]_i_3 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[0] ),
        .I2(p_0_in0),
        .I3(\round_ctr_reg_reg_n_0_[2] ),
        .I4(p_1_in[2]),
        .O(p_0_in));
  (* FSM_ENCODED_STATES = "CTRL_GENERATE:10,CTRL_INIT:01,CTRL_IDLE:00,CTRL_DONE:11" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_key_mem_ctrl_reg_reg[0] 
       (.C(clk_i),
        .CE(\FSM_sequential_key_mem_ctrl_reg[1]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_ctrl_new[0]),
        .Q(key_mem_ctrl_reg[0]));
  (* FSM_ENCODED_STATES = "CTRL_GENERATE:10,CTRL_INIT:01,CTRL_IDLE:00,CTRL_DONE:11" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_key_mem_ctrl_reg_reg[1] 
       (.C(clk_i),
        .CE(\FSM_sequential_key_mem_ctrl_reg[1]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_ctrl_new[1]),
        .Q(key_mem_ctrl_reg[1]));
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT3 #(
    .INIT(8'h60)) 
    \block_w0_reg[0]_i_2__0 
       (.I0(round_key[64]),
        .I1(core_block[64]),
        .I2(\block_w0_reg_reg[0]_1 ),
        .O(\block_reg_reg[1][0] ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \block_w0_reg[0]_i_3 
       (.I0(\dec_block/op161_in [7]),
        .I1(\block_w1_reg_reg[16] ),
        .I2(\block_w2_reg[16]_i_6_n_0 ),
        .I3(\block_w0_reg[0]_i_5_n_0 ),
        .I4(\block_w0_reg_reg[0]_1 ),
        .I5(\block_w0_reg_reg[16]_0 [0]),
        .O(\block_w1_reg_reg[31]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[0]_i_3__0 
       (.I0(\block_w0_reg[0]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[0]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[0]_i_7_n_0 ),
        .O(round_key[96]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[0]_i_4 
       (.I0(\block_w0_reg[0]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[0]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[0]_i_5__0_n_0 ),
        .I5(dec_new_block[96]),
        .O(\block_w0_reg_reg[0] ));
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \block_w0_reg[0]_i_5 
       (.I0(\dec_block/op158_in [0]),
        .I1(\dec_block/op161_in [0]),
        .I2(\block_w1_reg[7]_i_4_n_0 ),
        .O(\block_w0_reg[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[0]_i_5__0 
       (.I0(\block_w0_reg[0]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [96]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [96]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [96]),
        .O(\block_w0_reg[0]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[0]_i_6 
       (.I0(\key_mem_reg[7]_7 [96]),
        .I1(\key_mem_reg[6]_6 [96]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [96]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [96]),
        .O(\block_w0_reg[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[0]_i_7 
       (.I0(\key_mem_reg[3]_3 [96]),
        .I1(\key_mem_reg[2]_2 [96]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [96]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [96]),
        .O(\block_w0_reg[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[0]_i_8 
       (.I0(\key_mem_reg[11]_11 [96]),
        .I1(\key_mem_reg[10]_10 [96]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [96]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [96]),
        .O(\block_w0_reg[0]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[10]_i_2__0 
       (.I0(\dec_block/op190_in [2]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[10] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[10]_i_3 
       (.I0(\block_w0_reg[10]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[10]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[10]_i_7_n_0 ),
        .O(round_key[106]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[10]_i_4 
       (.I0(\block_w0_reg[10]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[10]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[10]_i_5__0_n_0 ),
        .I5(dec_new_block[106]),
        .O(\dec_block/op190_in [2]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[10]_i_5 
       (.I0(round_key[42]),
        .I1(core_block[42]),
        .O(addroundkey_return[24]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[10]_i_5__0 
       (.I0(\block_w0_reg[10]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [106]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [106]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [106]),
        .O(\block_w0_reg[10]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[10]_i_6 
       (.I0(\block_w3_reg[21]_i_11_n_0 ),
        .I1(\block_w1_reg[0]_i_5_n_0 ),
        .I2(\dec_block/p_0_in38_in [2]),
        .I3(\dec_block/op127_in [7]),
        .I4(\block_w1_reg[3]_i_8_n_0 ),
        .I5(\block_w2_reg_reg[9] ),
        .O(inv_mixcolumns_return0142_out__55[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[10]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [106]),
        .I1(\key_mem_reg[6]_6 [106]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [106]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [106]),
        .O(\block_w0_reg[10]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[10]_i_7 
       (.I0(\key_mem_reg[3]_3 [106]),
        .I1(\key_mem_reg[2]_2 [106]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [106]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [106]),
        .O(\block_w0_reg[10]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[10]_i_8 
       (.I0(\key_mem_reg[11]_11 [106]),
        .I1(\key_mem_reg[10]_10 [106]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [106]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [106]),
        .O(\block_w0_reg[10]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[11]_i_3 
       (.I0(\block_w0_reg[11]_i_6_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w0_reg[11]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[11]_i_8_n_0 ),
        .O(round_key[107]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[11]_i_4__0 
       (.I0(\block_w3_reg[19]_i_9_n_0 ),
        .I1(\block_w3_reg[20]_i_10_n_0 ),
        .I2(\block_w3_reg[22]_i_14_n_0 ),
        .I3(\block_w0_reg[11]_i_5__0_n_0 ),
        .I4(\block_w3_reg[22]_i_12_n_0 ),
        .I5(\dec_block/op127_in [3]),
        .O(inv_mixcolumns_return0142_out__55[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[11]_i_5 
       (.I0(round_key[107]),
        .I1(core_block[107]),
        .O(p_0_out[56]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[11]_i_5__0 
       (.I0(\dec_block/op126_in [2]),
        .I1(\dec_block/p_0_in38_in [3]),
        .O(\block_w0_reg[11]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[11]_i_6 
       (.I0(\block_w0_reg[11]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [107]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [107]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [107]),
        .O(\block_w0_reg[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[11]_i_7 
       (.I0(\key_mem_reg[7]_7 [107]),
        .I1(\key_mem_reg[6]_6 [107]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [107]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [107]),
        .O(\block_w0_reg[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[11]_i_8 
       (.I0(\key_mem_reg[3]_3 [107]),
        .I1(\key_mem_reg[2]_2 [107]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [107]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [107]),
        .O(\block_w0_reg[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[11]_i_9 
       (.I0(\key_mem_reg[11]_11 [107]),
        .I1(\key_mem_reg[10]_10 [107]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [107]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [107]),
        .O(\block_w0_reg[11]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[12]_i_2__0 
       (.I0(\dec_block/op190_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[12] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[12]_i_3 
       (.I0(\block_w0_reg[12]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[12]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[12]_i_8_n_0 ),
        .O(round_key[108]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[12]_i_4__0 
       (.I0(\block_w0_reg[12]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[12]_i_7_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[12]_i_6__0_n_0 ),
        .I5(dec_new_block[108]),
        .O(\dec_block/op190_in [4]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[12]_i_5 
       (.I0(round_key[108]),
        .I1(core_block[108]),
        .O(p_0_out[57]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[12]_i_5__0 
       (.I0(\block_w3_reg[21]_i_10_n_0 ),
        .I1(\block_w3_reg[20]_i_10_n_0 ),
        .I2(\block_w3_reg[20]_i_11_n_0 ),
        .I3(\block_w0_reg[12]_i_6_n_0 ),
        .I4(\block_w3_reg[22]_i_10_n_0 ),
        .I5(\block_w3_reg[19]_i_11_n_0 ),
        .O(inv_mixcolumns_return0142_out__55[4]));
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w0_reg[12]_i_6 
       (.I0(\block_w2_reg[7]_i_4_n_0 ),
        .I1(round_key[43]),
        .I2(dec_new_block[43]),
        .I3(\dec_block/op129_in [4]),
        .O(\block_w0_reg[12]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[12]_i_6__0 
       (.I0(\block_w0_reg[12]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [108]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [108]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [108]),
        .O(\block_w0_reg[12]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[12]_i_7 
       (.I0(\key_mem_reg[7]_7 [108]),
        .I1(\key_mem_reg[6]_6 [108]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [108]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [108]),
        .O(\block_w0_reg[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[12]_i_8 
       (.I0(\key_mem_reg[3]_3 [108]),
        .I1(\key_mem_reg[2]_2 [108]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [108]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [108]),
        .O(\block_w0_reg[12]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[12]_i_9 
       (.I0(\key_mem_reg[11]_11 [108]),
        .I1(\key_mem_reg[10]_10 [108]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [108]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [108]),
        .O(\block_w0_reg[12]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[13]_i_2__0 
       (.I0(\dec_block/op190_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[13] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[13]_i_3 
       (.I0(\block_w0_reg[13]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[13]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[13]_i_7__0_n_0 ),
        .O(round_key[109]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[13]_i_4 
       (.I0(\block_w0_reg[13]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[13]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[13]_i_5__0_n_0 ),
        .I5(dec_new_block[109]),
        .O(\dec_block/op190_in [5]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[13]_i_5 
       (.I0(round_key[45]),
        .I1(core_block[45]),
        .O(addroundkey_return[27]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[13]_i_5__0 
       (.I0(\block_w0_reg[13]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [109]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [109]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [109]),
        .O(\block_w0_reg[13]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[13]_i_6 
       (.I0(\block_w3_reg[21]_i_10_n_0 ),
        .I1(\block_w3_reg[21]_i_11_n_0 ),
        .I2(\block_w0_reg[13]_i_7_n_0 ),
        .I3(\dec_block/op129_in [5]),
        .I4(\block_w3_reg[23]_i_12_n_0 ),
        .I5(\block_w2_reg[29]_i_8_n_0 ),
        .O(inv_mixcolumns_return0142_out__55[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[13]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [109]),
        .I1(\key_mem_reg[6]_6 [109]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [109]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [109]),
        .O(\block_w0_reg[13]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[13]_i_7 
       (.I0(\dec_block/p_0_in38_in [5]),
        .I1(\dec_block/op126_in [4]),
        .O(\block_w0_reg[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[13]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [109]),
        .I1(\key_mem_reg[2]_2 [109]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [109]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [109]),
        .O(\block_w0_reg[13]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[13]_i_8 
       (.I0(\key_mem_reg[11]_11 [109]),
        .I1(\key_mem_reg[10]_10 [109]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [109]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [109]),
        .O(\block_w0_reg[13]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[14]_i_2__0 
       (.I0(\dec_block/op190_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[14] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[14]_i_3 
       (.I0(\block_w0_reg[14]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[14]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[14]_i_7__0_n_0 ),
        .O(round_key[110]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[14]_i_4 
       (.I0(\block_w0_reg[14]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[14]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[14]_i_5__0_n_0 ),
        .I5(dec_new_block[110]),
        .O(\dec_block/op190_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[14]_i_5 
       (.I0(round_key[46]),
        .I1(core_block[46]),
        .O(addroundkey_return[28]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[14]_i_5__0 
       (.I0(\block_w0_reg[14]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [110]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [110]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [110]),
        .O(\block_w0_reg[14]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[14]_i_6 
       (.I0(\block_w3_reg[20]_i_9_n_0 ),
        .I1(\block_w3_reg[22]_i_11_n_0 ),
        .I2(\block_w3_reg[22]_i_12_n_0 ),
        .I3(\block_w0_reg[14]_i_7_n_0 ),
        .I4(\block_w2_reg[30]_i_8_n_0 ),
        .I5(\dec_block/op129_in [6]),
        .O(inv_mixcolumns_return0142_out__55[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[14]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [110]),
        .I1(\key_mem_reg[6]_6 [110]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [110]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [110]),
        .O(\block_w0_reg[14]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[14]_i_7 
       (.I0(\dec_block/p_0_in38_in [6]),
        .I1(\dec_block/op126_in [5]),
        .O(\block_w0_reg[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[14]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [110]),
        .I1(\key_mem_reg[2]_2 [110]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [110]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [110]),
        .O(\block_w0_reg[14]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[14]_i_8 
       (.I0(\key_mem_reg[11]_11 [110]),
        .I1(\key_mem_reg[10]_10 [110]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [110]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [110]),
        .O(\block_w0_reg[14]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[15]_i_2__0 
       (.I0(\dec_block/op190_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[15] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[15]_i_3 
       (.I0(\block_w0_reg[15]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[15]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[15]_i_7_n_0 ),
        .O(round_key[111]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[15]_i_4 
       (.I0(\block_w0_reg[15]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[15]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[15]_i_5__0_n_0 ),
        .I5(dec_new_block[111]),
        .O(\dec_block/op190_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[15]_i_5 
       (.I0(round_key[47]),
        .I1(core_block[47]),
        .O(addroundkey_return[29]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[15]_i_5__0 
       (.I0(\block_w0_reg[15]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [111]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [111]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [111]),
        .O(\block_w0_reg[15]_i_5__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[15]_i_6 
       (.I0(\block_w1_reg[7]_i_7_n_0 ),
        .I1(\dec_block/op126_in [6]),
        .I2(\dec_block/p_0_in38_in [7]),
        .I3(\block_w2_reg[7]_i_4_n_0 ),
        .I4(\block_w3_reg[21]_i_13_n_0 ),
        .O(inv_mixcolumns_return0142_out__55[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[15]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [111]),
        .I1(\key_mem_reg[6]_6 [111]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [111]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [111]),
        .O(\block_w0_reg[15]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[15]_i_7 
       (.I0(\key_mem_reg[3]_3 [111]),
        .I1(\key_mem_reg[2]_2 [111]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [111]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [111]),
        .O(\block_w0_reg[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[15]_i_8 
       (.I0(\key_mem_reg[11]_11 [111]),
        .I1(\key_mem_reg[10]_10 [111]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [111]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [111]),
        .O(\block_w0_reg[15]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'h60)) 
    \block_w0_reg[16]_i_2__0 
       (.I0(round_key[16]),
        .I1(core_block[16]),
        .I2(\block_w0_reg_reg[0]_1 ),
        .O(\block_reg_reg[3][16] ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \block_w0_reg[16]_i_3 
       (.I0(\block_w0_reg[16]_i_5_n_0 ),
        .I1(\block_w2_reg[0]_i_5_n_0 ),
        .I2(\block_w3_reg_reg[0] ),
        .I3(\block_w0_reg[16]_i_6_n_0 ),
        .I4(\block_w0_reg_reg[0]_1 ),
        .I5(\block_w0_reg_reg[16]_0 [2]),
        .O(\block_w3_reg_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[16]_i_3__0 
       (.I0(\block_w0_reg[16]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[16]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[16]_i_7_n_0 ),
        .O(round_key[112]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[16]_i_4 
       (.I0(\block_w0_reg[16]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[16]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[16]_i_5__0_n_0 ),
        .I5(dec_new_block[112]),
        .O(\block_w0_reg_reg[16] ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[16]_i_5 
       (.I0(\dec_block/op95_in [7]),
        .I1(\dec_block/op96_in [7]),
        .O(\block_w0_reg[16]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[16]_i_5__0 
       (.I0(\block_w0_reg[16]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [112]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [112]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [112]),
        .O(\block_w0_reg[16]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[16]_i_6 
       (.I0(\dec_block/op95_in [0]),
        .I1(\dec_block/op98_in [0]),
        .O(\block_w0_reg[16]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[16]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [112]),
        .I1(\key_mem_reg[6]_6 [112]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [112]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [112]),
        .O(\block_w0_reg[16]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[16]_i_7 
       (.I0(\key_mem_reg[3]_3 [112]),
        .I1(\key_mem_reg[2]_2 [112]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [112]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [112]),
        .O(\block_w0_reg[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[16]_i_8 
       (.I0(\key_mem_reg[11]_11 [112]),
        .I1(\key_mem_reg[10]_10 [112]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [112]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [112]),
        .O(\block_w0_reg[16]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[17]_i_2__0 
       (.I0(\dec_block/op191_in [1]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[17] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[17]_i_3 
       (.I0(\block_w0_reg[17]_i_6_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[17]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[17]_i_8_n_0 ),
        .O(round_key[113]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[17]_i_4__0 
       (.I0(\block_w0_reg[17]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[17]_i_7_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[17]_i_6_n_0 ),
        .I5(dec_new_block[113]),
        .O(\dec_block/op191_in [1]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[17]_i_5 
       (.I0(round_key[113]),
        .I1(core_block[113]),
        .O(p_0_out[61]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[17]_i_5__0 
       (.I0(\block_w3_reg_reg[16] ),
        .I1(\dec_block/p_0_in31_in [2]),
        .I2(\block_w3_reg[28]_i_9_n_0 ),
        .I3(\block_w3_reg[24]_i_13_n_0 ),
        .I4(\dec_block/op95_in [0]),
        .I5(\block_w1_reg[8]_i_7_n_0 ),
        .O(inv_mixcolumns_return0117_out__50[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[17]_i_6 
       (.I0(\block_w0_reg[17]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [113]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [113]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [113]),
        .O(\block_w0_reg[17]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[17]_i_7 
       (.I0(\key_mem_reg[7]_7 [113]),
        .I1(\key_mem_reg[6]_6 [113]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [113]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [113]),
        .O(\block_w0_reg[17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[17]_i_8 
       (.I0(\key_mem_reg[3]_3 [113]),
        .I1(\key_mem_reg[2]_2 [113]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [113]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [113]),
        .O(\block_w0_reg[17]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[17]_i_9 
       (.I0(\key_mem_reg[11]_11 [113]),
        .I1(\key_mem_reg[10]_10 [113]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [113]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [113]),
        .O(\block_w0_reg[17]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[18]_i_3 
       (.I0(\block_w0_reg[18]_i_5__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w0_reg[18]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[18]_i_7_n_0 ),
        .O(round_key[114]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[18]_i_4 
       (.I0(round_key[18]),
        .I1(core_block[18]),
        .O(addroundkey_return[16]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[18]_i_5 
       (.I0(\block_w0_reg[18]_i_6_n_0 ),
        .I1(\dec_block/p_0_in31_in [3]),
        .I2(\dec_block/op96_in [1]),
        .I3(\block_w2_reg[2]_i_7_n_0 ),
        .I4(\block_w3_reg[29]_i_10_n_0 ),
        .I5(\dec_block/op95_in [1]),
        .O(inv_mixcolumns_return0117_out__50[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[18]_i_5__0 
       (.I0(\block_w0_reg[18]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [114]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [114]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [114]),
        .O(\block_w0_reg[18]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w0_reg[18]_i_6 
       (.I0(\block_w3_reg_reg[0] ),
        .I1(\block_w3_reg_reg[16] ),
        .I2(\dec_block/op98_in [6]),
        .I3(\dec_block/op95_in [6]),
        .O(\block_w0_reg[18]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[18]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [114]),
        .I1(\key_mem_reg[6]_6 [114]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [114]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [114]),
        .O(\block_w0_reg[18]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[18]_i_7 
       (.I0(\key_mem_reg[3]_3 [114]),
        .I1(\key_mem_reg[2]_2 [114]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [114]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [114]),
        .O(\block_w0_reg[18]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[18]_i_8 
       (.I0(\key_mem_reg[11]_11 [114]),
        .I1(\key_mem_reg[10]_10 [114]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [114]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [114]),
        .O(\block_w0_reg[18]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[19]_i_2__0 
       (.I0(\dec_block/op191_in [3]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[19] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[19]_i_3 
       (.I0(\block_w0_reg[19]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w0_reg[19]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[19]_i_8__0_n_0 ),
        .O(round_key[115]));
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[19]_i_4__0 
       (.I0(round_key[115]),
        .I1(dec_new_block[115]),
        .O(\dec_block/op191_in [3]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[19]_i_5 
       (.I0(\block_w2_reg[0]_i_5_n_0 ),
        .I1(\block_w3_reg[27]_i_8_n_0 ),
        .I2(\block_w0_reg[19]_i_6_n_0 ),
        .I3(\block_w1_reg[9]_i_6__0_n_0 ),
        .I4(\block_w1_reg[12]_i_7_n_0 ),
        .O(inv_mixcolumns_return0117_out__50[2]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[19]_i_5__0 
       (.I0(round_key[115]),
        .I1(core_block[115]),
        .O(p_0_out[63]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[19]_i_6 
       (.I0(\dec_block/op96_in [2]),
        .I1(dec_new_block[11]),
        .I2(round_key[11]),
        .I3(\block_w3_reg[7]_i_4_n_0 ),
        .I4(\dec_block/op98_in [3]),
        .I5(\dec_block/op95_in [2]),
        .O(\block_w0_reg[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[19]_i_6__0 
       (.I0(\block_w0_reg[19]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [115]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [115]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [115]),
        .O(\block_w0_reg[19]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[19]_i_7 
       (.I0(\block_w3_reg[18]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[18]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[18]_i_5_n_0 ),
        .I5(dec_new_block[18]),
        .O(\dec_block/op96_in [2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[19]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [115]),
        .I1(\key_mem_reg[6]_6 [115]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [115]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [115]),
        .O(\block_w0_reg[19]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[19]_i_8 
       (.I0(\block_w3_reg[27]_i_8__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[27]_i_7_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w3_reg[27]_i_6_n_0 ),
        .I5(dec_new_block[27]),
        .O(\dec_block/op98_in [3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[19]_i_8__0 
       (.I0(\key_mem_reg[3]_3 [115]),
        .I1(\key_mem_reg[2]_2 [115]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [115]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [115]),
        .O(\block_w0_reg[19]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[19]_i_9 
       (.I0(\key_mem_reg[11]_11 [115]),
        .I1(\key_mem_reg[10]_10 [115]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [115]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [115]),
        .O(\block_w0_reg[19]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[1]_i_2__0 
       (.I0(\dec_block/p_0_in54_in [2]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[1] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[1]_i_3 
       (.I0(\block_w0_reg[1]_i_6_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[1]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[1]_i_8_n_0 ),
        .O(round_key[97]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[1]_i_4__0 
       (.I0(\block_w0_reg[1]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[1]_i_7_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[1]_i_6_n_0 ),
        .I5(dec_new_block[97]),
        .O(\dec_block/p_0_in54_in [2]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[1]_i_5 
       (.I0(round_key[97]),
        .I1(core_block[97]),
        .O(p_0_out[46]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[1]_i_5__0 
       (.I0(\block_w1_reg_reg[0] ),
        .I1(\dec_block/op159_in [1]),
        .I2(\block_w3_reg[12]_i_9_n_0 ),
        .I3(\block_w3_reg[11]_i_9_n_0 ),
        .I4(\dec_block/op161_in [0]),
        .I5(\block_w1_reg[24]_i_7_n_0 ),
        .O(inv_mixcolumns_return0166_out__55[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[1]_i_6 
       (.I0(\block_w0_reg[1]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [97]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [97]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [97]),
        .O(\block_w0_reg[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[1]_i_7 
       (.I0(\key_mem_reg[7]_7 [97]),
        .I1(\key_mem_reg[6]_6 [97]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [97]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [97]),
        .O(\block_w0_reg[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[1]_i_8 
       (.I0(\key_mem_reg[3]_3 [97]),
        .I1(\key_mem_reg[2]_2 [97]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [97]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [97]),
        .O(\block_w0_reg[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[1]_i_9 
       (.I0(\key_mem_reg[11]_11 [97]),
        .I1(\key_mem_reg[10]_10 [97]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [97]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [97]),
        .O(\block_w0_reg[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[20]_i_10 
       (.I0(\key_mem_reg[11]_11 [116]),
        .I1(\key_mem_reg[10]_10 [116]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [116]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [116]),
        .O(\block_w0_reg[20]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[20]_i_2__0 
       (.I0(\dec_block/op191_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[20] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[20]_i_3 
       (.I0(\block_w0_reg[20]_i_7_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[20]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[20]_i_9_n_0 ),
        .O(round_key[116]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[20]_i_4 
       (.I0(\block_w0_reg[20]_i_9_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[20]_i_8_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[20]_i_7_n_0 ),
        .I5(dec_new_block[116]),
        .O(\dec_block/op191_in [4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[20]_i_5__0 
       (.I0(\block_w3_reg[30]_i_10_n_0 ),
        .I1(\dec_block/p_0_in31_in [5]),
        .I2(\block_w3_reg[28]_i_9_n_0 ),
        .I3(\block_w1_reg[9]_i_6__0_n_0 ),
        .I4(\block_w3_reg[29]_i_11_n_0 ),
        .I5(\block_w3_reg[30]_i_11_n_0 ),
        .O(inv_mixcolumns_return0117_out__50[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[20]_i_6 
       (.I0(round_key[116]),
        .I1(core_block[116]),
        .O(p_0_out[64]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[20]_i_7 
       (.I0(\block_w0_reg[20]_i_10_n_0 ),
        .I1(\key_mem_reg[14]_14 [116]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [116]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [116]),
        .O(\block_w0_reg[20]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[20]_i_8 
       (.I0(\key_mem_reg[7]_7 [116]),
        .I1(\key_mem_reg[6]_6 [116]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [116]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [116]),
        .O(\block_w0_reg[20]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[20]_i_9 
       (.I0(\key_mem_reg[3]_3 [116]),
        .I1(\key_mem_reg[2]_2 [116]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [116]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [116]),
        .O(\block_w0_reg[20]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[21]_i_2__0 
       (.I0(\dec_block/op191_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[21] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[21]_i_3 
       (.I0(\block_w0_reg[21]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[21]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[21]_i_7__0_n_0 ),
        .O(round_key[117]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[21]_i_4 
       (.I0(\block_w0_reg[21]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[21]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[21]_i_5__0_n_0 ),
        .I5(dec_new_block[117]),
        .O(\dec_block/op191_in [5]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[21]_i_5 
       (.I0(round_key[21]),
        .I1(core_block[21]),
        .O(addroundkey_return[19]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[21]_i_5__0 
       (.I0(\block_w0_reg[21]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [117]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [117]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [117]),
        .O(\block_w0_reg[21]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[21]_i_6 
       (.I0(\block_w3_reg[29]_i_10_n_0 ),
        .I1(\block_w3_reg[29]_i_11_n_0 ),
        .I2(\block_w0_reg[21]_i_7_n_0 ),
        .I3(\dec_block/p_0_in31_in [6]),
        .I4(\block_w3_reg[31]_i_14_n_0 ),
        .I5(\block_w2_reg[5]_i_8_n_0 ),
        .O(inv_mixcolumns_return0117_out__50[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[21]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [117]),
        .I1(\key_mem_reg[6]_6 [117]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [117]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [117]),
        .O(\block_w0_reg[21]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[21]_i_7 
       (.I0(\dec_block/op96_in [4]),
        .I1(\dec_block/op95_in [4]),
        .O(\block_w0_reg[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[21]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [117]),
        .I1(\key_mem_reg[2]_2 [117]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [117]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [117]),
        .O(\block_w0_reg[21]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[21]_i_8 
       (.I0(\key_mem_reg[11]_11 [117]),
        .I1(\key_mem_reg[10]_10 [117]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [117]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [117]),
        .O(\block_w0_reg[21]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[22]_i_2__0 
       (.I0(\dec_block/op191_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[22] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[22]_i_3 
       (.I0(\block_w0_reg[22]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[22]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[22]_i_7__0_n_0 ),
        .O(round_key[118]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[22]_i_4 
       (.I0(\block_w0_reg[22]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[22]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[22]_i_5__0_n_0 ),
        .I5(dec_new_block[118]),
        .O(\dec_block/op191_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[22]_i_5 
       (.I0(round_key[22]),
        .I1(core_block[22]),
        .O(addroundkey_return[20]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[22]_i_5__0 
       (.I0(\block_w0_reg[22]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [118]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [118]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [118]),
        .O(\block_w0_reg[22]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[22]_i_6 
       (.I0(\block_w3_reg[28]_i_11_n_0 ),
        .I1(\block_w3_reg[30]_i_11_n_0 ),
        .I2(\block_w3_reg[30]_i_12_n_0 ),
        .I3(\block_w0_reg[22]_i_7_n_0 ),
        .I4(\block_w3_reg[24]_i_13_n_0 ),
        .I5(\dec_block/p_0_in31_in [7]),
        .O(inv_mixcolumns_return0117_out__50[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[22]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [118]),
        .I1(\key_mem_reg[6]_6 [118]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [118]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [118]),
        .O(\block_w0_reg[22]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[22]_i_7 
       (.I0(\dec_block/op95_in [5]),
        .I1(\dec_block/op96_in [5]),
        .O(\block_w0_reg[22]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[22]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [118]),
        .I1(\key_mem_reg[2]_2 [118]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [118]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [118]),
        .O(\block_w0_reg[22]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[22]_i_8 
       (.I0(\key_mem_reg[11]_11 [118]),
        .I1(\key_mem_reg[10]_10 [118]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [118]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [118]),
        .O(\block_w0_reg[22]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[23]_i_2__0 
       (.I0(\dec_block/op191_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[23] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[23]_i_3 
       (.I0(\block_w0_reg[23]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[23]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[23]_i_7_n_0 ),
        .O(round_key[119]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[23]_i_4 
       (.I0(\block_w0_reg[23]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[23]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[23]_i_5__0_n_0 ),
        .I5(dec_new_block[119]),
        .O(\dec_block/op191_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[23]_i_5 
       (.I0(round_key[23]),
        .I1(core_block[23]),
        .O(addroundkey_return[21]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[23]_i_5__0 
       (.I0(\block_w0_reg[23]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [119]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [119]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [119]),
        .O(\block_w0_reg[23]_i_5__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[23]_i_6 
       (.I0(\block_w3_reg[31]_i_13_n_0 ),
        .I1(\dec_block/op95_in [6]),
        .I2(\dec_block/op96_in [6]),
        .I3(\dec_block/op98_in [7]),
        .I4(\block_w3_reg[29]_i_13_n_0 ),
        .O(inv_mixcolumns_return0117_out__50[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[23]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [119]),
        .I1(\key_mem_reg[6]_6 [119]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [119]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [119]),
        .O(\block_w0_reg[23]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[23]_i_7 
       (.I0(\key_mem_reg[3]_3 [119]),
        .I1(\key_mem_reg[2]_2 [119]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [119]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [119]),
        .O(\block_w0_reg[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[23]_i_8 
       (.I0(\key_mem_reg[11]_11 [119]),
        .I1(\key_mem_reg[10]_10 [119]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [119]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [119]),
        .O(\block_w0_reg[23]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[24]_i_2__0 
       (.I0(\dec_block/op193_in [0]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[24] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[24]_i_3 
       (.I0(\block_w0_reg[24]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[24]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[24]_i_7_n_0 ),
        .O(round_key[120]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[24]_i_4 
       (.I0(\block_w0_reg[24]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[24]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[24]_i_5__0_n_0 ),
        .I5(dec_new_block[120]),
        .O(\dec_block/op193_in [0]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[24]_i_5 
       (.I0(round_key[120]),
        .I1(core_block[120]),
        .O(p_0_out[68]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[24]_i_5__0 
       (.I0(\block_w0_reg[24]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [120]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [120]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [120]),
        .O(\block_w0_reg[24]_i_5__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[24]_i_6 
       (.I0(\block_w2_reg[8]_i_7_n_0 ),
        .I1(\dec_block/op190_in [0]),
        .I2(\block_w3_reg[1]_i_9_n_0 ),
        .I3(\block_w3_reg[2]_i_11_n_0 ),
        .I4(\block_w3_reg[6]_i_14_n_0 ),
        .O(inv_mixcolumns_return0220_out__63[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[24]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [120]),
        .I1(\key_mem_reg[6]_6 [120]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [120]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [120]),
        .O(\block_w0_reg[24]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[24]_i_7 
       (.I0(\key_mem_reg[3]_3 [120]),
        .I1(\key_mem_reg[2]_2 [120]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [120]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [120]),
        .O(\block_w0_reg[24]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[24]_i_8 
       (.I0(\key_mem_reg[11]_11 [120]),
        .I1(\key_mem_reg[10]_10 [120]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [120]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [120]),
        .O(\block_w0_reg[24]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[25]_i_10 
       (.I0(\key_mem_reg[11]_11 [121]),
        .I1(\key_mem_reg[10]_10 [121]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [121]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [121]),
        .O(\block_w0_reg[25]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[25]_i_2__0 
       (.I0(\dec_block/op193_in [1]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[25] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[25]_i_3 
       (.I0(\block_w0_reg[25]_i_7_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[25]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[25]_i_9_n_0 ),
        .O(round_key[121]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[25]_i_4 
       (.I0(\block_w0_reg[25]_i_9_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[25]_i_8_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[25]_i_7_n_0 ),
        .I5(dec_new_block[121]),
        .O(\dec_block/op193_in [1]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[25]_i_5 
       (.I0(\block_w2_reg[9]_i_6_n_0 ),
        .I1(\block_w2_reg[14]_i_8_n_0 ),
        .I2(\dec_block/op193_in [0]),
        .I3(\block_w1_reg[16]_i_5_n_0 ),
        .I4(\block_w0_reg[25]_i_6_n_0 ),
        .I5(\block_w0_reg_reg[16] ),
        .O(inv_mixcolumns_return0220_out__63[1]));
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[25]_i_6 
       (.I0(\dec_block/op190_in [1]),
        .I1(\dec_block/op191_in [5]),
        .I2(\dec_block/p_0_in54_in [6]),
        .I3(\dec_block/op190_in [5]),
        .I4(\dec_block/op193_in [5]),
        .O(\block_w0_reg[25]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[25]_i_6__0 
       (.I0(round_key[121]),
        .I1(core_block[121]),
        .O(p_0_out[69]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[25]_i_7 
       (.I0(\block_w0_reg[25]_i_10_n_0 ),
        .I1(\key_mem_reg[14]_14 [121]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [121]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [121]),
        .O(\block_w0_reg[25]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[25]_i_8 
       (.I0(\key_mem_reg[7]_7 [121]),
        .I1(\key_mem_reg[6]_6 [121]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [121]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [121]),
        .O(\block_w0_reg[25]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[25]_i_9 
       (.I0(\key_mem_reg[3]_3 [121]),
        .I1(\key_mem_reg[2]_2 [121]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [121]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [121]),
        .O(\block_w0_reg[25]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[26]_i_3 
       (.I0(\block_w0_reg[26]_i_5__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w0_reg[26]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[26]_i_7_n_0 ),
        .O(round_key[122]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[26]_i_4 
       (.I0(round_key[122]),
        .I1(core_block[122]),
        .O(p_0_out[70]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[26]_i_5 
       (.I0(\block_w3_reg[0]_i_7_n_0 ),
        .I1(\block_w0_reg[26]_i_6_n_0 ),
        .I2(\dec_block/op191_in [7]),
        .I3(\block_w2_reg[14]_i_8_n_0 ),
        .I4(\block_w3_reg[5]_i_11_n_0 ),
        .I5(\dec_block/op193_in [1]),
        .O(inv_mixcolumns_return0220_out__63[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[26]_i_5__0 
       (.I0(\block_w0_reg[26]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [122]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [122]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [122]),
        .O(\block_w0_reg[26]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[26]_i_6 
       (.I0(\dec_block/op190_in [2]),
        .I1(\dec_block/op191_in [1]),
        .O(\block_w0_reg[26]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[26]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [122]),
        .I1(\key_mem_reg[6]_6 [122]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [122]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [122]),
        .O(\block_w0_reg[26]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[26]_i_7 
       (.I0(\key_mem_reg[3]_3 [122]),
        .I1(\key_mem_reg[2]_2 [122]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [122]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [122]),
        .O(\block_w0_reg[26]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[26]_i_8 
       (.I0(\key_mem_reg[11]_11 [122]),
        .I1(\key_mem_reg[10]_10 [122]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [122]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [122]),
        .O(\block_w0_reg[26]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[27]_i_10 
       (.I0(\key_mem_reg[11]_11 [123]),
        .I1(\key_mem_reg[10]_10 [123]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [123]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [123]),
        .O(\block_w0_reg[27]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[27]_i_3 
       (.I0(\block_w0_reg[27]_i_6_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w0_reg[27]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[27]_i_8_n_0 ),
        .O(round_key[123]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[27]_i_4 
       (.I0(\block_w3_reg[6]_i_11_n_0 ),
        .I1(\block_w3_reg[3]_i_9_n_0 ),
        .I2(\dec_block/op193_in [2]),
        .I3(\dec_block/p_0_in54_in [4]),
        .I4(\block_w3_reg[4]_i_10_n_0 ),
        .I5(\block_w3_reg[2]_i_12_n_0 ),
        .O(inv_mixcolumns_return0220_out__63[3]));
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[27]_i_5 
       (.I0(round_key[123]),
        .I1(core_block[123]),
        .O(p_0_out[71]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[27]_i_5__0 
       (.I0(\block_w0_reg[26]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[26]_i_6__0_n_0 ),
        .I3(muxed_round_nr[3]),
        .I4(\block_w0_reg[26]_i_5__0_n_0 ),
        .I5(dec_new_block[122]),
        .O(\dec_block/op193_in [2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[27]_i_6 
       (.I0(\block_w0_reg[27]_i_10_n_0 ),
        .I1(\key_mem_reg[14]_14 [123]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [123]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [123]),
        .O(\block_w0_reg[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[27]_i_7 
       (.I0(\key_mem_reg[7]_7 [123]),
        .I1(\key_mem_reg[6]_6 [123]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [123]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [123]),
        .O(\block_w0_reg[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[27]_i_8 
       (.I0(\key_mem_reg[3]_3 [123]),
        .I1(\key_mem_reg[2]_2 [123]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [123]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [123]),
        .O(\block_w0_reg[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[28]_i_10 
       (.I0(\key_mem_reg[11]_11 [124]),
        .I1(\key_mem_reg[10]_10 [124]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [124]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [124]),
        .O(\block_w0_reg[28]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[28]_i_2__0 
       (.I0(\dec_block/op193_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[28] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[28]_i_3 
       (.I0(\block_w0_reg[28]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[28]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[28]_i_8_n_0 ),
        .O(round_key[124]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[28]_i_4__0 
       (.I0(\block_w0_reg[28]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[28]_i_7_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[28]_i_6__0_n_0 ),
        .I5(dec_new_block[124]),
        .O(\dec_block/op193_in [4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[28]_i_5 
       (.I0(\block_w3_reg[5]_i_10_n_0 ),
        .I1(\block_w3_reg[4]_i_10_n_0 ),
        .I2(\block_w2_reg[9]_i_6_n_0 ),
        .I3(\block_w0_reg[28]_i_6_n_0 ),
        .I4(\block_w3_reg[6]_i_10_n_0 ),
        .I5(\block_w3_reg[3]_i_13_n_0 ),
        .O(inv_mixcolumns_return0220_out__63[4]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[28]_i_5__0 
       (.I0(round_key[124]),
        .I1(core_block[124]),
        .O(p_0_out[72]));
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w0_reg[28]_i_6 
       (.I0(\dec_block/op190_in [7]),
        .I1(round_key[115]),
        .I2(dec_new_block[115]),
        .I3(\dec_block/op190_in [4]),
        .O(\block_w0_reg[28]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[28]_i_6__0 
       (.I0(\block_w0_reg[28]_i_10_n_0 ),
        .I1(\key_mem_reg[14]_14 [124]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [124]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [124]),
        .O(\block_w0_reg[28]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[28]_i_7 
       (.I0(\key_mem_reg[7]_7 [124]),
        .I1(\key_mem_reg[6]_6 [124]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [124]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [124]),
        .O(\block_w0_reg[28]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[28]_i_8 
       (.I0(\key_mem_reg[3]_3 [124]),
        .I1(\key_mem_reg[2]_2 [124]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [124]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [124]),
        .O(\block_w0_reg[28]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[29]_i_2__0 
       (.I0(\dec_block/op193_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[29] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[29]_i_3 
       (.I0(\block_w0_reg[29]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[29]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[29]_i_7__0_n_0 ),
        .O(round_key[125]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[29]_i_4 
       (.I0(\block_w0_reg[29]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[29]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[29]_i_5__0_n_0 ),
        .I5(dec_new_block[125]),
        .O(\dec_block/op193_in [5]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[29]_i_5 
       (.I0(round_key[125]),
        .I1(core_block[125]),
        .O(p_0_out[73]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[29]_i_5__0 
       (.I0(\block_w0_reg[29]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [125]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [125]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [125]),
        .O(\block_w0_reg[29]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[29]_i_6 
       (.I0(\block_w3_reg[5]_i_10_n_0 ),
        .I1(\block_w3_reg[5]_i_11_n_0 ),
        .I2(\block_w0_reg[29]_i_7_n_0 ),
        .I3(\dec_block/op190_in [5]),
        .I4(\block_w3_reg[7]_i_12_n_0 ),
        .I5(\block_w2_reg[13]_i_8_n_0 ),
        .O(inv_mixcolumns_return0220_out__63[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[29]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [125]),
        .I1(\key_mem_reg[6]_6 [125]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [125]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [125]),
        .O(\block_w0_reg[29]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[29]_i_7 
       (.I0(\dec_block/op191_in [4]),
        .I1(\dec_block/op193_in [4]),
        .O(\block_w0_reg[29]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[29]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [125]),
        .I1(\key_mem_reg[2]_2 [125]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [125]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [125]),
        .O(\block_w0_reg[29]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[29]_i_8 
       (.I0(\key_mem_reg[11]_11 [125]),
        .I1(\key_mem_reg[10]_10 [125]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [125]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [125]),
        .O(\block_w0_reg[29]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[2]_i_2__0 
       (.I0(\dec_block/p_0_in54_in [3]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[2] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[2]_i_3 
       (.I0(\block_w0_reg[2]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[2]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[2]_i_7_n_0 ),
        .O(round_key[98]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[2]_i_4 
       (.I0(\block_w0_reg[2]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[2]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[2]_i_5__0_n_0 ),
        .I5(dec_new_block[98]),
        .O(\dec_block/p_0_in54_in [3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[2]_i_5 
       (.I0(round_key[66]),
        .I1(core_block[66]),
        .O(addroundkey_return[31]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[2]_i_5__0 
       (.I0(\block_w0_reg[2]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [98]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [98]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [98]),
        .O(\block_w0_reg[2]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[2]_i_6 
       (.I0(\block_w3_reg[13]_i_10_n_0 ),
        .I1(\dec_block/p_0_in46_in [2]),
        .I2(\dec_block/op161_in [1]),
        .I3(\block_w2_reg[18]_i_7_n_0 ),
        .I4(\block_w3_reg[8]_i_12_n_0 ),
        .I5(\block_w1_reg[27]_i_6_n_0 ),
        .O(inv_mixcolumns_return0166_out__55[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[2]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [98]),
        .I1(\key_mem_reg[6]_6 [98]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [98]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [98]),
        .O(\block_w0_reg[2]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[2]_i_7 
       (.I0(\key_mem_reg[3]_3 [98]),
        .I1(\key_mem_reg[2]_2 [98]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [98]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [98]),
        .O(\block_w0_reg[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[2]_i_8 
       (.I0(\key_mem_reg[11]_11 [98]),
        .I1(\key_mem_reg[10]_10 [98]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [98]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [98]),
        .O(\block_w0_reg[2]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[30]_i_2__0 
       (.I0(\dec_block/op193_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[30] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[30]_i_3 
       (.I0(\block_w0_reg[30]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[30]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[30]_i_7__0_n_0 ),
        .O(round_key[126]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[30]_i_4 
       (.I0(\block_w0_reg[30]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[30]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[30]_i_5__0_n_0 ),
        .I5(dec_new_block[126]),
        .O(\dec_block/op193_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[30]_i_5 
       (.I0(round_key[126]),
        .I1(core_block[126]),
        .O(p_0_out[74]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[30]_i_5__0 
       (.I0(\block_w0_reg[30]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [126]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [126]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [126]),
        .O(\block_w0_reg[30]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[30]_i_6 
       (.I0(\block_w3_reg[4]_i_9_n_0 ),
        .I1(\block_w3_reg[6]_i_11_n_0 ),
        .I2(\block_w3_reg[6]_i_12_n_0 ),
        .I3(\block_w0_reg[30]_i_7_n_0 ),
        .I4(\block_w2_reg[14]_i_8_n_0 ),
        .I5(\dec_block/op190_in [6]),
        .O(inv_mixcolumns_return0220_out__63[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[30]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [126]),
        .I1(\key_mem_reg[6]_6 [126]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [126]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [126]),
        .O(\block_w0_reg[30]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[30]_i_7 
       (.I0(\dec_block/op191_in [5]),
        .I1(\dec_block/op193_in [5]),
        .O(\block_w0_reg[30]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[30]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [126]),
        .I1(\key_mem_reg[2]_2 [126]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [126]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [126]),
        .O(\block_w0_reg[30]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[30]_i_8 
       (.I0(\key_mem_reg[11]_11 [126]),
        .I1(\key_mem_reg[10]_10 [126]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [126]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [126]),
        .O(\block_w0_reg[30]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[31]_i_3__0 
       (.I0(\dec_block/op193_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[31] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[31]_i_4 
       (.I0(\block_w0_reg[31]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[31]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[31]_i_8_n_0 ),
        .O(round_key[127]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[31]_i_5 
       (.I0(round_key[127]),
        .I1(core_block[127]),
        .O(p_0_out[75]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[31]_i_6 
       (.I0(\block_w1_reg[23]_i_7_n_0 ),
        .I1(\dec_block/op193_in [6]),
        .I2(\dec_block/op191_in [6]),
        .I3(\dec_block/op191_in [7]),
        .I4(\block_w3_reg[5]_i_13_n_0 ),
        .O(inv_mixcolumns_return0220_out__63[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[31]_i_6__0 
       (.I0(\block_w0_reg[31]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [127]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [127]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [127]),
        .O(\block_w0_reg[31]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[31]_i_7 
       (.I0(\key_mem_reg[7]_7 [127]),
        .I1(\key_mem_reg[6]_6 [127]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [127]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [127]),
        .O(\block_w0_reg[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[31]_i_8 
       (.I0(\key_mem_reg[3]_3 [127]),
        .I1(\key_mem_reg[2]_2 [127]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [127]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [127]),
        .O(\block_w0_reg[31]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[31]_i_9 
       (.I0(\key_mem_reg[11]_11 [127]),
        .I1(\key_mem_reg[10]_10 [127]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [127]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [127]),
        .O(\block_w0_reg[31]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[3]_i_2__0 
       (.I0(\dec_block/p_0_in54_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[3] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[3]_i_3 
       (.I0(\block_w0_reg[3]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w0_reg[3]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[3]_i_8_n_0 ),
        .O(round_key[99]));
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[3]_i_4__0 
       (.I0(round_key[99]),
        .I1(dec_new_block[99]),
        .O(\dec_block/p_0_in54_in [4]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[3]_i_5 
       (.I0(round_key[99]),
        .I1(core_block[99]),
        .O(p_0_out[48]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[3]_i_5__0 
       (.I0(\block_w3_reg[11]_i_8_n_0 ),
        .I1(\block_w3_reg[12]_i_10_n_0 ),
        .I2(\block_w0_reg[3]_i_6_n_0 ),
        .I3(\block_w0_reg[3]_i_7_n_0 ),
        .I4(\block_w3_reg[10]_i_10_n_0 ),
        .I5(\block_w1_reg[28]_i_7_n_0 ),
        .O(inv_mixcolumns_return0166_out__55[2]));
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[3]_i_6 
       (.I0(\dec_block/op158_in [7]),
        .I1(round_key[83]),
        .I2(dec_new_block[83]),
        .I3(dec_new_block[75]),
        .I4(round_key[75]),
        .O(\block_w0_reg[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[3]_i_6__0 
       (.I0(\block_w0_reg[3]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [99]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [99]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [99]),
        .O(\block_w0_reg[3]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[3]_i_7 
       (.I0(\dec_block/p_0_in46_in [3]),
        .I1(\dec_block/op159_in [5]),
        .I2(\dec_block/p_0_in46_in [6]),
        .I3(\dec_block/op161_in [5]),
        .I4(\dec_block/op158_in [5]),
        .O(\block_w0_reg[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[3]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [99]),
        .I1(\key_mem_reg[6]_6 [99]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [99]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [99]),
        .O(\block_w0_reg[3]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[3]_i_8 
       (.I0(\key_mem_reg[3]_3 [99]),
        .I1(\key_mem_reg[2]_2 [99]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [99]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [99]),
        .O(\block_w0_reg[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[3]_i_9 
       (.I0(\key_mem_reg[11]_11 [99]),
        .I1(\key_mem_reg[10]_10 [99]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [99]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [99]),
        .O(\block_w0_reg[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[4]_i_10 
       (.I0(\key_mem_reg[11]_11 [100]),
        .I1(\key_mem_reg[10]_10 [100]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [100]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [100]),
        .O(\block_w0_reg[4]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[4]_i_2__0 
       (.I0(\dec_block/p_0_in54_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[4] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[4]_i_3 
       (.I0(\block_w0_reg[4]_i_7_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[4]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[4]_i_9_n_0 ),
        .O(round_key[100]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[4]_i_4 
       (.I0(\block_w0_reg[4]_i_9_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[4]_i_8_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[4]_i_7_n_0 ),
        .I5(dec_new_block[100]),
        .O(\dec_block/p_0_in54_in [5]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[4]_i_5__0 
       (.I0(\block_w3_reg[14]_i_10_n_0 ),
        .I1(\dec_block/op159_in [4]),
        .I2(\block_w3_reg[12]_i_9_n_0 ),
        .I3(\block_w3_reg[12]_i_10_n_0 ),
        .I4(\block_w3_reg[13]_i_11_n_0 ),
        .I5(\block_w3_reg[14]_i_12_n_0 ),
        .O(inv_mixcolumns_return0166_out__55[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[4]_i_6 
       (.I0(round_key[100]),
        .I1(core_block[100]),
        .O(p_0_out[49]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[4]_i_7 
       (.I0(\block_w0_reg[4]_i_10_n_0 ),
        .I1(\key_mem_reg[14]_14 [100]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [100]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [100]),
        .O(\block_w0_reg[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[4]_i_8 
       (.I0(\key_mem_reg[7]_7 [100]),
        .I1(\key_mem_reg[6]_6 [100]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [100]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [100]),
        .O(\block_w0_reg[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[4]_i_9 
       (.I0(\key_mem_reg[3]_3 [100]),
        .I1(\key_mem_reg[2]_2 [100]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [100]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [100]),
        .O(\block_w0_reg[4]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[5]_i_2__0 
       (.I0(\dec_block/p_0_in54_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[5] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[5]_i_3 
       (.I0(\block_w0_reg[5]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[5]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[5]_i_7__0_n_0 ),
        .O(round_key[101]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[5]_i_4 
       (.I0(\block_w0_reg[5]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[5]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[5]_i_5__0_n_0 ),
        .I5(dec_new_block[101]),
        .O(\dec_block/p_0_in54_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[5]_i_5 
       (.I0(round_key[69]),
        .I1(core_block[69]),
        .O(addroundkey_return[34]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[5]_i_5__0 
       (.I0(\block_w0_reg[5]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [101]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [101]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [101]),
        .O(\block_w0_reg[5]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[5]_i_6 
       (.I0(\block_w3_reg[13]_i_10_n_0 ),
        .I1(\block_w3_reg[13]_i_11_n_0 ),
        .I2(\block_w0_reg[5]_i_7_n_0 ),
        .I3(\dec_block/op159_in [5]),
        .I4(\block_w3_reg[15]_i_12_n_0 ),
        .I5(\block_w2_reg[21]_i_8_n_0 ),
        .O(inv_mixcolumns_return0166_out__55[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[5]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [101]),
        .I1(\key_mem_reg[6]_6 [101]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [101]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [101]),
        .O(\block_w0_reg[5]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[5]_i_7 
       (.I0(\dec_block/p_0_in46_in [5]),
        .I1(\dec_block/op161_in [4]),
        .O(\block_w0_reg[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[5]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [101]),
        .I1(\key_mem_reg[2]_2 [101]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [101]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [101]),
        .O(\block_w0_reg[5]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[5]_i_8 
       (.I0(\key_mem_reg[11]_11 [101]),
        .I1(\key_mem_reg[10]_10 [101]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [101]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [101]),
        .O(\block_w0_reg[5]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[6]_i_2__0 
       (.I0(\dec_block/p_0_in54_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[6] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[6]_i_3 
       (.I0(\block_w0_reg[6]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[6]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[6]_i_7__0_n_0 ),
        .O(round_key[102]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[6]_i_4 
       (.I0(\block_w0_reg[6]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[6]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[6]_i_5__0_n_0 ),
        .I5(dec_new_block[102]),
        .O(\dec_block/p_0_in54_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[6]_i_5 
       (.I0(round_key[70]),
        .I1(core_block[70]),
        .O(addroundkey_return[35]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[6]_i_5__0 
       (.I0(\block_w0_reg[6]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [102]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [102]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [102]),
        .O(\block_w0_reg[6]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[6]_i_6 
       (.I0(\block_w3_reg[12]_i_12_n_0 ),
        .I1(\block_w3_reg[14]_i_11_n_0 ),
        .I2(\block_w3_reg[14]_i_12_n_0 ),
        .I3(\block_w0_reg[6]_i_7_n_0 ),
        .I4(\block_w3_reg[11]_i_9_n_0 ),
        .I5(\dec_block/op159_in [6]),
        .O(inv_mixcolumns_return0166_out__55[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[6]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [102]),
        .I1(\key_mem_reg[6]_6 [102]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [102]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [102]),
        .O(\block_w0_reg[6]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[6]_i_7 
       (.I0(\dec_block/op161_in [5]),
        .I1(\dec_block/p_0_in46_in [6]),
        .O(\block_w0_reg[6]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[6]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [102]),
        .I1(\key_mem_reg[2]_2 [102]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [102]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [102]),
        .O(\block_w0_reg[6]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[6]_i_8 
       (.I0(\key_mem_reg[11]_11 [102]),
        .I1(\key_mem_reg[10]_10 [102]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [102]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [102]),
        .O(\block_w0_reg[6]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[7]_i_2__0 
       (.I0(\block_w0_reg[7]_i_4_n_0 ),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[7] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[7]_i_3 
       (.I0(\block_w0_reg[7]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[7]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[7]_i_7_n_0 ),
        .O(round_key[103]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[7]_i_4 
       (.I0(\block_w0_reg[7]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[7]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[7]_i_5__0_n_0 ),
        .I5(dec_new_block[103]),
        .O(\block_w0_reg[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[7]_i_5 
       (.I0(round_key[71]),
        .I1(core_block[71]),
        .O(addroundkey_return[36]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[7]_i_5__0 
       (.I0(\block_w0_reg[7]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [103]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [103]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [103]),
        .O(\block_w0_reg[7]_i_5__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[7]_i_6 
       (.I0(\block_w3_reg[15]_i_11_n_0 ),
        .I1(\dec_block/op161_in [6]),
        .I2(\dec_block/p_0_in46_in [7]),
        .I3(\dec_block/op158_in [7]),
        .I4(\block_w3_reg[13]_i_13_n_0 ),
        .O(inv_mixcolumns_return0166_out__55[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[7]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [103]),
        .I1(\key_mem_reg[6]_6 [103]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [103]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [103]),
        .O(\block_w0_reg[7]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[7]_i_7 
       (.I0(\key_mem_reg[3]_3 [103]),
        .I1(\key_mem_reg[2]_2 [103]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [103]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [103]),
        .O(\block_w0_reg[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[7]_i_8 
       (.I0(\key_mem_reg[11]_11 [103]),
        .I1(\key_mem_reg[10]_10 [103]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [103]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [103]),
        .O(\block_w0_reg[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[8]_i_2__0 
       (.I0(\dec_block/op190_in [0]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[8] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[8]_i_3 
       (.I0(\block_w0_reg[8]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[8]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[8]_i_7_n_0 ),
        .O(round_key[104]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[8]_i_4 
       (.I0(round_key[40]),
        .I1(core_block[40]),
        .O(addroundkey_return[22]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[8]_i_5 
       (.I0(\block_w2_reg[24]_i_7_n_0 ),
        .I1(\dec_block/op129_in [0]),
        .I2(\block_w3_reg[17]_i_9_n_0 ),
        .I3(\block_w2_reg[24]_i_9_n_0 ),
        .I4(\block_w3_reg[22]_i_14_n_0 ),
        .O(inv_mixcolumns_return0142_out__55[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[8]_i_5__0 
       (.I0(\block_w0_reg[8]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [104]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [104]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [104]),
        .O(\block_w0_reg[8]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[8]_i_6 
       (.I0(\key_mem_reg[7]_7 [104]),
        .I1(\key_mem_reg[6]_6 [104]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [104]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [104]),
        .O(\block_w0_reg[8]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[8]_i_7 
       (.I0(\key_mem_reg[3]_3 [104]),
        .I1(\key_mem_reg[2]_2 [104]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [104]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [104]),
        .O(\block_w0_reg[8]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[8]_i_8 
       (.I0(\key_mem_reg[11]_11 [104]),
        .I1(\key_mem_reg[10]_10 [104]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [104]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [104]),
        .O(\block_w0_reg[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[9]_i_10 
       (.I0(\key_mem_reg[11]_11 [105]),
        .I1(\key_mem_reg[10]_10 [105]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [105]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [105]),
        .O(\block_w0_reg[9]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w0_reg[9]_i_2__0 
       (.I0(\dec_block/op190_in [1]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w0_reg_reg[9] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w0_reg[9]_i_3 
       (.I0(\block_w0_reg[9]_i_7__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w0_reg[9]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w0_reg[9]_i_9_n_0 ),
        .O(round_key[105]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w0_reg[9]_i_4 
       (.I0(\block_w0_reg[9]_i_9_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[9]_i_8_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[9]_i_7__0_n_0 ),
        .I5(dec_new_block[105]),
        .O(\dec_block/op190_in [1]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w0_reg[9]_i_5__0 
       (.I0(\block_w3_reg[20]_i_11_n_0 ),
        .I1(\block_w2_reg[30]_i_8_n_0 ),
        .I2(\dec_block/op126_in [0]),
        .I3(\block_w0_reg[9]_i_6__0_n_0 ),
        .I4(\block_w0_reg[9]_i_7_n_0 ),
        .I5(\block_w2_reg_reg[0] ),
        .O(inv_mixcolumns_return0142_out__55[1]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[9]_i_6 
       (.I0(round_key[105]),
        .I1(core_block[105]),
        .O(p_0_out[54]));
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w0_reg[9]_i_6__0 
       (.I0(\block_w2_reg[7]_i_4_n_0 ),
        .I1(\dec_block/op129_in [7]),
        .O(\block_w0_reg[9]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w0_reg[9]_i_7 
       (.I0(\dec_block/op129_in [1]),
        .I1(\dec_block/op129_in [5]),
        .I2(\dec_block/op126_in [5]),
        .I3(\dec_block/p_0_in38_in [6]),
        .I4(\dec_block/op127_in [5]),
        .O(\block_w0_reg[9]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[9]_i_7__0 
       (.I0(\block_w0_reg[9]_i_10_n_0 ),
        .I1(\key_mem_reg[14]_14 [105]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [105]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [105]),
        .O(\block_w0_reg[9]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[9]_i_8 
       (.I0(\key_mem_reg[7]_7 [105]),
        .I1(\key_mem_reg[6]_6 [105]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[5]_5 [105]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[4]_4 [105]),
        .O(\block_w0_reg[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w0_reg[9]_i_9 
       (.I0(\key_mem_reg[3]_3 [105]),
        .I1(\key_mem_reg[2]_2 [105]),
        .I2(muxed_round_nr[1]),
        .I3(\key_mem_reg[1]_1 [105]),
        .I4(muxed_round_nr[0]),
        .I5(\key_mem_reg[0]_0 [105]),
        .O(\block_w0_reg[9]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'h60)) 
    \block_w1_reg[0]_i_2__0 
       (.I0(round_key[32]),
        .I1(core_block[32]),
        .I2(\block_w0_reg_reg[0]_1 ),
        .O(\block_reg_reg[2][0] ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \block_w1_reg[0]_i_3 
       (.I0(\dec_block/op129_in [7]),
        .I1(\block_w2_reg_reg[16] ),
        .I2(\block_w3_reg[16]_i_7_n_0 ),
        .I3(\block_w1_reg[0]_i_5_n_0 ),
        .I4(\block_w0_reg_reg[0]_1 ),
        .I5(\block_w0_reg_reg[16]_0 [0]),
        .O(\block_w2_reg_reg[31]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[0]_i_3__0 
       (.I0(\block_w1_reg[0]_i_5__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w1_reg[0]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[0]_i_7_n_0 ),
        .O(round_key[64]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[0]_i_4 
       (.I0(\block_w1_reg[0]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[0]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[0]_i_5__0_n_0 ),
        .I5(dec_new_block[64]),
        .O(\block_w1_reg_reg[0] ));
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \block_w1_reg[0]_i_5 
       (.I0(\dec_block/op126_in [0]),
        .I1(\dec_block/op129_in [0]),
        .I2(\block_w2_reg[7]_i_4_n_0 ),
        .O(\block_w1_reg[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[0]_i_5__0 
       (.I0(\block_w1_reg[0]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [64]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [64]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [64]),
        .O(\block_w1_reg[0]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[0]_i_6 
       (.I0(\key_mem_reg[7]_7 [64]),
        .I1(\key_mem_reg[6]_6 [64]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [64]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [64]),
        .O(\block_w1_reg[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[0]_i_7 
       (.I0(\key_mem_reg[3]_3 [64]),
        .I1(\key_mem_reg[2]_2 [64]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [64]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [64]),
        .O(\block_w1_reg[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[0]_i_8 
       (.I0(\key_mem_reg[11]_11 [64]),
        .I1(\key_mem_reg[10]_10 [64]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [64]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [64]),
        .O(\block_w1_reg[0]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[10]_i_2__0 
       (.I0(\dec_block/op158_in [2]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[10] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[10]_i_3 
       (.I0(\block_w1_reg[10]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[10]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[10]_i_7_n_0 ),
        .O(round_key[74]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[10]_i_4 
       (.I0(\block_w1_reg[10]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[10]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[10]_i_5__0_n_0 ),
        .I5(dec_new_block[74]),
        .O(\dec_block/op158_in [2]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[10]_i_5 
       (.I0(round_key[10]),
        .I1(core_block[10]),
        .O(addroundkey_return[9]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[10]_i_5__0 
       (.I0(\block_w1_reg[10]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [74]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [74]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [74]),
        .O(\block_w1_reg[10]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[10]_i_6 
       (.I0(\block_w3_reg[29]_i_11_n_0 ),
        .I1(\block_w2_reg[0]_i_6_n_0 ),
        .I2(\dec_block/p_0_in31_in [2]),
        .I3(\dec_block/op96_in [7]),
        .I4(\block_w2_reg[3]_i_8_n_0 ),
        .I5(\dec_block/op95_in [1]),
        .O(inv_mixcolumns_return0110_out__47[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[10]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [74]),
        .I1(\key_mem_reg[6]_6 [74]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [74]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [74]),
        .O(\block_w1_reg[10]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[10]_i_7 
       (.I0(\key_mem_reg[3]_3 [74]),
        .I1(\key_mem_reg[2]_2 [74]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [74]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [74]),
        .O(\block_w1_reg[10]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[10]_i_8 
       (.I0(\key_mem_reg[11]_11 [74]),
        .I1(\key_mem_reg[10]_10 [74]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [74]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [74]),
        .O(\block_w1_reg[10]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[11]_i_3 
       (.I0(\block_w1_reg[11]_i_6_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w1_reg[11]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[11]_i_8_n_0 ),
        .O(round_key[75]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[11]_i_4 
       (.I0(\block_w3_reg[27]_i_8_n_0 ),
        .I1(\block_w3_reg[28]_i_9_n_0 ),
        .I2(\block_w3_reg[24]_i_13_n_0 ),
        .I3(\block_w1_reg[11]_i_5__0_n_0 ),
        .I4(\block_w3_reg[30]_i_12_n_0 ),
        .I5(\dec_block/op96_in [3]),
        .O(inv_mixcolumns_return0110_out__47[2]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[11]_i_5 
       (.I0(round_key[75]),
        .I1(core_block[75]),
        .O(p_0_out[33]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[11]_i_5__0 
       (.I0(\dec_block/op95_in [2]),
        .I1(\dec_block/p_0_in31_in [3]),
        .O(\block_w1_reg[11]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[11]_i_6 
       (.I0(\block_w1_reg[11]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [75]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [75]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [75]),
        .O(\block_w1_reg[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[11]_i_7 
       (.I0(\key_mem_reg[7]_7 [75]),
        .I1(\key_mem_reg[6]_6 [75]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [75]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [75]),
        .O(\block_w1_reg[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[11]_i_8 
       (.I0(\key_mem_reg[3]_3 [75]),
        .I1(\key_mem_reg[2]_2 [75]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [75]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [75]),
        .O(\block_w1_reg[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[11]_i_9 
       (.I0(\key_mem_reg[11]_11 [75]),
        .I1(\key_mem_reg[10]_10 [75]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [75]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [75]),
        .O(\block_w1_reg[11]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[12]_i_2__0 
       (.I0(\dec_block/op158_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[12] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[12]_i_3 
       (.I0(\block_w1_reg[12]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[12]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[12]_i_8_n_0 ),
        .O(round_key[76]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[12]_i_4__0 
       (.I0(\block_w1_reg[12]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[12]_i_7__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[12]_i_6__0_n_0 ),
        .I5(dec_new_block[76]),
        .O(\dec_block/op158_in [4]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[12]_i_5 
       (.I0(round_key[76]),
        .I1(core_block[76]),
        .O(p_0_out[34]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[12]_i_5__0 
       (.I0(\block_w3_reg[29]_i_10_n_0 ),
        .I1(\block_w3_reg[28]_i_9_n_0 ),
        .I2(\block_w1_reg[9]_i_6__0_n_0 ),
        .I3(\block_w1_reg[12]_i_6_n_0 ),
        .I4(\block_w3_reg[28]_i_11_n_0 ),
        .I5(\block_w1_reg[12]_i_7_n_0 ),
        .O(inv_mixcolumns_return0110_out__47[3]));
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w1_reg[12]_i_6 
       (.I0(\block_w3_reg[7]_i_4_n_0 ),
        .I1(round_key[11]),
        .I2(dec_new_block[11]),
        .I3(\dec_block/op98_in [4]),
        .O(\block_w1_reg[12]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[12]_i_6__0 
       (.I0(\block_w1_reg[12]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [76]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [76]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [76]),
        .O(\block_w1_reg[12]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \block_w1_reg[12]_i_7 
       (.I0(dec_new_block[3]),
        .I1(round_key[3]),
        .I2(\dec_block/op98_in [7]),
        .O(\block_w1_reg[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[12]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [76]),
        .I1(\key_mem_reg[6]_6 [76]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [76]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [76]),
        .O(\block_w1_reg[12]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[12]_i_8 
       (.I0(\key_mem_reg[3]_3 [76]),
        .I1(\key_mem_reg[2]_2 [76]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [76]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [76]),
        .O(\block_w1_reg[12]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[12]_i_9 
       (.I0(\key_mem_reg[11]_11 [76]),
        .I1(\key_mem_reg[10]_10 [76]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [76]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [76]),
        .O(\block_w1_reg[12]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[13]_i_2__0 
       (.I0(\dec_block/op158_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[13] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[13]_i_3 
       (.I0(\block_w1_reg[13]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[13]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[13]_i_7__0_n_0 ),
        .O(round_key[77]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[13]_i_4 
       (.I0(\block_w1_reg[13]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[13]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[13]_i_5__0_n_0 ),
        .I5(dec_new_block[77]),
        .O(\dec_block/op158_in [5]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[13]_i_5 
       (.I0(round_key[13]),
        .I1(core_block[13]),
        .O(addroundkey_return[12]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[13]_i_5__0 
       (.I0(\block_w1_reg[13]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [77]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [77]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [77]),
        .O(\block_w1_reg[13]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[13]_i_6 
       (.I0(\block_w3_reg[29]_i_10_n_0 ),
        .I1(\block_w3_reg[29]_i_11_n_0 ),
        .I2(\block_w1_reg[13]_i_7_n_0 ),
        .I3(\dec_block/op98_in [5]),
        .I4(\block_w3_reg[29]_i_13_n_0 ),
        .I5(\block_w3_reg[29]_i_14_n_0 ),
        .O(inv_mixcolumns_return0110_out__47[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[13]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [77]),
        .I1(\key_mem_reg[6]_6 [77]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [77]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [77]),
        .O(\block_w1_reg[13]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[13]_i_7 
       (.I0(\dec_block/op95_in [4]),
        .I1(\dec_block/p_0_in31_in [5]),
        .O(\block_w1_reg[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[13]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [77]),
        .I1(\key_mem_reg[2]_2 [77]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [77]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [77]),
        .O(\block_w1_reg[13]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[13]_i_8 
       (.I0(\key_mem_reg[11]_11 [77]),
        .I1(\key_mem_reg[10]_10 [77]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [77]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [77]),
        .O(\block_w1_reg[13]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[14]_i_2__0 
       (.I0(\dec_block/op158_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[14] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[14]_i_3 
       (.I0(\block_w1_reg[14]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[14]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[14]_i_7__0_n_0 ),
        .O(round_key[78]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[14]_i_4 
       (.I0(\block_w1_reg[14]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[14]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[14]_i_5__0_n_0 ),
        .I5(dec_new_block[78]),
        .O(\dec_block/op158_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[14]_i_5 
       (.I0(round_key[14]),
        .I1(core_block[14]),
        .O(addroundkey_return[13]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[14]_i_5__0 
       (.I0(\block_w1_reg[14]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [78]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [78]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [78]),
        .O(\block_w1_reg[14]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[14]_i_6 
       (.I0(\block_w3_reg[30]_i_10_n_0 ),
        .I1(\block_w3_reg[30]_i_11_n_0 ),
        .I2(\block_w3_reg[30]_i_12_n_0 ),
        .I3(\block_w1_reg[14]_i_7_n_0 ),
        .I4(\block_w3_reg[30]_i_14_n_0 ),
        .I5(\dec_block/op98_in [6]),
        .O(inv_mixcolumns_return0110_out__47[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[14]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [78]),
        .I1(\key_mem_reg[6]_6 [78]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [78]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [78]),
        .O(\block_w1_reg[14]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[14]_i_7 
       (.I0(\dec_block/op95_in [5]),
        .I1(\dec_block/p_0_in31_in [6]),
        .O(\block_w1_reg[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[14]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [78]),
        .I1(\key_mem_reg[2]_2 [78]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [78]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [78]),
        .O(\block_w1_reg[14]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[14]_i_8 
       (.I0(\key_mem_reg[11]_11 [78]),
        .I1(\key_mem_reg[10]_10 [78]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [78]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [78]),
        .O(\block_w1_reg[14]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[15]_i_2__0 
       (.I0(\dec_block/op158_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[15] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[15]_i_3 
       (.I0(\block_w1_reg[15]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[15]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[15]_i_7_n_0 ),
        .O(round_key[79]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[15]_i_4 
       (.I0(\block_w1_reg[15]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[15]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[15]_i_5__0_n_0 ),
        .I5(dec_new_block[79]),
        .O(\dec_block/op158_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[15]_i_5 
       (.I0(round_key[15]),
        .I1(core_block[15]),
        .O(addroundkey_return[14]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[15]_i_5__0 
       (.I0(\block_w1_reg[15]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [79]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [79]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [79]),
        .O(\block_w1_reg[15]_i_5__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[15]_i_6 
       (.I0(\block_w2_reg[7]_i_7_n_0 ),
        .I1(\dec_block/op95_in [6]),
        .I2(\dec_block/p_0_in31_in [7]),
        .I3(\block_w3_reg[7]_i_4_n_0 ),
        .I4(\block_w3_reg[31]_i_14_n_0 ),
        .O(inv_mixcolumns_return0110_out__47[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[15]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [79]),
        .I1(\key_mem_reg[6]_6 [79]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [79]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [79]),
        .O(\block_w1_reg[15]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[15]_i_7 
       (.I0(\key_mem_reg[3]_3 [79]),
        .I1(\key_mem_reg[2]_2 [79]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [79]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [79]),
        .O(\block_w1_reg[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[15]_i_8 
       (.I0(\key_mem_reg[11]_11 [79]),
        .I1(\key_mem_reg[10]_10 [79]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [79]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [79]),
        .O(\block_w1_reg[15]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT3 #(
    .INIT(8'h60)) 
    \block_w1_reg[16]_i_2__0 
       (.I0(round_key[112]),
        .I1(core_block[112]),
        .I2(\block_w0_reg_reg[0]_1 ),
        .O(\block_reg_reg[0][16] ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \block_w1_reg[16]_i_3 
       (.I0(\block_w1_reg[16]_i_5_n_0 ),
        .I1(\block_w3_reg[0]_i_6_n_0 ),
        .I2(\block_w0_reg_reg[0] ),
        .I3(\block_w1_reg[16]_i_6_n_0 ),
        .I4(\block_w0_reg_reg[0]_1 ),
        .I5(\block_w0_reg_reg[16]_0 [2]),
        .O(\block_w0_reg_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[16]_i_3__0 
       (.I0(\block_w1_reg[16]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[16]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[16]_i_7_n_0 ),
        .O(round_key[80]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[16]_i_4 
       (.I0(\block_w1_reg[16]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[16]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[16]_i_5__0_n_0 ),
        .I5(dec_new_block[80]),
        .O(\block_w1_reg_reg[16] ));
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[16]_i_5 
       (.I0(\dec_block/op190_in [7]),
        .I1(\dec_block/op191_in [7]),
        .O(\block_w1_reg[16]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[16]_i_5__0 
       (.I0(\block_w1_reg[16]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [80]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [80]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [80]),
        .O(\block_w1_reg[16]_i_5__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[16]_i_6 
       (.I0(\dec_block/op190_in [0]),
        .I1(\dec_block/op193_in [0]),
        .O(\block_w1_reg[16]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[16]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [80]),
        .I1(\key_mem_reg[6]_6 [80]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [80]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [80]),
        .O(\block_w1_reg[16]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[16]_i_7 
       (.I0(\key_mem_reg[3]_3 [80]),
        .I1(\key_mem_reg[2]_2 [80]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [80]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [80]),
        .O(\block_w1_reg[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[16]_i_8 
       (.I0(\key_mem_reg[11]_11 [80]),
        .I1(\key_mem_reg[10]_10 [80]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [80]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [80]),
        .O(\block_w1_reg[16]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[17]_i_2__0 
       (.I0(\dec_block/op159_in [1]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[17] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[17]_i_3 
       (.I0(\block_w1_reg[17]_i_6_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[17]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[17]_i_8_n_0 ),
        .O(round_key[81]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[17]_i_4__0 
       (.I0(\block_w1_reg[17]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[17]_i_7_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[17]_i_6_n_0 ),
        .I5(dec_new_block[81]),
        .O(\dec_block/op159_in [1]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[17]_i_5 
       (.I0(\block_w0_reg_reg[16] ),
        .I1(\dec_block/p_0_in54_in [2]),
        .I2(\block_w3_reg[4]_i_10_n_0 ),
        .I3(\block_w3_reg[6]_i_14_n_0 ),
        .I4(\dec_block/op190_in [0]),
        .I5(\block_w2_reg[8]_i_8_n_0 ),
        .O(inv_mixcolumns_return0213_out__55[0]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[17]_i_5__0 
       (.I0(round_key[81]),
        .I1(core_block[81]),
        .O(addroundkey_return[37]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[17]_i_6 
       (.I0(\block_w1_reg[17]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [81]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [81]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [81]),
        .O(\block_w1_reg[17]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[17]_i_7 
       (.I0(\key_mem_reg[7]_7 [81]),
        .I1(\key_mem_reg[6]_6 [81]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [81]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [81]),
        .O(\block_w1_reg[17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[17]_i_8 
       (.I0(\key_mem_reg[3]_3 [81]),
        .I1(\key_mem_reg[2]_2 [81]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [81]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [81]),
        .O(\block_w1_reg[17]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[17]_i_9 
       (.I0(\key_mem_reg[11]_11 [81]),
        .I1(\key_mem_reg[10]_10 [81]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [81]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [81]),
        .O(\block_w1_reg[17]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[18]_i_3 
       (.I0(\block_w1_reg[18]_i_5__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w1_reg[18]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[18]_i_7_n_0 ),
        .O(round_key[82]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[18]_i_4 
       (.I0(round_key[114]),
        .I1(core_block[114]),
        .O(p_0_out[62]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[18]_i_5 
       (.I0(\block_w1_reg[18]_i_6_n_0 ),
        .I1(\dec_block/p_0_in54_in [3]),
        .I2(\dec_block/op191_in [1]),
        .I3(\block_w3_reg[2]_i_10_n_0 ),
        .I4(\block_w3_reg[5]_i_10_n_0 ),
        .I5(\dec_block/op190_in [1]),
        .O(inv_mixcolumns_return0213_out__55[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[18]_i_5__0 
       (.I0(\block_w1_reg[18]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [82]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [82]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [82]),
        .O(\block_w1_reg[18]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w1_reg[18]_i_6 
       (.I0(\block_w0_reg_reg[0] ),
        .I1(\block_w0_reg_reg[16] ),
        .I2(\dec_block/op193_in [6]),
        .I3(\dec_block/op190_in [6]),
        .O(\block_w1_reg[18]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[18]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [82]),
        .I1(\key_mem_reg[6]_6 [82]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [82]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [82]),
        .O(\block_w1_reg[18]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[18]_i_7 
       (.I0(\key_mem_reg[3]_3 [82]),
        .I1(\key_mem_reg[2]_2 [82]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [82]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [82]),
        .O(\block_w1_reg[18]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[18]_i_8 
       (.I0(\key_mem_reg[11]_11 [82]),
        .I1(\key_mem_reg[10]_10 [82]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [82]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [82]),
        .O(\block_w1_reg[18]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[19]_i_2__0 
       (.I0(\dec_block/op159_in [3]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[19] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[19]_i_3 
       (.I0(\block_w1_reg[19]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w1_reg[19]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[19]_i_8__0_n_0 ),
        .O(round_key[83]));
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[19]_i_4__0 
       (.I0(round_key[83]),
        .I1(dec_new_block[83]),
        .O(\dec_block/op159_in [3]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[19]_i_5 
       (.I0(\block_w3_reg[0]_i_6_n_0 ),
        .I1(\block_w3_reg[3]_i_9_n_0 ),
        .I2(\block_w1_reg[19]_i_6_n_0 ),
        .I3(\block_w2_reg[9]_i_6_n_0 ),
        .I4(\block_w2_reg[12]_i_7_n_0 ),
        .O(inv_mixcolumns_return0213_out__55[2]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[19]_i_5__0 
       (.I0(round_key[83]),
        .I1(core_block[83]),
        .O(addroundkey_return[39]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[19]_i_6 
       (.I0(\dec_block/op191_in [2]),
        .I1(dec_new_block[107]),
        .I2(round_key[107]),
        .I3(\block_w0_reg[7]_i_4_n_0 ),
        .I4(\dec_block/op190_in [2]),
        .I5(\dec_block/op193_in [3]),
        .O(\block_w1_reg[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[19]_i_6__0 
       (.I0(\block_w1_reg[19]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [83]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [83]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [83]),
        .O(\block_w1_reg[19]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[19]_i_7 
       (.I0(\block_w0_reg[18]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[18]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[18]_i_5__0_n_0 ),
        .I5(dec_new_block[114]),
        .O(\dec_block/op191_in [2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[19]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [83]),
        .I1(\key_mem_reg[6]_6 [83]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [83]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [83]),
        .O(\block_w1_reg[19]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[19]_i_8 
       (.I0(\block_w0_reg[27]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[27]_i_7_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[27]_i_6_n_0 ),
        .I5(dec_new_block[123]),
        .O(\dec_block/op193_in [3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[19]_i_8__0 
       (.I0(\key_mem_reg[3]_3 [83]),
        .I1(\key_mem_reg[2]_2 [83]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [83]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [83]),
        .O(\block_w1_reg[19]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[19]_i_9 
       (.I0(\key_mem_reg[11]_11 [83]),
        .I1(\key_mem_reg[10]_10 [83]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [83]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [83]),
        .O(\block_w1_reg[19]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[1]_i_2__0 
       (.I0(\dec_block/p_0_in46_in [2]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[1] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[1]_i_3 
       (.I0(\block_w1_reg[1]_i_6_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[1]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[1]_i_8_n_0 ),
        .O(round_key[65]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[1]_i_4__0 
       (.I0(\block_w1_reg[1]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[1]_i_7_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[1]_i_6_n_0 ),
        .I5(dec_new_block[65]),
        .O(\dec_block/p_0_in46_in [2]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[1]_i_5 
       (.I0(round_key[65]),
        .I1(core_block[65]),
        .O(addroundkey_return[30]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[1]_i_5__0 
       (.I0(\block_w2_reg_reg[0] ),
        .I1(\dec_block/op127_in [1]),
        .I2(\block_w3_reg[20]_i_10_n_0 ),
        .I3(\block_w3_reg[22]_i_14_n_0 ),
        .I4(\dec_block/op129_in [0]),
        .I5(\block_w2_reg[24]_i_8_n_0 ),
        .O(inv_mixcolumns_return0134_out__63[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[1]_i_6 
       (.I0(\block_w1_reg[1]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [65]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [65]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [65]),
        .O(\block_w1_reg[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[1]_i_7 
       (.I0(\key_mem_reg[7]_7 [65]),
        .I1(\key_mem_reg[6]_6 [65]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [65]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [65]),
        .O(\block_w1_reg[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[1]_i_8 
       (.I0(\key_mem_reg[3]_3 [65]),
        .I1(\key_mem_reg[2]_2 [65]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [65]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [65]),
        .O(\block_w1_reg[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[1]_i_9 
       (.I0(\key_mem_reg[11]_11 [65]),
        .I1(\key_mem_reg[10]_10 [65]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [65]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [65]),
        .O(\block_w1_reg[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[20]_i_10 
       (.I0(\key_mem_reg[11]_11 [84]),
        .I1(\key_mem_reg[10]_10 [84]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [84]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [84]),
        .O(\block_w1_reg[20]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[20]_i_2__0 
       (.I0(\dec_block/op159_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[20] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[20]_i_3 
       (.I0(\block_w1_reg[20]_i_7_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[20]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[20]_i_9_n_0 ),
        .O(round_key[84]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[20]_i_4 
       (.I0(\block_w1_reg[20]_i_9_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[20]_i_8_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[20]_i_7_n_0 ),
        .I5(dec_new_block[84]),
        .O(\dec_block/op159_in [4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[20]_i_5 
       (.I0(\block_w3_reg[4]_i_9_n_0 ),
        .I1(\dec_block/p_0_in54_in [5]),
        .I2(\block_w3_reg[4]_i_10_n_0 ),
        .I3(\block_w2_reg[9]_i_6_n_0 ),
        .I4(\block_w3_reg[5]_i_11_n_0 ),
        .I5(\block_w3_reg[6]_i_11_n_0 ),
        .O(inv_mixcolumns_return0213_out__55[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[20]_i_6 
       (.I0(round_key[84]),
        .I1(core_block[84]),
        .O(addroundkey_return[40]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[20]_i_7 
       (.I0(\block_w1_reg[20]_i_10_n_0 ),
        .I1(\key_mem_reg[14]_14 [84]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [84]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [84]),
        .O(\block_w1_reg[20]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[20]_i_8 
       (.I0(\key_mem_reg[7]_7 [84]),
        .I1(\key_mem_reg[6]_6 [84]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [84]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [84]),
        .O(\block_w1_reg[20]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[20]_i_9 
       (.I0(\key_mem_reg[3]_3 [84]),
        .I1(\key_mem_reg[2]_2 [84]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [84]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [84]),
        .O(\block_w1_reg[20]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[21]_i_2__0 
       (.I0(\dec_block/op159_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[21] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[21]_i_3 
       (.I0(\block_w1_reg[21]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[21]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[21]_i_7__0_n_0 ),
        .O(round_key[85]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[21]_i_4 
       (.I0(\block_w1_reg[21]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[21]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[21]_i_5__0_n_0 ),
        .I5(dec_new_block[85]),
        .O(\dec_block/op159_in [5]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[21]_i_5 
       (.I0(round_key[117]),
        .I1(core_block[117]),
        .O(p_0_out[65]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[21]_i_5__0 
       (.I0(\block_w1_reg[21]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [85]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [85]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [85]),
        .O(\block_w1_reg[21]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[21]_i_6 
       (.I0(\block_w3_reg[5]_i_10_n_0 ),
        .I1(\block_w3_reg[5]_i_11_n_0 ),
        .I2(\block_w1_reg[21]_i_7_n_0 ),
        .I3(\dec_block/p_0_in54_in [6]),
        .I4(\block_w3_reg[5]_i_13_n_0 ),
        .I5(\block_w3_reg[5]_i_14_n_0 ),
        .O(inv_mixcolumns_return0213_out__55[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[21]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [85]),
        .I1(\key_mem_reg[6]_6 [85]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [85]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [85]),
        .O(\block_w1_reg[21]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[21]_i_7 
       (.I0(\dec_block/op191_in [4]),
        .I1(\dec_block/op190_in [4]),
        .O(\block_w1_reg[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[21]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [85]),
        .I1(\key_mem_reg[2]_2 [85]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [85]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [85]),
        .O(\block_w1_reg[21]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[21]_i_8 
       (.I0(\key_mem_reg[11]_11 [85]),
        .I1(\key_mem_reg[10]_10 [85]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [85]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [85]),
        .O(\block_w1_reg[21]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[22]_i_2__0 
       (.I0(\dec_block/op159_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[22] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[22]_i_3 
       (.I0(\block_w1_reg[22]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[22]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[22]_i_7__0_n_0 ),
        .O(round_key[86]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[22]_i_4 
       (.I0(\block_w1_reg[22]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[22]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[22]_i_5__0_n_0 ),
        .I5(dec_new_block[86]),
        .O(\dec_block/op159_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[22]_i_5 
       (.I0(round_key[118]),
        .I1(core_block[118]),
        .O(p_0_out[66]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[22]_i_5__0 
       (.I0(\block_w1_reg[22]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [86]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [86]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [86]),
        .O(\block_w1_reg[22]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[22]_i_6 
       (.I0(\block_w3_reg[6]_i_10_n_0 ),
        .I1(\block_w3_reg[6]_i_11_n_0 ),
        .I2(\block_w3_reg[6]_i_12_n_0 ),
        .I3(\block_w1_reg[22]_i_7_n_0 ),
        .I4(\block_w3_reg[6]_i_14_n_0 ),
        .I5(\dec_block/p_0_in54_in [7]),
        .O(inv_mixcolumns_return0213_out__55[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[22]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [86]),
        .I1(\key_mem_reg[6]_6 [86]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [86]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [86]),
        .O(\block_w1_reg[22]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[22]_i_7 
       (.I0(\dec_block/op190_in [5]),
        .I1(\dec_block/op191_in [5]),
        .O(\block_w1_reg[22]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[22]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [86]),
        .I1(\key_mem_reg[2]_2 [86]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [86]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [86]),
        .O(\block_w1_reg[22]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[22]_i_8 
       (.I0(\key_mem_reg[11]_11 [86]),
        .I1(\key_mem_reg[10]_10 [86]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [86]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [86]),
        .O(\block_w1_reg[22]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[23]_i_2__0 
       (.I0(\dec_block/op159_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[23] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[23]_i_3 
       (.I0(\block_w1_reg[23]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[23]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[23]_i_7__0_n_0 ),
        .O(round_key[87]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[23]_i_4 
       (.I0(\block_w1_reg[23]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[23]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[23]_i_5__0_n_0 ),
        .I5(dec_new_block[87]),
        .O(\dec_block/op159_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[23]_i_5 
       (.I0(round_key[119]),
        .I1(core_block[119]),
        .O(p_0_out[67]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[23]_i_5__0 
       (.I0(\block_w1_reg[23]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [87]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [87]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [87]),
        .O(\block_w1_reg[23]_i_5__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[23]_i_6 
       (.I0(\block_w1_reg[23]_i_7_n_0 ),
        .I1(\dec_block/op190_in [6]),
        .I2(\dec_block/op191_in [6]),
        .I3(\dec_block/op193_in [7]),
        .I4(\block_w3_reg[7]_i_12_n_0 ),
        .O(inv_mixcolumns_return0213_out__55[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[23]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [87]),
        .I1(\key_mem_reg[6]_6 [87]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [87]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [87]),
        .O(\block_w1_reg[23]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[23]_i_7 
       (.I0(\dec_block/op191_in [4]),
        .I1(\dec_block/p_0_in54_in [5]),
        .I2(\dec_block/op190_in [4]),
        .I3(\dec_block/op193_in [4]),
        .I4(\block_w0_reg[7]_i_4_n_0 ),
        .I5(\dec_block/op190_in [7]),
        .O(\block_w1_reg[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[23]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [87]),
        .I1(\key_mem_reg[2]_2 [87]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [87]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [87]),
        .O(\block_w1_reg[23]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[23]_i_8 
       (.I0(\key_mem_reg[11]_11 [87]),
        .I1(\key_mem_reg[10]_10 [87]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [87]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [87]),
        .O(\block_w1_reg[23]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[24]_i_2__0 
       (.I0(\dec_block/op161_in [0]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[24] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[24]_i_3 
       (.I0(\block_w1_reg[24]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[24]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[24]_i_7__0_n_0 ),
        .O(round_key[88]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[24]_i_4 
       (.I0(\block_w1_reg[24]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[24]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[24]_i_5__0_n_0 ),
        .I5(dec_new_block[88]),
        .O(\dec_block/op161_in [0]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[24]_i_5 
       (.I0(round_key[88]),
        .I1(core_block[88]),
        .O(p_0_out[38]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[24]_i_5__0 
       (.I0(\block_w1_reg[24]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [88]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [88]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [88]),
        .O(\block_w1_reg[24]_i_5__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[24]_i_6 
       (.I0(\block_w3_reg[8]_i_10_n_0 ),
        .I1(\dec_block/op158_in [0]),
        .I2(\block_w1_reg[24]_i_7_n_0 ),
        .I3(\block_w3_reg[8]_i_12_n_0 ),
        .I4(\block_w3_reg[11]_i_9_n_0 ),
        .O(inv_mixcolumns_return0188_out__55[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[24]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [88]),
        .I1(\key_mem_reg[6]_6 [88]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [88]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [88]),
        .O(\block_w1_reg[24]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[24]_i_7 
       (.I0(\dec_block/op159_in [7]),
        .I1(\dec_block/op161_in [7]),
        .O(\block_w1_reg[24]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[24]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [88]),
        .I1(\key_mem_reg[2]_2 [88]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [88]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [88]),
        .O(\block_w1_reg[24]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[24]_i_8 
       (.I0(\key_mem_reg[11]_11 [88]),
        .I1(\key_mem_reg[10]_10 [88]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [88]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [88]),
        .O(\block_w1_reg[24]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[25]_i_10 
       (.I0(\key_mem_reg[11]_11 [89]),
        .I1(\key_mem_reg[10]_10 [89]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [89]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [89]),
        .O(\block_w1_reg[25]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[25]_i_2__0 
       (.I0(\dec_block/op161_in [1]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[25] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[25]_i_3 
       (.I0(\block_w1_reg[25]_i_7_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[25]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[25]_i_9_n_0 ),
        .O(round_key[89]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[25]_i_4 
       (.I0(\block_w1_reg[25]_i_9_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[25]_i_8_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[25]_i_7_n_0 ),
        .I5(dec_new_block[89]),
        .O(\dec_block/op161_in [1]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[25]_i_5 
       (.I0(\block_w2_reg[16]_i_6_n_0 ),
        .I1(\block_w1_reg_reg[9] ),
        .I2(\block_w1_reg_reg[16] ),
        .I3(\block_w2_reg[16]_i_5_n_0 ),
        .I4(\block_w3_reg[12]_i_10_n_0 ),
        .I5(\dec_block/op161_in [0]),
        .O(inv_mixcolumns_return0188_out__55[1]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[25]_i_6 
       (.I0(round_key[89]),
        .I1(core_block[89]),
        .O(p_0_out[39]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[25]_i_7 
       (.I0(\block_w1_reg[25]_i_10_n_0 ),
        .I1(\key_mem_reg[14]_14 [89]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [89]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [89]),
        .O(\block_w1_reg[25]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[25]_i_8 
       (.I0(\key_mem_reg[7]_7 [89]),
        .I1(\key_mem_reg[6]_6 [89]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [89]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [89]),
        .O(\block_w1_reg[25]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[25]_i_9 
       (.I0(\key_mem_reg[3]_3 [89]),
        .I1(\key_mem_reg[2]_2 [89]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [89]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [89]),
        .O(\block_w1_reg[25]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[26]_i_3 
       (.I0(\block_w1_reg[26]_i_5__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w1_reg[26]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[26]_i_7_n_0 ),
        .O(round_key[90]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[26]_i_4 
       (.I0(round_key[90]),
        .I1(core_block[90]),
        .O(p_0_out[40]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[26]_i_5 
       (.I0(\block_w0_reg[0]_i_5_n_0 ),
        .I1(\block_w1_reg[26]_i_6_n_0 ),
        .I2(\dec_block/op159_in [7]),
        .I3(\block_w3_reg[14]_i_14_n_0 ),
        .I4(\block_w3_reg[13]_i_11_n_0 ),
        .I5(\dec_block/op161_in [1]),
        .O(inv_mixcolumns_return0188_out__55[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[26]_i_5__0 
       (.I0(\block_w1_reg[26]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [90]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [90]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [90]),
        .O(\block_w1_reg[26]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[26]_i_6 
       (.I0(\dec_block/op159_in [1]),
        .I1(\dec_block/op158_in [2]),
        .O(\block_w1_reg[26]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[26]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [90]),
        .I1(\key_mem_reg[6]_6 [90]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [90]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [90]),
        .O(\block_w1_reg[26]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[26]_i_7 
       (.I0(\key_mem_reg[3]_3 [90]),
        .I1(\key_mem_reg[2]_2 [90]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [90]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [90]),
        .O(\block_w1_reg[26]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[26]_i_8 
       (.I0(\key_mem_reg[11]_11 [90]),
        .I1(\key_mem_reg[10]_10 [90]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [90]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [90]),
        .O(\block_w1_reg[26]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[27]_i_10 
       (.I0(\key_mem_reg[11]_11 [91]),
        .I1(\key_mem_reg[10]_10 [91]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [91]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [91]),
        .O(\block_w1_reg[27]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[27]_i_3 
       (.I0(\block_w1_reg[27]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w1_reg[27]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[27]_i_8_n_0 ),
        .O(round_key[91]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[27]_i_4 
       (.I0(\block_w3_reg[14]_i_11_n_0 ),
        .I1(\block_w3_reg[11]_i_8_n_0 ),
        .I2(\dec_block/p_0_in46_in [4]),
        .I3(\dec_block/op161_in [2]),
        .I4(\block_w3_reg[12]_i_9_n_0 ),
        .I5(\block_w1_reg[27]_i_6_n_0 ),
        .O(inv_mixcolumns_return0188_out__55[3]));
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[27]_i_5 
       (.I0(round_key[91]),
        .I1(core_block[91]),
        .O(p_0_out[41]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[27]_i_5__0 
       (.I0(\block_w1_reg[26]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[26]_i_6__0_n_0 ),
        .I3(muxed_round_nr[3]),
        .I4(\block_w1_reg[26]_i_5__0_n_0 ),
        .I5(dec_new_block[90]),
        .O(\dec_block/op161_in [2]));
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w1_reg[27]_i_6 
       (.I0(dec_new_block[82]),
        .I1(round_key[82]),
        .I2(\dec_block/op158_in [6]),
        .I3(\dec_block/op161_in [6]),
        .O(\block_w1_reg[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[27]_i_6__0 
       (.I0(\block_w1_reg[27]_i_10_n_0 ),
        .I1(\key_mem_reg[14]_14 [91]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [91]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [91]),
        .O(\block_w1_reg[27]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[27]_i_7 
       (.I0(\key_mem_reg[7]_7 [91]),
        .I1(\key_mem_reg[6]_6 [91]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [91]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [91]),
        .O(\block_w1_reg[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[27]_i_8 
       (.I0(\key_mem_reg[3]_3 [91]),
        .I1(\key_mem_reg[2]_2 [91]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [91]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [91]),
        .O(\block_w1_reg[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[28]_i_10 
       (.I0(\key_mem_reg[11]_11 [92]),
        .I1(\key_mem_reg[10]_10 [92]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [92]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [92]),
        .O(\block_w1_reg[28]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[28]_i_2__0 
       (.I0(\dec_block/op161_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[28] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[28]_i_3 
       (.I0(\block_w1_reg[28]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[28]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[28]_i_8_n_0 ),
        .O(round_key[92]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[28]_i_4__0 
       (.I0(\block_w1_reg[28]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[28]_i_7__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[28]_i_6__0_n_0 ),
        .I5(dec_new_block[92]),
        .O(\dec_block/op161_in [4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[28]_i_5 
       (.I0(\block_w3_reg[13]_i_10_n_0 ),
        .I1(\block_w3_reg[12]_i_9_n_0 ),
        .I2(\block_w3_reg[12]_i_10_n_0 ),
        .I3(\block_w1_reg[28]_i_6_n_0 ),
        .I4(\block_w3_reg[12]_i_12_n_0 ),
        .I5(\block_w1_reg[28]_i_7_n_0 ),
        .O(inv_mixcolumns_return0188_out__55[4]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[28]_i_5__0 
       (.I0(round_key[92]),
        .I1(core_block[92]),
        .O(p_0_out[42]));
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w1_reg[28]_i_6 
       (.I0(\dec_block/op158_in [7]),
        .I1(round_key[83]),
        .I2(dec_new_block[83]),
        .I3(\dec_block/op158_in [4]),
        .O(\block_w1_reg[28]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[28]_i_6__0 
       (.I0(\block_w1_reg[28]_i_10_n_0 ),
        .I1(\key_mem_reg[14]_14 [92]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [92]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [92]),
        .O(\block_w1_reg[28]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \block_w1_reg[28]_i_7 
       (.I0(dec_new_block[91]),
        .I1(round_key[91]),
        .I2(\dec_block/op159_in [7]),
        .O(\block_w1_reg[28]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[28]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [92]),
        .I1(\key_mem_reg[6]_6 [92]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [92]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [92]),
        .O(\block_w1_reg[28]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[28]_i_8 
       (.I0(\key_mem_reg[3]_3 [92]),
        .I1(\key_mem_reg[2]_2 [92]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [92]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [92]),
        .O(\block_w1_reg[28]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[29]_i_2__0 
       (.I0(\dec_block/op161_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[29] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[29]_i_3 
       (.I0(\block_w1_reg[29]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[29]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[29]_i_7__0_n_0 ),
        .O(round_key[93]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[29]_i_4 
       (.I0(\block_w1_reg[29]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[29]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[29]_i_5__0_n_0 ),
        .I5(dec_new_block[93]),
        .O(\dec_block/op161_in [5]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[29]_i_5 
       (.I0(round_key[93]),
        .I1(core_block[93]),
        .O(p_0_out[43]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[29]_i_5__0 
       (.I0(\block_w1_reg[29]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [93]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [93]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [93]),
        .O(\block_w1_reg[29]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[29]_i_6 
       (.I0(\block_w3_reg[13]_i_10_n_0 ),
        .I1(\block_w3_reg[13]_i_11_n_0 ),
        .I2(\block_w1_reg[29]_i_7_n_0 ),
        .I3(\dec_block/op158_in [5]),
        .I4(\block_w3_reg[13]_i_13_n_0 ),
        .I5(\block_w3_reg[13]_i_14_n_0 ),
        .O(inv_mixcolumns_return0188_out__55[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[29]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [93]),
        .I1(\key_mem_reg[6]_6 [93]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [93]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [93]),
        .O(\block_w1_reg[29]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[29]_i_7 
       (.I0(\dec_block/op159_in [4]),
        .I1(\dec_block/op161_in [4]),
        .O(\block_w1_reg[29]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[29]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [93]),
        .I1(\key_mem_reg[2]_2 [93]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [93]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [93]),
        .O(\block_w1_reg[29]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[29]_i_8 
       (.I0(\key_mem_reg[11]_11 [93]),
        .I1(\key_mem_reg[10]_10 [93]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [93]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [93]),
        .O(\block_w1_reg[29]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[2]_i_2__0 
       (.I0(\dec_block/p_0_in46_in [3]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[2] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[2]_i_3 
       (.I0(\block_w1_reg[2]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[2]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[2]_i_7_n_0 ),
        .O(round_key[66]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[2]_i_4 
       (.I0(\block_w1_reg[2]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[2]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[2]_i_5__0_n_0 ),
        .I5(dec_new_block[66]),
        .O(\dec_block/p_0_in46_in [3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[2]_i_5 
       (.I0(round_key[34]),
        .I1(core_block[34]),
        .O(p_0_out[9]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[2]_i_5__0 
       (.I0(\block_w1_reg[2]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [66]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [66]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [66]),
        .O(\block_w1_reg[2]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[2]_i_6 
       (.I0(\block_w3_reg[21]_i_10_n_0 ),
        .I1(\dec_block/p_0_in38_in [2]),
        .I2(\dec_block/op129_in [1]),
        .I3(\block_w3_reg[18]_i_10_n_0 ),
        .I4(\block_w2_reg[24]_i_9_n_0 ),
        .I5(\block_w2_reg[27]_i_6_n_0 ),
        .O(inv_mixcolumns_return0134_out__63[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[2]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [66]),
        .I1(\key_mem_reg[6]_6 [66]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [66]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [66]),
        .O(\block_w1_reg[2]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[2]_i_7 
       (.I0(\key_mem_reg[3]_3 [66]),
        .I1(\key_mem_reg[2]_2 [66]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [66]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [66]),
        .O(\block_w1_reg[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[2]_i_8 
       (.I0(\key_mem_reg[11]_11 [66]),
        .I1(\key_mem_reg[10]_10 [66]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [66]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [66]),
        .O(\block_w1_reg[2]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[30]_i_2__0 
       (.I0(\dec_block/op161_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[30] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[30]_i_3 
       (.I0(\block_w1_reg[30]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[30]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[30]_i_7__0_n_0 ),
        .O(round_key[94]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[30]_i_4 
       (.I0(\block_w1_reg[30]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[30]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[30]_i_5__0_n_0 ),
        .I5(dec_new_block[94]),
        .O(\dec_block/op161_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[30]_i_5 
       (.I0(round_key[94]),
        .I1(core_block[94]),
        .O(p_0_out[44]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[30]_i_5__0 
       (.I0(\block_w1_reg[30]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [94]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [94]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [94]),
        .O(\block_w1_reg[30]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[30]_i_6 
       (.I0(\block_w3_reg[14]_i_10_n_0 ),
        .I1(\block_w3_reg[14]_i_11_n_0 ),
        .I2(\block_w3_reg[14]_i_12_n_0 ),
        .I3(\block_w1_reg[30]_i_7_n_0 ),
        .I4(\block_w3_reg[14]_i_14_n_0 ),
        .I5(\dec_block/op158_in [6]),
        .O(inv_mixcolumns_return0188_out__55[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[30]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [94]),
        .I1(\key_mem_reg[6]_6 [94]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [94]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [94]),
        .O(\block_w1_reg[30]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[30]_i_7 
       (.I0(\dec_block/op161_in [5]),
        .I1(\dec_block/op159_in [5]),
        .O(\block_w1_reg[30]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[30]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [94]),
        .I1(\key_mem_reg[2]_2 [94]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [94]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [94]),
        .O(\block_w1_reg[30]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[30]_i_8 
       (.I0(\key_mem_reg[11]_11 [94]),
        .I1(\key_mem_reg[10]_10 [94]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [94]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [94]),
        .O(\block_w1_reg[30]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[31]_i_3__0 
       (.I0(\dec_block/op161_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[31] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[31]_i_4 
       (.I0(\block_w1_reg[31]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[31]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[31]_i_8_n_0 ),
        .O(round_key[95]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[31]_i_5 
       (.I0(\block_w1_reg[31]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[31]_i_7__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[31]_i_6__0_n_0 ),
        .I5(dec_new_block[95]),
        .O(\dec_block/op161_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[31]_i_6 
       (.I0(round_key[95]),
        .I1(core_block[95]),
        .O(p_0_out[45]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[31]_i_6__0 
       (.I0(\block_w1_reg[31]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [95]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [95]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [95]),
        .O(\block_w1_reg[31]_i_6__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[31]_i_7 
       (.I0(\block_w2_reg[23]_i_7_n_0 ),
        .I1(\dec_block/op161_in [6]),
        .I2(\dec_block/op159_in [6]),
        .I3(\dec_block/op159_in [7]),
        .I4(\block_w3_reg[15]_i_12_n_0 ),
        .O(inv_mixcolumns_return0188_out__55[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[31]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [95]),
        .I1(\key_mem_reg[6]_6 [95]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [95]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [95]),
        .O(\block_w1_reg[31]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[31]_i_8 
       (.I0(\key_mem_reg[3]_3 [95]),
        .I1(\key_mem_reg[2]_2 [95]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [95]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [95]),
        .O(\block_w1_reg[31]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[31]_i_9 
       (.I0(\key_mem_reg[11]_11 [95]),
        .I1(\key_mem_reg[10]_10 [95]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [95]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [95]),
        .O(\block_w1_reg[31]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[3]_i_2__0 
       (.I0(\dec_block/p_0_in46_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[3] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[3]_i_3 
       (.I0(\block_w1_reg[3]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w1_reg[3]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[3]_i_8__0_n_0 ),
        .O(round_key[67]));
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[3]_i_4__0 
       (.I0(round_key[67]),
        .I1(dec_new_block[67]),
        .O(\dec_block/p_0_in46_in [4]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[3]_i_5 
       (.I0(round_key[67]),
        .I1(core_block[67]),
        .O(addroundkey_return[32]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[3]_i_5__0 
       (.I0(\block_w3_reg[19]_i_9_n_0 ),
        .I1(\block_w3_reg[20]_i_11_n_0 ),
        .I2(\block_w1_reg[3]_i_6_n_0 ),
        .I3(\block_w1_reg[3]_i_7_n_0 ),
        .I4(\block_w1_reg[3]_i_8_n_0 ),
        .I5(\block_w2_reg[28]_i_7_n_0 ),
        .O(inv_mixcolumns_return0134_out__63[2]));
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[3]_i_6 
       (.I0(\dec_block/op126_in [7]),
        .I1(round_key[51]),
        .I2(dec_new_block[51]),
        .I3(dec_new_block[43]),
        .I4(round_key[43]),
        .O(\block_w1_reg[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[3]_i_6__0 
       (.I0(\block_w1_reg[3]_i_9_n_0 ),
        .I1(\key_mem_reg[14]_14 [67]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [67]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [67]),
        .O(\block_w1_reg[3]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[3]_i_7 
       (.I0(\dec_block/p_0_in38_in [3]),
        .I1(\dec_block/op129_in [5]),
        .I2(\dec_block/op126_in [5]),
        .I3(\dec_block/p_0_in38_in [6]),
        .I4(\dec_block/op127_in [5]),
        .O(\block_w1_reg[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[3]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [67]),
        .I1(\key_mem_reg[6]_6 [67]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [67]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [67]),
        .O(\block_w1_reg[3]_i_7__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w1_reg[3]_i_8 
       (.I0(dec_new_block[58]),
        .I1(round_key[58]),
        .I2(\dec_block/op127_in [6]),
        .I3(\dec_block/p_0_in38_in [7]),
        .O(\block_w1_reg[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[3]_i_8__0 
       (.I0(\key_mem_reg[3]_3 [67]),
        .I1(\key_mem_reg[2]_2 [67]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [67]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [67]),
        .O(\block_w1_reg[3]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[3]_i_9 
       (.I0(\key_mem_reg[11]_11 [67]),
        .I1(\key_mem_reg[10]_10 [67]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [67]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [67]),
        .O(\block_w1_reg[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[4]_i_10 
       (.I0(\key_mem_reg[11]_11 [68]),
        .I1(\key_mem_reg[10]_10 [68]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [68]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [68]),
        .O(\block_w1_reg[4]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[4]_i_2__0 
       (.I0(\dec_block/p_0_in46_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[4] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[4]_i_3 
       (.I0(\block_w1_reg[4]_i_7_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[4]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[4]_i_9_n_0 ),
        .O(round_key[68]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[4]_i_4 
       (.I0(\block_w1_reg[4]_i_9_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[4]_i_8_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[4]_i_7_n_0 ),
        .I5(dec_new_block[68]),
        .O(\dec_block/p_0_in46_in [5]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[4]_i_5__0 
       (.I0(\block_w3_reg[20]_i_9_n_0 ),
        .I1(\dec_block/op127_in [4]),
        .I2(\block_w3_reg[20]_i_10_n_0 ),
        .I3(\block_w3_reg[20]_i_11_n_0 ),
        .I4(\block_w3_reg[21]_i_11_n_0 ),
        .I5(\block_w3_reg[22]_i_12_n_0 ),
        .O(inv_mixcolumns_return0134_out__63[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[4]_i_6 
       (.I0(round_key[68]),
        .I1(core_block[68]),
        .O(addroundkey_return[33]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[4]_i_7 
       (.I0(\block_w1_reg[4]_i_10_n_0 ),
        .I1(\key_mem_reg[14]_14 [68]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [68]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [68]),
        .O(\block_w1_reg[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[4]_i_8 
       (.I0(\key_mem_reg[7]_7 [68]),
        .I1(\key_mem_reg[6]_6 [68]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [68]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [68]),
        .O(\block_w1_reg[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[4]_i_9 
       (.I0(\key_mem_reg[3]_3 [68]),
        .I1(\key_mem_reg[2]_2 [68]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [68]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [68]),
        .O(\block_w1_reg[4]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[5]_i_2__0 
       (.I0(\dec_block/p_0_in46_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[5] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[5]_i_3 
       (.I0(\block_w1_reg[5]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[5]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[5]_i_7__0_n_0 ),
        .O(round_key[69]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[5]_i_4 
       (.I0(\block_w1_reg[5]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[5]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[5]_i_5__0_n_0 ),
        .I5(dec_new_block[69]),
        .O(\dec_block/p_0_in46_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[5]_i_5 
       (.I0(round_key[37]),
        .I1(core_block[37]),
        .O(p_0_out[12]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[5]_i_5__0 
       (.I0(\block_w1_reg[5]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [69]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [69]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [69]),
        .O(\block_w1_reg[5]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[5]_i_6 
       (.I0(\block_w3_reg[21]_i_10_n_0 ),
        .I1(\block_w3_reg[21]_i_11_n_0 ),
        .I2(\block_w1_reg[5]_i_7_n_0 ),
        .I3(\dec_block/op127_in [5]),
        .I4(\block_w3_reg[21]_i_13_n_0 ),
        .I5(\block_w3_reg[21]_i_14_n_0 ),
        .O(inv_mixcolumns_return0134_out__63[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[5]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [69]),
        .I1(\key_mem_reg[6]_6 [69]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [69]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [69]),
        .O(\block_w1_reg[5]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[5]_i_7 
       (.I0(\dec_block/p_0_in38_in [5]),
        .I1(\dec_block/op129_in [4]),
        .O(\block_w1_reg[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[5]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [69]),
        .I1(\key_mem_reg[2]_2 [69]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [69]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [69]),
        .O(\block_w1_reg[5]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[5]_i_8 
       (.I0(\key_mem_reg[11]_11 [69]),
        .I1(\key_mem_reg[10]_10 [69]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [69]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [69]),
        .O(\block_w1_reg[5]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[6]_i_2__0 
       (.I0(\dec_block/p_0_in46_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[6] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[6]_i_3 
       (.I0(\block_w1_reg[6]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[6]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[6]_i_7__0_n_0 ),
        .O(round_key[70]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[6]_i_4 
       (.I0(\block_w1_reg[6]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[6]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[6]_i_5__0_n_0 ),
        .I5(dec_new_block[70]),
        .O(\dec_block/p_0_in46_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[6]_i_5 
       (.I0(round_key[38]),
        .I1(core_block[38]),
        .O(p_0_out[13]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[6]_i_5__0 
       (.I0(\block_w1_reg[6]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [70]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [70]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [70]),
        .O(\block_w1_reg[6]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[6]_i_6 
       (.I0(\block_w3_reg[22]_i_10_n_0 ),
        .I1(\block_w3_reg[22]_i_11_n_0 ),
        .I2(\block_w3_reg[22]_i_12_n_0 ),
        .I3(\block_w1_reg[6]_i_7_n_0 ),
        .I4(\block_w3_reg[22]_i_14_n_0 ),
        .I5(\dec_block/op127_in [6]),
        .O(inv_mixcolumns_return0134_out__63[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[6]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [70]),
        .I1(\key_mem_reg[6]_6 [70]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [70]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [70]),
        .O(\block_w1_reg[6]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[6]_i_7 
       (.I0(\dec_block/op129_in [5]),
        .I1(\dec_block/p_0_in38_in [6]),
        .O(\block_w1_reg[6]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[6]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [70]),
        .I1(\key_mem_reg[2]_2 [70]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [70]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [70]),
        .O(\block_w1_reg[6]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[6]_i_8 
       (.I0(\key_mem_reg[11]_11 [70]),
        .I1(\key_mem_reg[10]_10 [70]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [70]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [70]),
        .O(\block_w1_reg[6]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[7]_i_2__0 
       (.I0(\block_w1_reg[7]_i_4_n_0 ),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[7] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[7]_i_3 
       (.I0(\block_w1_reg[7]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[7]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[7]_i_7__0_n_0 ),
        .O(round_key[71]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[7]_i_4 
       (.I0(\block_w1_reg[7]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[7]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[7]_i_5__0_n_0 ),
        .I5(dec_new_block[71]),
        .O(\block_w1_reg[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[7]_i_5 
       (.I0(round_key[39]),
        .I1(core_block[39]),
        .O(p_0_out[14]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[7]_i_5__0 
       (.I0(\block_w1_reg[7]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [71]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [71]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [71]),
        .O(\block_w1_reg[7]_i_5__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[7]_i_6 
       (.I0(\block_w1_reg[7]_i_7_n_0 ),
        .I1(\dec_block/op129_in [6]),
        .I2(\dec_block/p_0_in38_in [7]),
        .I3(\dec_block/op126_in [7]),
        .I4(\block_w3_reg[23]_i_12_n_0 ),
        .O(inv_mixcolumns_return0134_out__63[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[7]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [71]),
        .I1(\key_mem_reg[6]_6 [71]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [71]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [71]),
        .O(\block_w1_reg[7]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w1_reg[7]_i_7 
       (.I0(\dec_block/p_0_in38_in [5]),
        .I1(\dec_block/op127_in [4]),
        .I2(\dec_block/op126_in [4]),
        .I3(\dec_block/op129_in [4]),
        .I4(\dec_block/op129_in [7]),
        .I5(\dec_block/op127_in [7]),
        .O(\block_w1_reg[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[7]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [71]),
        .I1(\key_mem_reg[2]_2 [71]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [71]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [71]),
        .O(\block_w1_reg[7]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[7]_i_8 
       (.I0(\key_mem_reg[11]_11 [71]),
        .I1(\key_mem_reg[10]_10 [71]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [71]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [71]),
        .O(\block_w1_reg[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w1_reg[8]_i_2__0 
       (.I0(\dec_block/op158_in [0]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w1_reg_reg[8] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[8]_i_3 
       (.I0(\block_w1_reg[8]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[8]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[8]_i_7__0_n_0 ),
        .O(round_key[72]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[8]_i_4 
       (.I0(\block_w1_reg[8]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[8]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[8]_i_5__0_n_0 ),
        .I5(dec_new_block[72]),
        .O(\dec_block/op158_in [0]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[8]_i_5 
       (.I0(round_key[8]),
        .I1(core_block[8]),
        .O(addroundkey_return[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[8]_i_5__0 
       (.I0(\block_w1_reg[8]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [72]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [72]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [72]),
        .O(\block_w1_reg[8]_i_5__0_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w1_reg[8]_i_6 
       (.I0(\block_w3_reg[24]_i_10_n_0 ),
        .I1(\dec_block/op98_in [0]),
        .I2(\block_w1_reg[8]_i_7_n_0 ),
        .I3(\block_w3_reg[24]_i_12_n_0 ),
        .I4(\block_w3_reg[24]_i_13_n_0 ),
        .O(inv_mixcolumns_return0110_out__47[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[8]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [72]),
        .I1(\key_mem_reg[6]_6 [72]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [72]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [72]),
        .O(\block_w1_reg[8]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[8]_i_7 
       (.I0(\dec_block/op95_in [7]),
        .I1(\block_w3_reg[7]_i_4_n_0 ),
        .O(\block_w1_reg[8]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[8]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [72]),
        .I1(\key_mem_reg[2]_2 [72]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [72]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [72]),
        .O(\block_w1_reg[8]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[8]_i_8 
       (.I0(\key_mem_reg[11]_11 [72]),
        .I1(\key_mem_reg[10]_10 [72]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [72]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [72]),
        .O(\block_w1_reg[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[9]_i_10 
       (.I0(\key_mem_reg[11]_11 [73]),
        .I1(\key_mem_reg[10]_10 [73]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [73]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [73]),
        .O(\block_w1_reg[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \block_w1_reg[9]_i_3 
       (.I0(\block_w2_reg[0]_i_5_n_0 ),
        .I1(\block_w1_reg[9]_i_5_n_0 ),
        .I2(\block_w1_reg[9]_i_6__0_n_0 ),
        .I3(\dec_block/op95_in [0]),
        .I4(\block_w0_reg_reg[0]_1 ),
        .I5(\block_w0_reg_reg[16]_0 [1]),
        .O(\block_w3_reg_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w1_reg[9]_i_3__0 
       (.I0(\block_w1_reg[9]_i_7_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w1_reg[9]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w1_reg[9]_i_9_n_0 ),
        .O(round_key[73]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w1_reg[9]_i_4 
       (.I0(\block_w1_reg[9]_i_9_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[9]_i_8_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[9]_i_7_n_0 ),
        .I5(dec_new_block[73]),
        .O(\block_w1_reg_reg[9] ));
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w1_reg[9]_i_5 
       (.I0(\block_w3_reg_reg[0] ),
        .I1(\dec_block/op98_in [1]),
        .I2(\dec_block/op98_in [7]),
        .I3(\block_w3_reg[7]_i_4_n_0 ),
        .O(\block_w1_reg[9]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[9]_i_6 
       (.I0(round_key[73]),
        .I1(core_block[73]),
        .O(p_0_out[31]));
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w1_reg[9]_i_6__0 
       (.I0(\dec_block/op96_in [1]),
        .I1(\dec_block/p_0_in31_in [2]),
        .O(\block_w1_reg[9]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[9]_i_7 
       (.I0(\block_w1_reg[9]_i_10_n_0 ),
        .I1(\key_mem_reg[14]_14 [73]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [73]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [73]),
        .O(\block_w1_reg[9]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[9]_i_8 
       (.I0(\key_mem_reg[7]_7 [73]),
        .I1(\key_mem_reg[6]_6 [73]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [73]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [73]),
        .O(\block_w1_reg[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w1_reg[9]_i_9 
       (.I0(\key_mem_reg[3]_3 [73]),
        .I1(\key_mem_reg[2]_2 [73]),
        .I2(\block_w1_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [73]),
        .I4(\block_w1_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [73]),
        .O(\block_w1_reg[9]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[0]_i_11 
       (.I0(\key_mem_reg[11]_11 [32]),
        .I1(\key_mem_reg[10]_10 [32]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [32]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [32]),
        .O(\block_w2_reg[0]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT3 #(
    .INIT(8'h60)) 
    \block_w2_reg[0]_i_2__0 
       (.I0(round_key[0]),
        .I1(core_block[0]),
        .I2(\block_w0_reg_reg[0]_1 ),
        .O(\block_reg_reg[3][0] ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \block_w2_reg[0]_i_3 
       (.I0(\dec_block/op98_in [7]),
        .I1(\block_w3_reg_reg[16] ),
        .I2(\block_w2_reg[0]_i_5_n_0 ),
        .I3(\block_w2_reg[0]_i_6_n_0 ),
        .I4(\block_w0_reg_reg[0]_1 ),
        .I5(\block_w0_reg_reg[16]_0 [0]),
        .O(\block_w3_reg_reg[31]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[0]_i_3__0 
       (.I0(\block_w2_reg[0]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[0]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[0]_i_8_n_0 ),
        .O(round_key[32]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[0]_i_4 
       (.I0(\block_w2_reg[0]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[0]_i_7_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[0]_i_6__0_n_0 ),
        .I5(dec_new_block[32]),
        .O(\block_w2_reg_reg[0] ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[0]_i_5 
       (.I0(\dec_block/op95_in [5]),
        .I1(\dec_block/op98_in [5]),
        .I2(\dec_block/op96_in [5]),
        .I3(\dec_block/p_0_in31_in [6]),
        .I4(\dec_block/p_0_in31_in [7]),
        .I5(\dec_block/op96_in [6]),
        .O(\block_w2_reg[0]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \block_w2_reg[0]_i_6 
       (.I0(\dec_block/op98_in [0]),
        .I1(\dec_block/op95_in [0]),
        .I2(\block_w3_reg[7]_i_4_n_0 ),
        .O(\block_w2_reg[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[0]_i_6__0 
       (.I0(\block_w2_reg[0]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [32]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [32]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [32]),
        .O(\block_w2_reg[0]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[0]_i_7 
       (.I0(\key_mem_reg[7]_7 [32]),
        .I1(\key_mem_reg[6]_6 [32]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [32]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [32]),
        .O(\block_w2_reg[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[0]_i_8 
       (.I0(\key_mem_reg[3]_3 [32]),
        .I1(\key_mem_reg[2]_2 [32]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [32]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [32]),
        .O(\block_w2_reg[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[10]_i_11 
       (.I0(\key_mem_reg[11]_11 [42]),
        .I1(\key_mem_reg[10]_10 [42]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [42]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [42]),
        .O(\block_w2_reg[10]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[10]_i_2__0 
       (.I0(\dec_block/op126_in [2]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[10] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[10]_i_3 
       (.I0(\block_w2_reg[10]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[10]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[10]_i_8_n_0 ),
        .O(round_key[42]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[10]_i_4 
       (.I0(\block_w2_reg[10]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[10]_i_7_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[10]_i_6__0_n_0 ),
        .I5(dec_new_block[42]),
        .O(\dec_block/op126_in [2]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[10]_i_5 
       (.I0(round_key[106]),
        .I1(core_block[106]),
        .O(p_0_out[55]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[10]_i_6 
       (.I0(\block_w3_reg[5]_i_11_n_0 ),
        .I1(\block_w3_reg[0]_i_7_n_0 ),
        .I2(\dec_block/p_0_in54_in [2]),
        .I3(\dec_block/op191_in [7]),
        .I4(\block_w3_reg[3]_i_12_n_0 ),
        .I5(\dec_block/op190_in [1]),
        .O(inv_mixcolumns_return0206_out__55[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[10]_i_6__0 
       (.I0(\block_w2_reg[10]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [42]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [42]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [42]),
        .O(\block_w2_reg[10]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[10]_i_7 
       (.I0(\key_mem_reg[7]_7 [42]),
        .I1(\key_mem_reg[6]_6 [42]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [42]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [42]),
        .O(\block_w2_reg[10]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[10]_i_8 
       (.I0(\key_mem_reg[3]_3 [42]),
        .I1(\key_mem_reg[2]_2 [42]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [42]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [42]),
        .O(\block_w2_reg[10]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[11]_i_12 
       (.I0(\key_mem_reg[11]_11 [43]),
        .I1(\key_mem_reg[10]_10 [43]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [43]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [43]),
        .O(\block_w2_reg[11]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[11]_i_3 
       (.I0(\block_w2_reg[11]_i_7_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w2_reg[11]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[11]_i_9_n_0 ),
        .O(round_key[43]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[11]_i_4 
       (.I0(\block_w3_reg[3]_i_9_n_0 ),
        .I1(\block_w3_reg[4]_i_10_n_0 ),
        .I2(\block_w3_reg[6]_i_14_n_0 ),
        .I3(\block_w2_reg[11]_i_5_n_0 ),
        .I4(\block_w3_reg[6]_i_12_n_0 ),
        .I5(\dec_block/op191_in [3]),
        .O(inv_mixcolumns_return0206_out__55[2]));
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[11]_i_5 
       (.I0(\dec_block/op190_in [2]),
        .I1(\dec_block/p_0_in54_in [3]),
        .O(\block_w2_reg[11]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[11]_i_6 
       (.I0(round_key[43]),
        .I1(core_block[43]),
        .O(addroundkey_return[25]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[11]_i_7 
       (.I0(\block_w2_reg[11]_i_12_n_0 ),
        .I1(\key_mem_reg[14]_14 [43]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [43]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [43]),
        .O(\block_w2_reg[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[11]_i_8 
       (.I0(\key_mem_reg[7]_7 [43]),
        .I1(\key_mem_reg[6]_6 [43]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [43]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [43]),
        .O(\block_w2_reg[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[11]_i_9 
       (.I0(\key_mem_reg[3]_3 [43]),
        .I1(\key_mem_reg[2]_2 [43]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [43]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [43]),
        .O(\block_w2_reg[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[12]_i_12 
       (.I0(\key_mem_reg[11]_11 [44]),
        .I1(\key_mem_reg[10]_10 [44]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [44]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [44]),
        .O(\block_w2_reg[12]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[12]_i_2__0 
       (.I0(\dec_block/op126_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[12] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[12]_i_3 
       (.I0(\block_w2_reg[12]_i_7__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[12]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[12]_i_9_n_0 ),
        .O(round_key[44]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[12]_i_4__0 
       (.I0(\block_w2_reg[12]_i_9_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[12]_i_8_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[12]_i_7__0_n_0 ),
        .I5(dec_new_block[44]),
        .O(\dec_block/op126_in [4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[12]_i_5 
       (.I0(\block_w3_reg[5]_i_10_n_0 ),
        .I1(\block_w3_reg[4]_i_10_n_0 ),
        .I2(\block_w2_reg[9]_i_6_n_0 ),
        .I3(\block_w2_reg[12]_i_6_n_0 ),
        .I4(\block_w3_reg[6]_i_10_n_0 ),
        .I5(\block_w2_reg[12]_i_7_n_0 ),
        .O(inv_mixcolumns_return0206_out__55[3]));
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w2_reg[12]_i_6 
       (.I0(\block_w0_reg[7]_i_4_n_0 ),
        .I1(round_key[107]),
        .I2(dec_new_block[107]),
        .I3(\dec_block/op193_in [4]),
        .O(\block_w2_reg[12]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[12]_i_6__0 
       (.I0(round_key[44]),
        .I1(core_block[44]),
        .O(addroundkey_return[26]));
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \block_w2_reg[12]_i_7 
       (.I0(dec_new_block[99]),
        .I1(round_key[99]),
        .I2(\dec_block/op193_in [7]),
        .O(\block_w2_reg[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[12]_i_7__0 
       (.I0(\block_w2_reg[12]_i_12_n_0 ),
        .I1(\key_mem_reg[14]_14 [44]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [44]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [44]),
        .O(\block_w2_reg[12]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[12]_i_8 
       (.I0(\key_mem_reg[7]_7 [44]),
        .I1(\key_mem_reg[6]_6 [44]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [44]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [44]),
        .O(\block_w2_reg[12]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[12]_i_9 
       (.I0(\key_mem_reg[3]_3 [44]),
        .I1(\key_mem_reg[2]_2 [44]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [44]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [44]),
        .O(\block_w2_reg[12]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[13]_i_11 
       (.I0(\key_mem_reg[11]_11 [45]),
        .I1(\key_mem_reg[10]_10 [45]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [45]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [45]),
        .O(\block_w2_reg[13]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[13]_i_2__0 
       (.I0(\dec_block/op126_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[13] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[13]_i_3 
       (.I0(\block_w2_reg[13]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[13]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[13]_i_8__0_n_0 ),
        .O(round_key[45]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[13]_i_4 
       (.I0(\block_w2_reg[13]_i_8__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[13]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[13]_i_6__0_n_0 ),
        .I5(dec_new_block[45]),
        .O(\dec_block/op126_in [5]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[13]_i_5 
       (.I0(round_key[109]),
        .I1(core_block[109]),
        .O(p_0_out[58]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[13]_i_6 
       (.I0(\block_w3_reg[5]_i_10_n_0 ),
        .I1(\block_w3_reg[5]_i_11_n_0 ),
        .I2(\block_w2_reg[13]_i_7_n_0 ),
        .I3(\dec_block/op193_in [5]),
        .I4(\block_w3_reg[7]_i_12_n_0 ),
        .I5(\block_w2_reg[13]_i_8_n_0 ),
        .O(inv_mixcolumns_return0206_out__55[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[13]_i_6__0 
       (.I0(\block_w2_reg[13]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [45]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [45]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [45]),
        .O(\block_w2_reg[13]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[13]_i_7 
       (.I0(\dec_block/op190_in [4]),
        .I1(\dec_block/p_0_in54_in [5]),
        .O(\block_w2_reg[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[13]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [45]),
        .I1(\key_mem_reg[6]_6 [45]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [45]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [45]),
        .O(\block_w2_reg[13]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[13]_i_8 
       (.I0(\dec_block/op191_in [7]),
        .I1(round_key[123]),
        .I2(dec_new_block[123]),
        .I3(\block_w0_reg[7]_i_4_n_0 ),
        .I4(round_key[107]),
        .I5(dec_new_block[107]),
        .O(\block_w2_reg[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[13]_i_8__0 
       (.I0(\key_mem_reg[3]_3 [45]),
        .I1(\key_mem_reg[2]_2 [45]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [45]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [45]),
        .O(\block_w2_reg[13]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[14]_i_11 
       (.I0(\key_mem_reg[11]_11 [46]),
        .I1(\key_mem_reg[10]_10 [46]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [46]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [46]),
        .O(\block_w2_reg[14]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[14]_i_2__0 
       (.I0(\dec_block/op126_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[14] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[14]_i_3 
       (.I0(\block_w2_reg[14]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[14]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[14]_i_8__0_n_0 ),
        .O(round_key[46]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[14]_i_4 
       (.I0(\block_w2_reg[14]_i_8__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[14]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[14]_i_6__0_n_0 ),
        .I5(dec_new_block[46]),
        .O(\dec_block/op126_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[14]_i_5 
       (.I0(round_key[110]),
        .I1(core_block[110]),
        .O(p_0_out[59]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[14]_i_6 
       (.I0(\block_w3_reg[4]_i_9_n_0 ),
        .I1(\block_w3_reg[6]_i_11_n_0 ),
        .I2(\block_w3_reg[6]_i_12_n_0 ),
        .I3(\block_w2_reg[14]_i_7_n_0 ),
        .I4(\block_w2_reg[14]_i_8_n_0 ),
        .I5(\dec_block/op193_in [6]),
        .O(inv_mixcolumns_return0206_out__55[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[14]_i_6__0 
       (.I0(\block_w2_reg[14]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [46]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [46]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [46]),
        .O(\block_w2_reg[14]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[14]_i_7 
       (.I0(\dec_block/op190_in [5]),
        .I1(\dec_block/p_0_in54_in [6]),
        .O(\block_w2_reg[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[14]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [46]),
        .I1(\key_mem_reg[6]_6 [46]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [46]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [46]),
        .O(\block_w2_reg[14]_i_7__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[14]_i_8 
       (.I0(\dec_block/op191_in [6]),
        .I1(\dec_block/p_0_in54_in [7]),
        .O(\block_w2_reg[14]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[14]_i_8__0 
       (.I0(\key_mem_reg[3]_3 [46]),
        .I1(\key_mem_reg[2]_2 [46]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [46]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [46]),
        .O(\block_w2_reg[14]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[15]_i_12 
       (.I0(\key_mem_reg[11]_11 [47]),
        .I1(\key_mem_reg[10]_10 [47]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [47]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [47]),
        .O(\block_w2_reg[15]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[15]_i_2__0 
       (.I0(\dec_block/op126_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[15] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[15]_i_3 
       (.I0(\block_w2_reg[15]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[15]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[15]_i_8_n_0 ),
        .O(round_key[47]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[15]_i_4 
       (.I0(\block_w2_reg[15]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[15]_i_7_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[15]_i_6__0_n_0 ),
        .I5(dec_new_block[47]),
        .O(\dec_block/op126_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[15]_i_5 
       (.I0(round_key[111]),
        .I1(core_block[111]),
        .O(p_0_out[60]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[15]_i_6 
       (.I0(\block_w3_reg[7]_i_11_n_0 ),
        .I1(\dec_block/op190_in [6]),
        .I2(\dec_block/p_0_in54_in [7]),
        .I3(\block_w0_reg[7]_i_4_n_0 ),
        .I4(\block_w3_reg[5]_i_13_n_0 ),
        .O(inv_mixcolumns_return0206_out__55[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[15]_i_6__0 
       (.I0(\block_w2_reg[15]_i_12_n_0 ),
        .I1(\key_mem_reg[14]_14 [47]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [47]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [47]),
        .O(\block_w2_reg[15]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[15]_i_7 
       (.I0(\key_mem_reg[7]_7 [47]),
        .I1(\key_mem_reg[6]_6 [47]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [47]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [47]),
        .O(\block_w2_reg[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[15]_i_8 
       (.I0(\key_mem_reg[3]_3 [47]),
        .I1(\key_mem_reg[2]_2 [47]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [47]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [47]),
        .O(\block_w2_reg[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[16]_i_11 
       (.I0(\key_mem_reg[11]_11 [48]),
        .I1(\key_mem_reg[10]_10 [48]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [48]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [48]),
        .O(\block_w2_reg[16]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT3 #(
    .INIT(8'h60)) 
    \block_w2_reg[16]_i_2__0 
       (.I0(round_key[80]),
        .I1(core_block[80]),
        .I2(\block_w0_reg_reg[0]_1 ),
        .O(\block_reg_reg[1][16] ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \block_w2_reg[16]_i_3 
       (.I0(\block_w2_reg[16]_i_5_n_0 ),
        .I1(\block_w2_reg[16]_i_6_n_0 ),
        .I2(\block_w1_reg_reg[0] ),
        .I3(\block_w2_reg[16]_i_7_n_0 ),
        .I4(\block_w0_reg_reg[0]_1 ),
        .I5(\block_w0_reg_reg[16]_0 [2]),
        .O(\block_w1_reg_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[16]_i_3__0 
       (.I0(\block_w2_reg[16]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w2_reg[16]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[16]_i_8_n_0 ),
        .O(round_key[48]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[16]_i_4 
       (.I0(\block_w2_reg[16]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[16]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[16]_i_6__0_n_0 ),
        .I5(dec_new_block[48]),
        .O(\block_w2_reg_reg[16] ));
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[16]_i_5 
       (.I0(\dec_block/op158_in [7]),
        .I1(\dec_block/op159_in [7]),
        .O(\block_w2_reg[16]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[16]_i_6 
       (.I0(\dec_block/op159_in [5]),
        .I1(\dec_block/p_0_in46_in [6]),
        .I2(\dec_block/op161_in [5]),
        .I3(\dec_block/op158_in [5]),
        .I4(\dec_block/p_0_in46_in [7]),
        .I5(\dec_block/op159_in [6]),
        .O(\block_w2_reg[16]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[16]_i_6__0 
       (.I0(\block_w2_reg[16]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [48]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [48]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [48]),
        .O(\block_w2_reg[16]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[16]_i_7 
       (.I0(\dec_block/op161_in [0]),
        .I1(\dec_block/op158_in [0]),
        .O(\block_w2_reg[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[16]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [48]),
        .I1(\key_mem_reg[6]_6 [48]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [48]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [48]),
        .O(\block_w2_reg[16]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[16]_i_8 
       (.I0(\key_mem_reg[3]_3 [48]),
        .I1(\key_mem_reg[2]_2 [48]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [48]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [48]),
        .O(\block_w2_reg[16]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[17]_i_12 
       (.I0(\key_mem_reg[11]_11 [49]),
        .I1(\key_mem_reg[10]_10 [49]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [49]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [49]),
        .O(\block_w2_reg[17]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[17]_i_2__0 
       (.I0(\dec_block/op127_in [1]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[17] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[17]_i_3 
       (.I0(\block_w2_reg[17]_i_7_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[17]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[17]_i_9_n_0 ),
        .O(round_key[49]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[17]_i_4__0 
       (.I0(\block_w2_reg[17]_i_9_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[17]_i_8_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[17]_i_7_n_0 ),
        .I5(dec_new_block[49]),
        .O(\dec_block/op127_in [1]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[17]_i_5 
       (.I0(\dec_block/op158_in [0]),
        .I1(\dec_block/p_0_in46_in [2]),
        .I2(\block_w3_reg[12]_i_9_n_0 ),
        .I3(\block_w3_reg[11]_i_9_n_0 ),
        .I4(\block_w1_reg_reg[16] ),
        .I5(\block_w3_reg[8]_i_11_n_0 ),
        .O(inv_mixcolumns_return0181_out__58[0]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[17]_i_6 
       (.I0(round_key[49]),
        .I1(core_block[49]),
        .O(p_0_out[15]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[17]_i_7 
       (.I0(\block_w2_reg[17]_i_12_n_0 ),
        .I1(\key_mem_reg[14]_14 [49]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [49]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [49]),
        .O(\block_w2_reg[17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[17]_i_8 
       (.I0(\key_mem_reg[7]_7 [49]),
        .I1(\key_mem_reg[6]_6 [49]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [49]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [49]),
        .O(\block_w2_reg[17]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[17]_i_9 
       (.I0(\key_mem_reg[3]_3 [49]),
        .I1(\key_mem_reg[2]_2 [49]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [49]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [49]),
        .O(\block_w2_reg[17]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[18]_i_11 
       (.I0(\key_mem_reg[11]_11 [50]),
        .I1(\key_mem_reg[10]_10 [50]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [50]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [50]),
        .O(\block_w2_reg[18]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[18]_i_3 
       (.I0(\block_w2_reg[18]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w2_reg[18]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[18]_i_8_n_0 ),
        .O(round_key[50]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[18]_i_4 
       (.I0(round_key[82]),
        .I1(core_block[82]),
        .O(addroundkey_return[38]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[18]_i_5 
       (.I0(\block_w2_reg[18]_i_6_n_0 ),
        .I1(\dec_block/p_0_in46_in [3]),
        .I2(\dec_block/op159_in [1]),
        .I3(\block_w2_reg[18]_i_7_n_0 ),
        .I4(\block_w3_reg[13]_i_10_n_0 ),
        .I5(\block_w1_reg_reg[9] ),
        .O(inv_mixcolumns_return0181_out__58[1]));
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w2_reg[18]_i_6 
       (.I0(\block_w1_reg_reg[0] ),
        .I1(\block_w1_reg_reg[16] ),
        .I2(\dec_block/op158_in [6]),
        .I3(\dec_block/op161_in [6]),
        .O(\block_w2_reg[18]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[18]_i_6__0 
       (.I0(\block_w2_reg[18]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [50]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [50]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [50]),
        .O(\block_w2_reg[18]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[18]_i_7 
       (.I0(\dec_block/op158_in [7]),
        .I1(\dec_block/op161_in [7]),
        .O(\block_w2_reg[18]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[18]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [50]),
        .I1(\key_mem_reg[6]_6 [50]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [50]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [50]),
        .O(\block_w2_reg[18]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[18]_i_8 
       (.I0(\key_mem_reg[3]_3 [50]),
        .I1(\key_mem_reg[2]_2 [50]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [50]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [50]),
        .O(\block_w2_reg[18]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[19]_i_12 
       (.I0(\key_mem_reg[11]_11 [51]),
        .I1(\key_mem_reg[10]_10 [51]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [51]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [51]),
        .O(\block_w2_reg[19]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[19]_i_2__0 
       (.I0(\dec_block/op127_in [3]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[19] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[19]_i_3 
       (.I0(\block_w2_reg[19]_i_7__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w2_reg[19]_i_8__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[19]_i_9_n_0 ),
        .O(round_key[51]));
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[19]_i_4__0 
       (.I0(round_key[51]),
        .I1(dec_new_block[51]),
        .O(\dec_block/op127_in [3]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[19]_i_5 
       (.I0(\block_w2_reg[16]_i_6_n_0 ),
        .I1(\block_w3_reg[11]_i_8_n_0 ),
        .I2(\block_w2_reg[19]_i_6_n_0 ),
        .I3(\block_w3_reg[12]_i_10_n_0 ),
        .I4(\block_w3_reg[12]_i_13_n_0 ),
        .O(inv_mixcolumns_return0181_out__58[2]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[19]_i_6 
       (.I0(\dec_block/op159_in [2]),
        .I1(dec_new_block[75]),
        .I2(round_key[75]),
        .I3(\block_w1_reg[7]_i_4_n_0 ),
        .I4(\dec_block/op158_in [2]),
        .I5(\dec_block/op161_in [3]),
        .O(\block_w2_reg[19]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[19]_i_6__0 
       (.I0(round_key[51]),
        .I1(core_block[51]),
        .O(p_0_out[17]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[19]_i_7 
       (.I0(\block_w1_reg[18]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[18]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[18]_i_5__0_n_0 ),
        .I5(dec_new_block[82]),
        .O(\dec_block/op159_in [2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[19]_i_7__0 
       (.I0(\block_w2_reg[19]_i_12_n_0 ),
        .I1(\key_mem_reg[14]_14 [51]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [51]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [51]),
        .O(\block_w2_reg[19]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[19]_i_8 
       (.I0(\block_w1_reg[27]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w1_reg[27]_i_7_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w1_reg[27]_i_6__0_n_0 ),
        .I5(dec_new_block[91]),
        .O(\dec_block/op161_in [3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[19]_i_8__0 
       (.I0(\key_mem_reg[7]_7 [51]),
        .I1(\key_mem_reg[6]_6 [51]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [51]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [51]),
        .O(\block_w2_reg[19]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[19]_i_9 
       (.I0(\key_mem_reg[3]_3 [51]),
        .I1(\key_mem_reg[2]_2 [51]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [51]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [51]),
        .O(\block_w2_reg[19]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[1]_i_12 
       (.I0(\key_mem_reg[11]_11 [33]),
        .I1(\key_mem_reg[10]_10 [33]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [33]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [33]),
        .O(\block_w2_reg[1]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[1]_i_2__0 
       (.I0(\dec_block/p_0_in38_in [2]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[1] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[1]_i_3 
       (.I0(\block_w2_reg[1]_i_7_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w2_reg[1]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[1]_i_9_n_0 ),
        .O(round_key[33]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[1]_i_4__0 
       (.I0(\block_w2_reg[1]_i_9_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[1]_i_8_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[1]_i_7_n_0 ),
        .I5(dec_new_block[33]),
        .O(\dec_block/p_0_in38_in [2]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[1]_i_5 
       (.I0(\block_w3_reg_reg[0] ),
        .I1(\dec_block/op96_in [1]),
        .I2(\block_w3_reg[28]_i_9_n_0 ),
        .I3(\block_w3_reg[24]_i_13_n_0 ),
        .I4(\dec_block/op98_in [0]),
        .I5(\block_w3_reg[24]_i_11_n_0 ),
        .O(inv_mixcolumns_return0__55[0]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[1]_i_6 
       (.I0(round_key[33]),
        .I1(core_block[33]),
        .O(p_0_out[8]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[1]_i_7 
       (.I0(\block_w2_reg[1]_i_12_n_0 ),
        .I1(\key_mem_reg[14]_14 [33]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [33]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [33]),
        .O(\block_w2_reg[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[1]_i_8 
       (.I0(\key_mem_reg[7]_7 [33]),
        .I1(\key_mem_reg[6]_6 [33]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [33]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [33]),
        .O(\block_w2_reg[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[1]_i_9 
       (.I0(\key_mem_reg[3]_3 [33]),
        .I1(\key_mem_reg[2]_2 [33]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [33]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [33]),
        .O(\block_w2_reg[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[20]_i_10 
       (.I0(\key_mem_reg[3]_3 [52]),
        .I1(\key_mem_reg[2]_2 [52]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [52]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [52]),
        .O(\block_w2_reg[20]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[20]_i_13 
       (.I0(\key_mem_reg[11]_11 [52]),
        .I1(\key_mem_reg[10]_10 [52]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [52]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [52]),
        .O(\block_w2_reg[20]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[20]_i_2__0 
       (.I0(\dec_block/op127_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[20] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[20]_i_3 
       (.I0(\block_w2_reg[20]_i_8_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[20]_i_9_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[20]_i_10_n_0 ),
        .O(round_key[52]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[20]_i_4 
       (.I0(\block_w2_reg[20]_i_10_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[20]_i_9_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[20]_i_8_n_0 ),
        .I5(dec_new_block[52]),
        .O(\dec_block/op127_in [4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[20]_i_5 
       (.I0(\block_w3_reg[14]_i_10_n_0 ),
        .I1(\dec_block/p_0_in46_in [5]),
        .I2(\block_w3_reg[12]_i_9_n_0 ),
        .I3(\block_w3_reg[12]_i_10_n_0 ),
        .I4(\block_w3_reg[13]_i_11_n_0 ),
        .I5(\block_w3_reg[14]_i_11_n_0 ),
        .O(inv_mixcolumns_return0181_out__58[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[20]_i_7 
       (.I0(round_key[52]),
        .I1(core_block[52]),
        .O(p_0_out[18]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[20]_i_8 
       (.I0(\block_w2_reg[20]_i_13_n_0 ),
        .I1(\key_mem_reg[14]_14 [52]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [52]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [52]),
        .O(\block_w2_reg[20]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[20]_i_9 
       (.I0(\key_mem_reg[7]_7 [52]),
        .I1(\key_mem_reg[6]_6 [52]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [52]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [52]),
        .O(\block_w2_reg[20]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[21]_i_11 
       (.I0(\key_mem_reg[11]_11 [53]),
        .I1(\key_mem_reg[10]_10 [53]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [53]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [53]),
        .O(\block_w2_reg[21]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[21]_i_2__0 
       (.I0(\dec_block/op127_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[21] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[21]_i_3 
       (.I0(\block_w2_reg[21]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[21]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[21]_i_8__0_n_0 ),
        .O(round_key[53]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[21]_i_4 
       (.I0(\block_w2_reg[21]_i_8__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[21]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[21]_i_6__0_n_0 ),
        .I5(dec_new_block[53]),
        .O(\dec_block/op127_in [5]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[21]_i_5 
       (.I0(round_key[85]),
        .I1(core_block[85]),
        .O(addroundkey_return[41]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[21]_i_6 
       (.I0(\block_w3_reg[13]_i_10_n_0 ),
        .I1(\block_w3_reg[13]_i_11_n_0 ),
        .I2(\block_w2_reg[21]_i_7_n_0 ),
        .I3(\dec_block/p_0_in46_in [6]),
        .I4(\block_w3_reg[15]_i_12_n_0 ),
        .I5(\block_w2_reg[21]_i_8_n_0 ),
        .O(inv_mixcolumns_return0181_out__58[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[21]_i_6__0 
       (.I0(\block_w2_reg[21]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [53]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [53]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [53]),
        .O(\block_w2_reg[21]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[21]_i_7 
       (.I0(\dec_block/op158_in [4]),
        .I1(\dec_block/op159_in [4]),
        .O(\block_w2_reg[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[21]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [53]),
        .I1(\key_mem_reg[6]_6 [53]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [53]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [53]),
        .O(\block_w2_reg[21]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[21]_i_8 
       (.I0(\dec_block/op161_in [7]),
        .I1(round_key[67]),
        .I2(dec_new_block[67]),
        .I3(\dec_block/op158_in [7]),
        .I4(round_key[83]),
        .I5(dec_new_block[83]),
        .O(\block_w2_reg[21]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[21]_i_8__0 
       (.I0(\key_mem_reg[3]_3 [53]),
        .I1(\key_mem_reg[2]_2 [53]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [53]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [53]),
        .O(\block_w2_reg[21]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[22]_i_11 
       (.I0(\key_mem_reg[11]_11 [54]),
        .I1(\key_mem_reg[10]_10 [54]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [54]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [54]),
        .O(\block_w2_reg[22]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[22]_i_2__0 
       (.I0(\dec_block/op127_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[22] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[22]_i_3 
       (.I0(\block_w2_reg[22]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[22]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[22]_i_8_n_0 ),
        .O(round_key[54]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[22]_i_4 
       (.I0(\block_w2_reg[22]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[22]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[22]_i_6__0_n_0 ),
        .I5(dec_new_block[54]),
        .O(\dec_block/op127_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[22]_i_5 
       (.I0(round_key[86]),
        .I1(core_block[86]),
        .O(addroundkey_return[42]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[22]_i_6 
       (.I0(\block_w3_reg[12]_i_12_n_0 ),
        .I1(\block_w3_reg[14]_i_11_n_0 ),
        .I2(\block_w3_reg[14]_i_12_n_0 ),
        .I3(\block_w2_reg[22]_i_7_n_0 ),
        .I4(\block_w3_reg[11]_i_9_n_0 ),
        .I5(\dec_block/p_0_in46_in [7]),
        .O(inv_mixcolumns_return0181_out__58[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[22]_i_6__0 
       (.I0(\block_w2_reg[22]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [54]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [54]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [54]),
        .O(\block_w2_reg[22]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[22]_i_7 
       (.I0(\dec_block/op159_in [5]),
        .I1(\dec_block/op158_in [5]),
        .O(\block_w2_reg[22]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[22]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [54]),
        .I1(\key_mem_reg[6]_6 [54]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [54]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [54]),
        .O(\block_w2_reg[22]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[22]_i_8 
       (.I0(\key_mem_reg[3]_3 [54]),
        .I1(\key_mem_reg[2]_2 [54]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [54]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [54]),
        .O(\block_w2_reg[22]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[23]_i_12 
       (.I0(\key_mem_reg[11]_11 [55]),
        .I1(\key_mem_reg[10]_10 [55]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [55]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [55]),
        .O(\block_w2_reg[23]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[23]_i_2__0 
       (.I0(\dec_block/op127_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[23] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[23]_i_3 
       (.I0(\block_w2_reg[23]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[23]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[23]_i_8_n_0 ),
        .O(round_key[55]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[23]_i_4 
       (.I0(\block_w2_reg[23]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[23]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[23]_i_6__0_n_0 ),
        .I5(dec_new_block[55]),
        .O(\dec_block/op127_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[23]_i_5 
       (.I0(round_key[87]),
        .I1(core_block[87]),
        .O(addroundkey_return[43]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[23]_i_6 
       (.I0(\block_w2_reg[23]_i_7_n_0 ),
        .I1(\dec_block/op158_in [6]),
        .I2(\dec_block/op159_in [6]),
        .I3(\dec_block/op161_in [7]),
        .I4(\block_w3_reg[13]_i_13_n_0 ),
        .O(inv_mixcolumns_return0181_out__58[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[23]_i_6__0 
       (.I0(\block_w2_reg[23]_i_12_n_0 ),
        .I1(\key_mem_reg[14]_14 [55]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [55]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [55]),
        .O(\block_w2_reg[23]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[23]_i_7 
       (.I0(\dec_block/op159_in [4]),
        .I1(\dec_block/p_0_in46_in [5]),
        .I2(\dec_block/op158_in [4]),
        .I3(\dec_block/op161_in [4]),
        .I4(\dec_block/op158_in [7]),
        .I5(\block_w1_reg[7]_i_4_n_0 ),
        .O(\block_w2_reg[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[23]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [55]),
        .I1(\key_mem_reg[6]_6 [55]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [55]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [55]),
        .O(\block_w2_reg[23]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[23]_i_8 
       (.I0(\key_mem_reg[3]_3 [55]),
        .I1(\key_mem_reg[2]_2 [55]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [55]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [55]),
        .O(\block_w2_reg[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[24]_i_11 
       (.I0(\key_mem_reg[11]_11 [56]),
        .I1(\key_mem_reg[10]_10 [56]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [56]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [56]),
        .O(\block_w2_reg[24]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[24]_i_2__0 
       (.I0(\dec_block/op129_in [0]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[24] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[24]_i_3 
       (.I0(\block_w2_reg[24]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[24]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[24]_i_8__0_n_0 ),
        .O(round_key[56]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[24]_i_4 
       (.I0(\block_w2_reg[24]_i_8__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[24]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[24]_i_6__0_n_0 ),
        .I5(dec_new_block[56]),
        .O(\dec_block/op129_in [0]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[24]_i_5 
       (.I0(round_key[56]),
        .I1(core_block[56]),
        .O(p_0_out[22]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[24]_i_6 
       (.I0(\block_w2_reg[24]_i_7_n_0 ),
        .I1(\dec_block/op126_in [0]),
        .I2(\block_w2_reg[24]_i_8_n_0 ),
        .I3(\block_w2_reg[24]_i_9_n_0 ),
        .I4(\block_w3_reg[22]_i_14_n_0 ),
        .O(inv_mixcolumns_return0156_out__63[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[24]_i_6__0 
       (.I0(\block_w2_reg[24]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [56]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [56]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [56]),
        .O(\block_w2_reg[24]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w2_reg[24]_i_7 
       (.I0(\dec_block/op127_in [5]),
        .I1(\dec_block/p_0_in38_in [6]),
        .I2(\dec_block/op126_in [5]),
        .I3(\dec_block/op129_in [5]),
        .O(\block_w2_reg[24]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[24]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [56]),
        .I1(\key_mem_reg[6]_6 [56]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [56]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [56]),
        .O(\block_w2_reg[24]_i_7__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[24]_i_8 
       (.I0(\dec_block/op127_in [7]),
        .I1(\dec_block/op129_in [7]),
        .O(\block_w2_reg[24]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[24]_i_8__0 
       (.I0(\key_mem_reg[3]_3 [56]),
        .I1(\key_mem_reg[2]_2 [56]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [56]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [56]),
        .O(\block_w2_reg[24]_i_8__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[24]_i_9 
       (.I0(\block_w2_reg_reg[0] ),
        .I1(\block_w2_reg_reg[16] ),
        .O(\block_w2_reg[24]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[25]_i_10 
       (.I0(\key_mem_reg[3]_3 [57]),
        .I1(\key_mem_reg[2]_2 [57]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [57]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [57]),
        .O(\block_w2_reg[25]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[25]_i_13 
       (.I0(\key_mem_reg[11]_11 [57]),
        .I1(\key_mem_reg[10]_10 [57]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [57]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [57]),
        .O(\block_w2_reg[25]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[25]_i_2__0 
       (.I0(\dec_block/op129_in [1]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[25] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[25]_i_3 
       (.I0(\block_w2_reg[25]_i_8_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[25]_i_9_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[25]_i_10_n_0 ),
        .O(round_key[57]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[25]_i_4 
       (.I0(\block_w2_reg[25]_i_10_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[25]_i_9_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[25]_i_8_n_0 ),
        .I5(dec_new_block[57]),
        .O(\dec_block/op129_in [1]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[25]_i_5 
       (.I0(\block_w3_reg[16]_i_7_n_0 ),
        .I1(\block_w2_reg_reg[16] ),
        .I2(\block_w2_reg_reg[9] ),
        .I3(\block_w3_reg[16]_i_6_n_0 ),
        .I4(\block_w3_reg[20]_i_11_n_0 ),
        .I5(\dec_block/op129_in [0]),
        .O(inv_mixcolumns_return0156_out__63[1]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[25]_i_7 
       (.I0(round_key[57]),
        .I1(core_block[57]),
        .O(p_0_out[23]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[25]_i_8 
       (.I0(\block_w2_reg[25]_i_13_n_0 ),
        .I1(\key_mem_reg[14]_14 [57]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [57]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [57]),
        .O(\block_w2_reg[25]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[25]_i_9 
       (.I0(\key_mem_reg[7]_7 [57]),
        .I1(\key_mem_reg[6]_6 [57]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [57]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [57]),
        .O(\block_w2_reg[25]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[26]_i_11 
       (.I0(\key_mem_reg[11]_11 [58]),
        .I1(\key_mem_reg[10]_10 [58]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [58]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [58]),
        .O(\block_w2_reg[26]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[26]_i_3 
       (.I0(\block_w2_reg[26]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w2_reg[26]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[26]_i_8_n_0 ),
        .O(round_key[58]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[26]_i_4 
       (.I0(round_key[58]),
        .I1(core_block[58]),
        .O(p_0_out[24]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[26]_i_5 
       (.I0(\block_w1_reg[0]_i_5_n_0 ),
        .I1(\block_w2_reg[26]_i_6_n_0 ),
        .I2(\dec_block/op127_in [7]),
        .I3(\block_w2_reg[30]_i_8_n_0 ),
        .I4(\block_w3_reg[21]_i_11_n_0 ),
        .I5(\dec_block/op129_in [1]),
        .O(inv_mixcolumns_return0156_out__63[2]));
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[26]_i_6 
       (.I0(\dec_block/op126_in [2]),
        .I1(\dec_block/op127_in [1]),
        .O(\block_w2_reg[26]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[26]_i_6__0 
       (.I0(\block_w2_reg[26]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [58]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [58]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [58]),
        .O(\block_w2_reg[26]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[26]_i_7 
       (.I0(\key_mem_reg[7]_7 [58]),
        .I1(\key_mem_reg[6]_6 [58]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [58]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [58]),
        .O(\block_w2_reg[26]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[26]_i_8 
       (.I0(\key_mem_reg[3]_3 [58]),
        .I1(\key_mem_reg[2]_2 [58]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [58]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [58]),
        .O(\block_w2_reg[26]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[27]_i_10 
       (.I0(\key_mem_reg[3]_3 [59]),
        .I1(\key_mem_reg[2]_2 [59]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [59]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [59]),
        .O(\block_w2_reg[27]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[27]_i_14 
       (.I0(\key_mem_reg[11]_11 [59]),
        .I1(\key_mem_reg[10]_10 [59]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [59]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [59]),
        .O(\block_w2_reg[27]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[27]_i_3 
       (.I0(\block_w2_reg[27]_i_7_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w2_reg[27]_i_9_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[27]_i_10_n_0 ),
        .O(round_key[59]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[27]_i_4 
       (.I0(\block_w3_reg[22]_i_11_n_0 ),
        .I1(\block_w3_reg[19]_i_9_n_0 ),
        .I2(\dec_block/p_0_in38_in [4]),
        .I3(\dec_block/op129_in [2]),
        .I4(\block_w3_reg[20]_i_10_n_0 ),
        .I5(\block_w2_reg[27]_i_6_n_0 ),
        .O(inv_mixcolumns_return0156_out__63[3]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[27]_i_5 
       (.I0(\block_w2_reg[26]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[26]_i_7_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[26]_i_6__0_n_0 ),
        .I5(dec_new_block[58]),
        .O(\dec_block/op129_in [2]));
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w2_reg[27]_i_6 
       (.I0(dec_new_block[50]),
        .I1(round_key[50]),
        .I2(\dec_block/op126_in [6]),
        .I3(\dec_block/op129_in [6]),
        .O(\block_w2_reg[27]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[27]_i_6__0 
       (.I0(round_key[59]),
        .I1(core_block[59]),
        .O(p_0_out[25]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[27]_i_7 
       (.I0(\block_w2_reg[27]_i_14_n_0 ),
        .I1(\key_mem_reg[14]_14 [59]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [59]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [59]),
        .O(\block_w2_reg[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[27]_i_9 
       (.I0(\key_mem_reg[7]_7 [59]),
        .I1(\key_mem_reg[6]_6 [59]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [59]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [59]),
        .O(\block_w2_reg[27]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[28]_i_13 
       (.I0(\key_mem_reg[11]_11 [60]),
        .I1(\key_mem_reg[10]_10 [60]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [60]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [60]),
        .O(\block_w2_reg[28]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[28]_i_2__0 
       (.I0(\dec_block/op129_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[28] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[28]_i_3 
       (.I0(\block_w2_reg[28]_i_7__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[28]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[28]_i_9_n_0 ),
        .O(round_key[60]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[28]_i_4__0 
       (.I0(\block_w2_reg[28]_i_9_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[28]_i_8_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[28]_i_7__0_n_0 ),
        .I5(dec_new_block[60]),
        .O(\dec_block/op129_in [4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[28]_i_5 
       (.I0(\block_w3_reg[21]_i_10_n_0 ),
        .I1(\block_w3_reg[20]_i_10_n_0 ),
        .I2(\block_w3_reg[20]_i_11_n_0 ),
        .I3(\block_w2_reg[28]_i_6__0_n_0 ),
        .I4(\block_w3_reg[22]_i_10_n_0 ),
        .I5(\block_w2_reg[28]_i_7_n_0 ),
        .O(inv_mixcolumns_return0156_out__63[4]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[28]_i_6 
       (.I0(round_key[60]),
        .I1(core_block[60]),
        .O(p_0_out[26]));
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w2_reg[28]_i_6__0 
       (.I0(\dec_block/op126_in [7]),
        .I1(round_key[51]),
        .I2(dec_new_block[51]),
        .I3(\dec_block/op126_in [4]),
        .O(\block_w2_reg[28]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \block_w2_reg[28]_i_7 
       (.I0(dec_new_block[59]),
        .I1(round_key[59]),
        .I2(\dec_block/op127_in [7]),
        .O(\block_w2_reg[28]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[28]_i_7__0 
       (.I0(\block_w2_reg[28]_i_13_n_0 ),
        .I1(\key_mem_reg[14]_14 [60]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [60]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [60]),
        .O(\block_w2_reg[28]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[28]_i_8 
       (.I0(\key_mem_reg[7]_7 [60]),
        .I1(\key_mem_reg[6]_6 [60]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [60]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [60]),
        .O(\block_w2_reg[28]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[28]_i_9 
       (.I0(\key_mem_reg[3]_3 [60]),
        .I1(\key_mem_reg[2]_2 [60]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [60]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [60]),
        .O(\block_w2_reg[28]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[29]_i_11 
       (.I0(\key_mem_reg[11]_11 [61]),
        .I1(\key_mem_reg[10]_10 [61]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [61]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [61]),
        .O(\block_w2_reg[29]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[29]_i_2__0 
       (.I0(\dec_block/op129_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[29] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[29]_i_3 
       (.I0(\block_w2_reg[29]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[29]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[29]_i_8__0_n_0 ),
        .O(round_key[61]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[29]_i_4 
       (.I0(\block_w2_reg[29]_i_8__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[29]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[29]_i_6__0_n_0 ),
        .I5(dec_new_block[61]),
        .O(\dec_block/op129_in [5]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[29]_i_5 
       (.I0(round_key[61]),
        .I1(core_block[61]),
        .O(p_0_out[27]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[29]_i_6 
       (.I0(\block_w3_reg[21]_i_10_n_0 ),
        .I1(\block_w3_reg[21]_i_11_n_0 ),
        .I2(\block_w2_reg[29]_i_7_n_0 ),
        .I3(\dec_block/op126_in [5]),
        .I4(\block_w3_reg[23]_i_12_n_0 ),
        .I5(\block_w2_reg[29]_i_8_n_0 ),
        .O(inv_mixcolumns_return0156_out__63[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[29]_i_6__0 
       (.I0(\block_w2_reg[29]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [61]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [61]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [61]),
        .O(\block_w2_reg[29]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[29]_i_7 
       (.I0(\dec_block/op127_in [4]),
        .I1(\dec_block/op129_in [4]),
        .O(\block_w2_reg[29]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[29]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [61]),
        .I1(\key_mem_reg[6]_6 [61]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [61]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [61]),
        .O(\block_w2_reg[29]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[29]_i_8 
       (.I0(\dec_block/op127_in [7]),
        .I1(round_key[59]),
        .I2(dec_new_block[59]),
        .I3(\block_w2_reg[7]_i_4_n_0 ),
        .I4(round_key[43]),
        .I5(dec_new_block[43]),
        .O(\block_w2_reg[29]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[29]_i_8__0 
       (.I0(\key_mem_reg[3]_3 [61]),
        .I1(\key_mem_reg[2]_2 [61]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [61]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [61]),
        .O(\block_w2_reg[29]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[2]_i_11 
       (.I0(\key_mem_reg[11]_11 [34]),
        .I1(\key_mem_reg[10]_10 [34]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [34]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [34]),
        .O(\block_w2_reg[2]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[2]_i_2__0 
       (.I0(\dec_block/p_0_in38_in [3]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[2] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[2]_i_3 
       (.I0(\block_w2_reg[2]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[2]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[2]_i_8_n_0 ),
        .O(round_key[34]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[2]_i_4 
       (.I0(\block_w2_reg[2]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[2]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[2]_i_6__0_n_0 ),
        .I5(dec_new_block[34]),
        .O(\dec_block/p_0_in38_in [3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[2]_i_5 
       (.I0(round_key[2]),
        .I1(core_block[2]),
        .O(addroundkey_return[1]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[2]_i_6 
       (.I0(\block_w3_reg[29]_i_10_n_0 ),
        .I1(\dec_block/p_0_in31_in [2]),
        .I2(\dec_block/op98_in [1]),
        .I3(\block_w2_reg[2]_i_7_n_0 ),
        .I4(\block_w3_reg[24]_i_12_n_0 ),
        .I5(\block_w3_reg[27]_i_10_n_0 ),
        .O(inv_mixcolumns_return0__55[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[2]_i_6__0 
       (.I0(\block_w2_reg[2]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [34]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [34]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [34]),
        .O(\block_w2_reg[2]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[2]_i_7 
       (.I0(\dec_block/op95_in [7]),
        .I1(\dec_block/op98_in [7]),
        .O(\block_w2_reg[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[2]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [34]),
        .I1(\key_mem_reg[6]_6 [34]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [34]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [34]),
        .O(\block_w2_reg[2]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[2]_i_8 
       (.I0(\key_mem_reg[3]_3 [34]),
        .I1(\key_mem_reg[2]_2 [34]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [34]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [34]),
        .O(\block_w2_reg[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[30]_i_11 
       (.I0(\key_mem_reg[11]_11 [62]),
        .I1(\key_mem_reg[10]_10 [62]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [62]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [62]),
        .O(\block_w2_reg[30]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[30]_i_2__0 
       (.I0(\dec_block/op129_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[30] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[30]_i_3 
       (.I0(\block_w2_reg[30]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[30]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[30]_i_8__0_n_0 ),
        .O(round_key[62]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[30]_i_4 
       (.I0(\block_w2_reg[30]_i_8__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[30]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[30]_i_6__0_n_0 ),
        .I5(dec_new_block[62]),
        .O(\dec_block/op129_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[30]_i_5 
       (.I0(round_key[62]),
        .I1(core_block[62]),
        .O(p_0_out[28]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[30]_i_6 
       (.I0(\block_w3_reg[20]_i_9_n_0 ),
        .I1(\block_w3_reg[22]_i_11_n_0 ),
        .I2(\block_w3_reg[22]_i_12_n_0 ),
        .I3(\block_w2_reg[30]_i_7_n_0 ),
        .I4(\block_w2_reg[30]_i_8_n_0 ),
        .I5(\dec_block/op126_in [6]),
        .O(inv_mixcolumns_return0156_out__63[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[30]_i_6__0 
       (.I0(\block_w2_reg[30]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [62]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [62]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [62]),
        .O(\block_w2_reg[30]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[30]_i_7 
       (.I0(\dec_block/op129_in [5]),
        .I1(\dec_block/op127_in [5]),
        .O(\block_w2_reg[30]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[30]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [62]),
        .I1(\key_mem_reg[6]_6 [62]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [62]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [62]),
        .O(\block_w2_reg[30]_i_7__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[30]_i_8 
       (.I0(\dec_block/p_0_in38_in [7]),
        .I1(\dec_block/op127_in [6]),
        .O(\block_w2_reg[30]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[30]_i_8__0 
       (.I0(\key_mem_reg[3]_3 [62]),
        .I1(\key_mem_reg[2]_2 [62]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [62]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [62]),
        .O(\block_w2_reg[30]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[31]_i_11 
       (.I0(\block_w2_reg[31]_i_19_n_0 ),
        .I1(\key_mem_reg[14]_14 [63]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [63]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [63]),
        .O(\block_w2_reg[31]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[31]_i_13 
       (.I0(\key_mem_reg[7]_7 [63]),
        .I1(\key_mem_reg[6]_6 [63]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [63]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [63]),
        .O(\block_w2_reg[31]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[31]_i_15 
       (.I0(\key_mem_reg[3]_3 [63]),
        .I1(\key_mem_reg[2]_2 [63]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [63]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [63]),
        .O(\block_w2_reg[31]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[31]_i_19 
       (.I0(\key_mem_reg[11]_11 [63]),
        .I1(\key_mem_reg[10]_10 [63]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [63]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [63]),
        .O(\block_w2_reg[31]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \block_w2_reg[31]_i_21 
       (.I0(muxed_round_nr[2]),
        .I1(\block_w0_reg[31]_i_6__0_1 ),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .O(\block_w2_reg[31]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[31]_i_3__0 
       (.I0(\dec_block/op129_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[31] ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[31]_i_5 
       (.I0(\block_w2_reg[31]_i_15_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[31]_i_13_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[31]_i_11_n_0 ),
        .I5(dec_new_block[63]),
        .O(\dec_block/op129_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[31]_i_6__0 
       (.I0(round_key[63]),
        .I1(core_block[63]),
        .O(p_0_out[29]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[31]_i_7 
       (.I0(\block_w3_reg[23]_i_11_n_0 ),
        .I1(\dec_block/op129_in [6]),
        .I2(\dec_block/op127_in [6]),
        .I3(\dec_block/op127_in [7]),
        .I4(\block_w3_reg[21]_i_13_n_0 ),
        .O(inv_mixcolumns_return0156_out__63[7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[31]_i_7__0 
       (.I0(\block_w2_reg[31]_i_11_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[31]_i_13_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[31]_i_15_n_0 ),
        .O(round_key[63]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[3]_i_12 
       (.I0(\key_mem_reg[11]_11 [35]),
        .I1(\key_mem_reg[10]_10 [35]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [35]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [35]),
        .O(\block_w2_reg[3]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[3]_i_2__0 
       (.I0(\dec_block/p_0_in38_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[3] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[3]_i_3 
       (.I0(\block_w2_reg[3]_i_7__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w2_reg[3]_i_8__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[3]_i_9_n_0 ),
        .O(round_key[35]));
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[3]_i_4__0 
       (.I0(round_key[35]),
        .I1(dec_new_block[35]),
        .O(\dec_block/p_0_in38_in [4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[3]_i_5 
       (.I0(\block_w3_reg[27]_i_8_n_0 ),
        .I1(\block_w1_reg[9]_i_6__0_n_0 ),
        .I2(\block_w2_reg[3]_i_6__0_n_0 ),
        .I3(\block_w2_reg[3]_i_7_n_0 ),
        .I4(\block_w2_reg[3]_i_8_n_0 ),
        .I5(\block_w3_reg[28]_i_12_n_0 ),
        .O(inv_mixcolumns_return0__55[2]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[3]_i_6 
       (.I0(round_key[35]),
        .I1(core_block[35]),
        .O(p_0_out[10]));
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[3]_i_6__0 
       (.I0(\dec_block/op95_in [7]),
        .I1(round_key[19]),
        .I2(dec_new_block[19]),
        .I3(dec_new_block[11]),
        .I4(round_key[11]),
        .O(\block_w2_reg[3]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[3]_i_7 
       (.I0(\dec_block/p_0_in31_in [3]),
        .I1(\dec_block/op95_in [5]),
        .I2(\dec_block/op98_in [5]),
        .I3(\dec_block/op96_in [5]),
        .I4(\dec_block/p_0_in31_in [6]),
        .O(\block_w2_reg[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[3]_i_7__0 
       (.I0(\block_w2_reg[3]_i_12_n_0 ),
        .I1(\key_mem_reg[14]_14 [35]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [35]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [35]),
        .O(\block_w2_reg[3]_i_7__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w2_reg[3]_i_8 
       (.I0(dec_new_block[26]),
        .I1(round_key[26]),
        .I2(\dec_block/p_0_in31_in [7]),
        .I3(\dec_block/op96_in [6]),
        .O(\block_w2_reg[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[3]_i_8__0 
       (.I0(\key_mem_reg[7]_7 [35]),
        .I1(\key_mem_reg[6]_6 [35]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [35]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [35]),
        .O(\block_w2_reg[3]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[3]_i_9 
       (.I0(\key_mem_reg[3]_3 [35]),
        .I1(\key_mem_reg[2]_2 [35]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [35]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [35]),
        .O(\block_w2_reg[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[4]_i_10 
       (.I0(\key_mem_reg[3]_3 [36]),
        .I1(\key_mem_reg[2]_2 [36]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [36]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [36]),
        .O(\block_w2_reg[4]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[4]_i_13 
       (.I0(\key_mem_reg[11]_11 [36]),
        .I1(\key_mem_reg[10]_10 [36]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [36]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [36]),
        .O(\block_w2_reg[4]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[4]_i_2__0 
       (.I0(\dec_block/p_0_in38_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[4] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[4]_i_3 
       (.I0(\block_w2_reg[4]_i_8_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[4]_i_9_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[4]_i_10_n_0 ),
        .O(round_key[36]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[4]_i_4 
       (.I0(\block_w2_reg[4]_i_10_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[4]_i_9_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[4]_i_8_n_0 ),
        .I5(dec_new_block[36]),
        .O(\dec_block/p_0_in38_in [5]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[4]_i_5__0 
       (.I0(\block_w3_reg[30]_i_10_n_0 ),
        .I1(\dec_block/op96_in [4]),
        .I2(\block_w3_reg[28]_i_9_n_0 ),
        .I3(\block_w1_reg[9]_i_6__0_n_0 ),
        .I4(\block_w3_reg[29]_i_11_n_0 ),
        .I5(\block_w3_reg[30]_i_12_n_0 ),
        .O(inv_mixcolumns_return0__55[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[4]_i_7 
       (.I0(round_key[36]),
        .I1(core_block[36]),
        .O(p_0_out[11]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[4]_i_8 
       (.I0(\block_w2_reg[4]_i_13_n_0 ),
        .I1(\key_mem_reg[14]_14 [36]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [36]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [36]),
        .O(\block_w2_reg[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[4]_i_9 
       (.I0(\key_mem_reg[7]_7 [36]),
        .I1(\key_mem_reg[6]_6 [36]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [36]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [36]),
        .O(\block_w2_reg[4]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[5]_i_11 
       (.I0(\key_mem_reg[11]_11 [37]),
        .I1(\key_mem_reg[10]_10 [37]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [37]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [37]),
        .O(\block_w2_reg[5]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[5]_i_2__0 
       (.I0(\dec_block/p_0_in38_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[5] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[5]_i_3 
       (.I0(\block_w2_reg[5]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[5]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[5]_i_8__0_n_0 ),
        .O(round_key[37]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[5]_i_4 
       (.I0(\block_w2_reg[5]_i_8__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[5]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[5]_i_6__0_n_0 ),
        .I5(dec_new_block[37]),
        .O(\dec_block/p_0_in38_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[5]_i_5 
       (.I0(round_key[5]),
        .I1(core_block[5]),
        .O(addroundkey_return[4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[5]_i_6 
       (.I0(\block_w3_reg[29]_i_10_n_0 ),
        .I1(\block_w3_reg[29]_i_11_n_0 ),
        .I2(\block_w2_reg[5]_i_7_n_0 ),
        .I3(\dec_block/op96_in [5]),
        .I4(\block_w3_reg[31]_i_14_n_0 ),
        .I5(\block_w2_reg[5]_i_8_n_0 ),
        .O(inv_mixcolumns_return0__55[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[5]_i_6__0 
       (.I0(\block_w2_reg[5]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [37]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [37]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [37]),
        .O(\block_w2_reg[5]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[5]_i_7 
       (.I0(\dec_block/p_0_in31_in [5]),
        .I1(\dec_block/op98_in [4]),
        .O(\block_w2_reg[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[5]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [37]),
        .I1(\key_mem_reg[6]_6 [37]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [37]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [37]),
        .O(\block_w2_reg[5]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[5]_i_8 
       (.I0(\dec_block/op98_in [7]),
        .I1(round_key[3]),
        .I2(dec_new_block[3]),
        .I3(\dec_block/op95_in [7]),
        .I4(round_key[19]),
        .I5(dec_new_block[19]),
        .O(\block_w2_reg[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[5]_i_8__0 
       (.I0(\key_mem_reg[3]_3 [37]),
        .I1(\key_mem_reg[2]_2 [37]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [37]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [37]),
        .O(\block_w2_reg[5]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[6]_i_11 
       (.I0(\key_mem_reg[11]_11 [38]),
        .I1(\key_mem_reg[10]_10 [38]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [38]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [38]),
        .O(\block_w2_reg[6]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[6]_i_2__0 
       (.I0(\dec_block/p_0_in38_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[6] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[6]_i_3 
       (.I0(\block_w2_reg[6]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[6]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[6]_i_8_n_0 ),
        .O(round_key[38]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[6]_i_4 
       (.I0(\block_w2_reg[6]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[6]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[6]_i_6__0_n_0 ),
        .I5(dec_new_block[38]),
        .O(\dec_block/p_0_in38_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[6]_i_5 
       (.I0(round_key[6]),
        .I1(core_block[6]),
        .O(addroundkey_return[5]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[6]_i_6 
       (.I0(\block_w3_reg[28]_i_11_n_0 ),
        .I1(\block_w3_reg[30]_i_11_n_0 ),
        .I2(\block_w3_reg[30]_i_12_n_0 ),
        .I3(\block_w2_reg[6]_i_7_n_0 ),
        .I4(\block_w3_reg[24]_i_13_n_0 ),
        .I5(\dec_block/op96_in [6]),
        .O(inv_mixcolumns_return0__55[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[6]_i_6__0 
       (.I0(\block_w2_reg[6]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [38]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [38]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [38]),
        .O(\block_w2_reg[6]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[6]_i_7 
       (.I0(\dec_block/op98_in [5]),
        .I1(\dec_block/p_0_in31_in [6]),
        .O(\block_w2_reg[6]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[6]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [38]),
        .I1(\key_mem_reg[6]_6 [38]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [38]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [38]),
        .O(\block_w2_reg[6]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[6]_i_8 
       (.I0(\key_mem_reg[3]_3 [38]),
        .I1(\key_mem_reg[2]_2 [38]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [38]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [38]),
        .O(\block_w2_reg[6]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[7]_i_12 
       (.I0(\key_mem_reg[11]_11 [39]),
        .I1(\key_mem_reg[10]_10 [39]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [39]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [39]),
        .O(\block_w2_reg[7]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[7]_i_2__0 
       (.I0(\block_w2_reg[7]_i_4_n_0 ),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[7] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[7]_i_3 
       (.I0(\block_w2_reg[7]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[7]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[7]_i_8_n_0 ),
        .O(round_key[39]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[7]_i_4 
       (.I0(\block_w2_reg[7]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[7]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[7]_i_6__0_n_0 ),
        .I5(dec_new_block[39]),
        .O(\block_w2_reg[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[7]_i_5 
       (.I0(round_key[7]),
        .I1(core_block[7]),
        .O(addroundkey_return[6]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[7]_i_6 
       (.I0(\block_w2_reg[7]_i_7_n_0 ),
        .I1(\dec_block/op98_in [6]),
        .I2(\dec_block/p_0_in31_in [7]),
        .I3(\dec_block/op95_in [7]),
        .I4(\block_w3_reg[29]_i_13_n_0 ),
        .O(inv_mixcolumns_return0__55[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[7]_i_6__0 
       (.I0(\block_w2_reg[7]_i_12_n_0 ),
        .I1(\key_mem_reg[14]_14 [39]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [39]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [39]),
        .O(\block_w2_reg[7]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w2_reg[7]_i_7 
       (.I0(\dec_block/op96_in [4]),
        .I1(\dec_block/p_0_in31_in [5]),
        .I2(\dec_block/op95_in [4]),
        .I3(\dec_block/op98_in [4]),
        .I4(\dec_block/op98_in [7]),
        .I5(\dec_block/op96_in [7]),
        .O(\block_w2_reg[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[7]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [39]),
        .I1(\key_mem_reg[6]_6 [39]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [39]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [39]),
        .O(\block_w2_reg[7]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[7]_i_8 
       (.I0(\key_mem_reg[3]_3 [39]),
        .I1(\key_mem_reg[2]_2 [39]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [39]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [39]),
        .O(\block_w2_reg[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[8]_i_11 
       (.I0(\key_mem_reg[11]_11 [40]),
        .I1(\key_mem_reg[10]_10 [40]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [40]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [40]),
        .O(\block_w2_reg[8]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w2_reg[8]_i_2__0 
       (.I0(\dec_block/op126_in [0]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w2_reg_reg[8] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[8]_i_3 
       (.I0(\block_w2_reg[8]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w2_reg[8]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[8]_i_8__0_n_0 ),
        .O(round_key[40]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[8]_i_4 
       (.I0(\block_w2_reg[8]_i_8__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[8]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[8]_i_6__0_n_0 ),
        .I5(dec_new_block[40]),
        .O(\dec_block/op126_in [0]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[8]_i_5 
       (.I0(round_key[104]),
        .I1(core_block[104]),
        .O(p_0_out[53]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w2_reg[8]_i_6 
       (.I0(\block_w2_reg[8]_i_7_n_0 ),
        .I1(\dec_block/op193_in [0]),
        .I2(\block_w2_reg[8]_i_8_n_0 ),
        .I3(\block_w3_reg[2]_i_11_n_0 ),
        .I4(\block_w3_reg[6]_i_14_n_0 ),
        .O(inv_mixcolumns_return0206_out__55[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[8]_i_6__0 
       (.I0(\block_w2_reg[8]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [40]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [40]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [40]),
        .O(\block_w2_reg[8]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w2_reg[8]_i_7 
       (.I0(\dec_block/op193_in [5]),
        .I1(\dec_block/op190_in [5]),
        .I2(\dec_block/p_0_in54_in [6]),
        .I3(\dec_block/op191_in [5]),
        .O(\block_w2_reg[8]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[8]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [40]),
        .I1(\key_mem_reg[6]_6 [40]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [40]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [40]),
        .O(\block_w2_reg[8]_i_7__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[8]_i_8 
       (.I0(\dec_block/op190_in [7]),
        .I1(\block_w0_reg[7]_i_4_n_0 ),
        .O(\block_w2_reg[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[8]_i_8__0 
       (.I0(\key_mem_reg[3]_3 [40]),
        .I1(\key_mem_reg[2]_2 [40]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [40]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [40]),
        .O(\block_w2_reg[8]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[9]_i_10 
       (.I0(\key_mem_reg[3]_3 [41]),
        .I1(\key_mem_reg[2]_2 [41]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [41]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [41]),
        .O(\block_w2_reg[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[9]_i_13 
       (.I0(\key_mem_reg[11]_11 [41]),
        .I1(\key_mem_reg[10]_10 [41]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [41]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [41]),
        .O(\block_w2_reg[9]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \block_w2_reg[9]_i_3 
       (.I0(\block_w3_reg[0]_i_6_n_0 ),
        .I1(\block_w2_reg[9]_i_5_n_0 ),
        .I2(\block_w2_reg[9]_i_6_n_0 ),
        .I3(\dec_block/op190_in [0]),
        .I4(\block_w0_reg_reg[0]_1 ),
        .I5(\block_w0_reg_reg[16]_0 [1]),
        .O(\block_w0_reg_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w2_reg[9]_i_3__0 
       (.I0(\block_w2_reg[9]_i_8_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w2_reg[9]_i_9_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w2_reg[9]_i_10_n_0 ),
        .O(round_key[41]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[9]_i_4 
       (.I0(\block_w2_reg[9]_i_10_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[9]_i_9_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[9]_i_8_n_0 ),
        .I5(dec_new_block[41]),
        .O(\block_w2_reg_reg[9] ));
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w2_reg[9]_i_5 
       (.I0(\dec_block/op193_in [1]),
        .I1(\block_w0_reg_reg[0] ),
        .I2(\dec_block/op193_in [7]),
        .I3(\block_w0_reg[7]_i_4_n_0 ),
        .O(\block_w2_reg[9]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[9]_i_6 
       (.I0(\dec_block/op191_in [1]),
        .I1(\dec_block/p_0_in54_in [2]),
        .O(\block_w2_reg[9]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w2_reg[9]_i_7 
       (.I0(\block_w0_reg[8]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[8]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[8]_i_5__0_n_0 ),
        .I5(dec_new_block[104]),
        .O(\dec_block/op190_in [0]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w2_reg[9]_i_7__0 
       (.I0(round_key[41]),
        .I1(core_block[41]),
        .O(addroundkey_return[23]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[9]_i_8 
       (.I0(\block_w2_reg[9]_i_13_n_0 ),
        .I1(\key_mem_reg[14]_14 [41]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [41]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [41]),
        .O(\block_w2_reg[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w2_reg[9]_i_9 
       (.I0(\key_mem_reg[7]_7 [41]),
        .I1(\key_mem_reg[6]_6 [41]),
        .I2(\block_w2_reg[29]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [41]),
        .I4(\block_w2_reg[29]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [41]),
        .O(\block_w2_reg[9]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT3 #(
    .INIT(8'h60)) 
    \block_w3_reg[0]_i_2__0 
       (.I0(round_key[96]),
        .I1(core_block[96]),
        .I2(\block_w0_reg_reg[0]_1 ),
        .O(\block_reg_reg[0][0] ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \block_w3_reg[0]_i_3 
       (.I0(\dec_block/op193_in [7]),
        .I1(\block_w0_reg_reg[16] ),
        .I2(\block_w3_reg[0]_i_6_n_0 ),
        .I3(\block_w3_reg[0]_i_7_n_0 ),
        .I4(\block_w0_reg_reg[0]_1 ),
        .I5(\block_w0_reg_reg[16]_0 [0]),
        .O(\block_w0_reg_reg[31]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[0]_i_3__0 
       (.I0(\block_w3_reg[0]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[0]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[0]_i_7__0_n_0 ),
        .O(round_key[0]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[0]_i_4 
       (.I0(\block_w3_reg[0]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[0]_i_6__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w3_reg[0]_i_5__0_n_0 ),
        .I5(dec_new_block[0]),
        .O(\block_w3_reg_reg[0] ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[0]_i_5 
       (.I0(\block_w0_reg[31]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w0_reg[31]_i_7_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w0_reg[31]_i_6__0_n_0 ),
        .I5(dec_new_block[127]),
        .O(\dec_block/op193_in [7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[0]_i_5__0 
       (.I0(\block_w3_reg[0]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [0]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [0]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [0]),
        .O(\block_w3_reg[0]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[0]_i_6 
       (.I0(\dec_block/op191_in [5]),
        .I1(\dec_block/p_0_in54_in [6]),
        .I2(\dec_block/op190_in [5]),
        .I3(\dec_block/op193_in [5]),
        .I4(\dec_block/p_0_in54_in [7]),
        .I5(\dec_block/op191_in [6]),
        .O(\block_w3_reg[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[0]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [0]),
        .I1(\key_mem_reg[6]_6 [0]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [0]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [0]),
        .O(\block_w3_reg[0]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \block_w3_reg[0]_i_7 
       (.I0(\dec_block/op193_in [0]),
        .I1(\dec_block/op190_in [0]),
        .I2(\block_w0_reg[7]_i_4_n_0 ),
        .O(\block_w3_reg[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[0]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [0]),
        .I1(\key_mem_reg[2]_2 [0]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [0]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [0]),
        .O(\block_w3_reg[0]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[0]_i_8 
       (.I0(\key_mem_reg[11]_11 [0]),
        .I1(\key_mem_reg[10]_10 [0]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [0]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [0]),
        .O(\block_w3_reg[0]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w3_reg[10]_i_10 
       (.I0(dec_new_block[90]),
        .I1(round_key[90]),
        .I2(\dec_block/p_0_in46_in [7]),
        .I3(\dec_block/op159_in [6]),
        .O(\block_w3_reg[10]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[10]_i_2__0 
       (.I0(\dec_block/op95_in [2]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[10] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[10]_i_3 
       (.I0(\block_w3_reg[10]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[10]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[10]_i_7__0_n_0 ),
        .O(round_key[10]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[10]_i_4 
       (.I0(\block_w3_reg[10]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[10]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[10]_i_5__0_n_0 ),
        .I5(dec_new_block[10]),
        .O(\dec_block/op95_in [2]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[10]_i_5 
       (.I0(round_key[74]),
        .I1(core_block[74]),
        .O(p_0_out[32]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[10]_i_5__0 
       (.I0(\block_w3_reg[10]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [10]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [10]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [10]),
        .O(\block_w3_reg[10]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[10]_i_6 
       (.I0(\key_mem_reg[7]_7 [10]),
        .I1(\key_mem_reg[6]_6 [10]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [10]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [10]),
        .O(\block_w3_reg[10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[10]_i_7 
       (.I0(\block_w3_reg[13]_i_11_n_0 ),
        .I1(\block_w0_reg[0]_i_5_n_0 ),
        .I2(\dec_block/p_0_in46_in [2]),
        .I3(\dec_block/op159_in [7]),
        .I4(\block_w3_reg[10]_i_10_n_0 ),
        .I5(\block_w1_reg_reg[9] ),
        .O(inv_mixcolumns_return0174_out__63[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[10]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [10]),
        .I1(\key_mem_reg[2]_2 [10]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [10]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [10]),
        .O(\block_w3_reg[10]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[10]_i_8 
       (.I0(\key_mem_reg[11]_11 [10]),
        .I1(\key_mem_reg[10]_10 [10]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [10]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [10]),
        .O(\block_w3_reg[10]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[11]_i_10 
       (.I0(\dec_block/op158_in [2]),
        .I1(\dec_block/p_0_in46_in [3]),
        .O(\block_w3_reg[11]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[11]_i_3 
       (.I0(\block_w3_reg[11]_i_6_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w3_reg[11]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[11]_i_8__0_n_0 ),
        .O(round_key[11]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[11]_i_5 
       (.I0(\block_w3_reg[11]_i_8_n_0 ),
        .I1(\block_w3_reg[12]_i_9_n_0 ),
        .I2(\block_w3_reg[11]_i_9_n_0 ),
        .I3(\block_w3_reg[11]_i_10_n_0 ),
        .I4(\block_w3_reg[14]_i_12_n_0 ),
        .I5(\dec_block/op159_in [3]),
        .O(inv_mixcolumns_return0174_out__63[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[11]_i_5__0 
       (.I0(round_key[11]),
        .I1(core_block[11]),
        .O(addroundkey_return[10]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[11]_i_6 
       (.I0(\block_w3_reg[11]_i_9__0_n_0 ),
        .I1(\key_mem_reg[14]_14 [11]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [11]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [11]),
        .O(\block_w3_reg[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[11]_i_7 
       (.I0(\key_mem_reg[7]_7 [11]),
        .I1(\key_mem_reg[6]_6 [11]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [11]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [11]),
        .O(\block_w3_reg[11]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w3_reg[11]_i_8 
       (.I0(\dec_block/op158_in [0]),
        .I1(\dec_block/op161_in [0]),
        .I2(\block_w1_reg_reg[0] ),
        .I3(\block_w1_reg_reg[16] ),
        .O(\block_w3_reg[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[11]_i_8__0 
       (.I0(\key_mem_reg[3]_3 [11]),
        .I1(\key_mem_reg[2]_2 [11]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [11]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [11]),
        .O(\block_w3_reg[11]_i_8__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[11]_i_9 
       (.I0(\dec_block/op161_in [6]),
        .I1(\dec_block/op158_in [6]),
        .O(\block_w3_reg[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[11]_i_9__0 
       (.I0(\key_mem_reg[11]_11 [11]),
        .I1(\key_mem_reg[10]_10 [11]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [11]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [11]),
        .O(\block_w3_reg[11]_i_9__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[12]_i_10 
       (.I0(\dec_block/op159_in [1]),
        .I1(\dec_block/p_0_in46_in [2]),
        .O(\block_w3_reg[12]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w3_reg[12]_i_11 
       (.I0(\block_w1_reg[7]_i_4_n_0 ),
        .I1(round_key[75]),
        .I2(dec_new_block[75]),
        .I3(\dec_block/op161_in [4]),
        .O(\block_w3_reg[12]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[12]_i_12 
       (.I0(\dec_block/op159_in [4]),
        .I1(\dec_block/p_0_in46_in [5]),
        .O(\block_w3_reg[12]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \block_w3_reg[12]_i_13 
       (.I0(dec_new_block[67]),
        .I1(round_key[67]),
        .I2(\dec_block/op161_in [7]),
        .O(\block_w3_reg[12]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[12]_i_2__0 
       (.I0(\dec_block/op95_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[12] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[12]_i_3 
       (.I0(\block_w3_reg[12]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[12]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[12]_i_8_n_0 ),
        .O(round_key[12]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[12]_i_4__0 
       (.I0(\block_w3_reg[12]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[12]_i_7_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[12]_i_6__0_n_0 ),
        .I5(dec_new_block[12]),
        .O(\dec_block/op95_in [4]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[12]_i_5 
       (.I0(round_key[12]),
        .I1(core_block[12]),
        .O(addroundkey_return[11]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[12]_i_6 
       (.I0(\block_w3_reg[13]_i_10_n_0 ),
        .I1(\block_w3_reg[12]_i_9_n_0 ),
        .I2(\block_w3_reg[12]_i_10_n_0 ),
        .I3(\block_w3_reg[12]_i_11_n_0 ),
        .I4(\block_w3_reg[12]_i_12_n_0 ),
        .I5(\block_w3_reg[12]_i_13_n_0 ),
        .O(inv_mixcolumns_return0174_out__63[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[12]_i_6__0 
       (.I0(\block_w3_reg[12]_i_9__0_n_0 ),
        .I1(\key_mem_reg[14]_14 [12]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [12]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [12]),
        .O(\block_w3_reg[12]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[12]_i_7 
       (.I0(\key_mem_reg[7]_7 [12]),
        .I1(\key_mem_reg[6]_6 [12]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [12]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [12]),
        .O(\block_w3_reg[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[12]_i_8 
       (.I0(\key_mem_reg[3]_3 [12]),
        .I1(\key_mem_reg[2]_2 [12]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [12]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [12]),
        .O(\block_w3_reg[12]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[12]_i_9 
       (.I0(\dec_block/op158_in [5]),
        .I1(\dec_block/op161_in [5]),
        .I2(\dec_block/p_0_in46_in [6]),
        .I3(\dec_block/op159_in [5]),
        .I4(\dec_block/op161_in [1]),
        .I5(\block_w1_reg_reg[9] ),
        .O(\block_w3_reg[12]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[12]_i_9__0 
       (.I0(\key_mem_reg[11]_11 [12]),
        .I1(\key_mem_reg[10]_10 [12]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [12]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [12]),
        .O(\block_w3_reg[12]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[13]_i_10 
       (.I0(\dec_block/op159_in [6]),
        .I1(\dec_block/p_0_in46_in [7]),
        .I2(round_key[90]),
        .I3(dec_new_block[90]),
        .I4(\dec_block/op158_in [2]),
        .O(\block_w3_reg[13]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[13]_i_11 
       (.I0(\dec_block/op161_in [6]),
        .I1(\dec_block/op158_in [6]),
        .I2(round_key[82]),
        .I3(dec_new_block[82]),
        .I4(\dec_block/p_0_in46_in [3]),
        .O(\block_w3_reg[13]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[13]_i_12 
       (.I0(\dec_block/op158_in [4]),
        .I1(\dec_block/p_0_in46_in [5]),
        .O(\block_w3_reg[13]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[13]_i_13 
       (.I0(\dec_block/op159_in [5]),
        .I1(\dec_block/p_0_in46_in [6]),
        .O(\block_w3_reg[13]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[13]_i_14 
       (.I0(\dec_block/op159_in [7]),
        .I1(round_key[91]),
        .I2(dec_new_block[91]),
        .I3(\block_w1_reg[7]_i_4_n_0 ),
        .I4(round_key[75]),
        .I5(dec_new_block[75]),
        .O(\block_w3_reg[13]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[13]_i_2__0 
       (.I0(\dec_block/op95_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[13] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[13]_i_3 
       (.I0(\block_w3_reg[13]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[13]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[13]_i_7__0_n_0 ),
        .O(round_key[13]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[13]_i_4 
       (.I0(\block_w3_reg[13]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[13]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[13]_i_5__0_n_0 ),
        .I5(dec_new_block[13]),
        .O(\dec_block/op95_in [5]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[13]_i_5 
       (.I0(round_key[77]),
        .I1(core_block[77]),
        .O(p_0_out[35]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[13]_i_5__0 
       (.I0(\block_w3_reg[13]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [13]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [13]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [13]),
        .O(\block_w3_reg[13]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[13]_i_6 
       (.I0(\key_mem_reg[7]_7 [13]),
        .I1(\key_mem_reg[6]_6 [13]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [13]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [13]),
        .O(\block_w3_reg[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[13]_i_7 
       (.I0(\block_w3_reg[13]_i_10_n_0 ),
        .I1(\block_w3_reg[13]_i_11_n_0 ),
        .I2(\block_w3_reg[13]_i_12_n_0 ),
        .I3(\dec_block/op161_in [5]),
        .I4(\block_w3_reg[13]_i_13_n_0 ),
        .I5(\block_w3_reg[13]_i_14_n_0 ),
        .O(inv_mixcolumns_return0174_out__63[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[13]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [13]),
        .I1(\key_mem_reg[2]_2 [13]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [13]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [13]),
        .O(\block_w3_reg[13]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[13]_i_8 
       (.I0(\key_mem_reg[11]_11 [13]),
        .I1(\key_mem_reg[10]_10 [13]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [13]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [13]),
        .O(\block_w3_reg[13]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[14]_i_10 
       (.I0(\dec_block/op158_in [4]),
        .I1(\dec_block/op161_in [4]),
        .O(\block_w3_reg[14]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[14]_i_11 
       (.I0(\dec_block/op158_in [7]),
        .I1(round_key[83]),
        .I2(dec_new_block[83]),
        .I3(\block_w1_reg[7]_i_4_n_0 ),
        .I4(round_key[75]),
        .I5(dec_new_block[75]),
        .O(\block_w3_reg[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[14]_i_12 
       (.I0(\dec_block/op161_in [7]),
        .I1(round_key[67]),
        .I2(dec_new_block[67]),
        .I3(\dec_block/op159_in [7]),
        .I4(round_key[91]),
        .I5(dec_new_block[91]),
        .O(\block_w3_reg[14]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[14]_i_13 
       (.I0(\dec_block/p_0_in46_in [6]),
        .I1(\dec_block/op158_in [5]),
        .O(\block_w3_reg[14]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[14]_i_14 
       (.I0(\dec_block/op159_in [6]),
        .I1(\dec_block/p_0_in46_in [7]),
        .O(\block_w3_reg[14]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[14]_i_2__0 
       (.I0(\dec_block/op95_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[14] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[14]_i_3 
       (.I0(\block_w3_reg[14]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[14]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[14]_i_7__0_n_0 ),
        .O(round_key[14]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[14]_i_4 
       (.I0(\block_w3_reg[14]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[14]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[14]_i_5__0_n_0 ),
        .I5(dec_new_block[14]),
        .O(\dec_block/op95_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[14]_i_5 
       (.I0(round_key[78]),
        .I1(core_block[78]),
        .O(p_0_out[36]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[14]_i_5__0 
       (.I0(\block_w3_reg[14]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [14]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [14]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [14]),
        .O(\block_w3_reg[14]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[14]_i_6 
       (.I0(\key_mem_reg[7]_7 [14]),
        .I1(\key_mem_reg[6]_6 [14]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [14]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [14]),
        .O(\block_w3_reg[14]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[14]_i_7 
       (.I0(\block_w3_reg[14]_i_10_n_0 ),
        .I1(\block_w3_reg[14]_i_11_n_0 ),
        .I2(\block_w3_reg[14]_i_12_n_0 ),
        .I3(\block_w3_reg[14]_i_13_n_0 ),
        .I4(\block_w3_reg[14]_i_14_n_0 ),
        .I5(\dec_block/op161_in [6]),
        .O(inv_mixcolumns_return0174_out__63[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[14]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [14]),
        .I1(\key_mem_reg[2]_2 [14]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [14]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [14]),
        .O(\block_w3_reg[14]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[14]_i_8 
       (.I0(\key_mem_reg[11]_11 [14]),
        .I1(\key_mem_reg[10]_10 [14]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [14]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [14]),
        .O(\block_w3_reg[14]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[15]_i_11 
       (.I0(\dec_block/op159_in [4]),
        .I1(\dec_block/p_0_in46_in [5]),
        .I2(\dec_block/op158_in [4]),
        .I3(\dec_block/op161_in [4]),
        .I4(\dec_block/op161_in [7]),
        .I5(\dec_block/op159_in [7]),
        .O(\block_w3_reg[15]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[15]_i_12 
       (.I0(\dec_block/op161_in [5]),
        .I1(\dec_block/op158_in [5]),
        .O(\block_w3_reg[15]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[15]_i_2__0 
       (.I0(\dec_block/op95_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[15] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[15]_i_3 
       (.I0(\block_w3_reg[15]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[15]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[15]_i_7__0_n_0 ),
        .O(round_key[15]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[15]_i_4 
       (.I0(\block_w3_reg[15]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[15]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[15]_i_5__0_n_0 ),
        .I5(dec_new_block[15]),
        .O(\dec_block/op95_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[15]_i_5 
       (.I0(round_key[79]),
        .I1(core_block[79]),
        .O(p_0_out[37]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[15]_i_5__0 
       (.I0(\block_w3_reg[15]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [15]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [15]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [15]),
        .O(\block_w3_reg[15]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[15]_i_6 
       (.I0(\key_mem_reg[7]_7 [15]),
        .I1(\key_mem_reg[6]_6 [15]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [15]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [15]),
        .O(\block_w3_reg[15]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[15]_i_7 
       (.I0(\block_w3_reg[15]_i_11_n_0 ),
        .I1(\dec_block/op158_in [6]),
        .I2(\dec_block/p_0_in46_in [7]),
        .I3(\block_w1_reg[7]_i_4_n_0 ),
        .I4(\block_w3_reg[15]_i_12_n_0 ),
        .O(inv_mixcolumns_return0174_out__63[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[15]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [15]),
        .I1(\key_mem_reg[2]_2 [15]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [15]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [15]),
        .O(\block_w3_reg[15]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[15]_i_8 
       (.I0(\key_mem_reg[11]_11 [15]),
        .I1(\key_mem_reg[10]_10 [15]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [15]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [15]),
        .O(\block_w3_reg[15]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT3 #(
    .INIT(8'h60)) 
    \block_w3_reg[16]_i_2__0 
       (.I0(round_key[48]),
        .I1(core_block[48]),
        .I2(\block_w0_reg_reg[0]_1 ),
        .O(\block_reg_reg[2][16] ));
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \block_w3_reg[16]_i_3 
       (.I0(\block_w3_reg[16]_i_6_n_0 ),
        .I1(\block_w3_reg[16]_i_7_n_0 ),
        .I2(\block_w2_reg_reg[0] ),
        .I3(\block_w3_reg[16]_i_8_n_0 ),
        .I4(\block_w0_reg_reg[0]_1 ),
        .I5(\block_w0_reg_reg[16]_0 [2]),
        .O(\block_w2_reg_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[16]_i_3__0 
       (.I0(\block_w3_reg[16]_i_5_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w3_reg[16]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[16]_i_7__0_n_0 ),
        .O(round_key[16]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[16]_i_4 
       (.I0(\block_w3_reg[16]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[16]_i_6__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[16]_i_5_n_0 ),
        .I5(dec_new_block[16]),
        .O(\block_w3_reg_reg[16] ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[16]_i_5 
       (.I0(\block_w3_reg[16]_i_8__0_n_0 ),
        .I1(\key_mem_reg[14]_14 [16]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [16]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [16]),
        .O(\block_w3_reg[16]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[16]_i_6 
       (.I0(\dec_block/op126_in [7]),
        .I1(\dec_block/op127_in [7]),
        .O(\block_w3_reg[16]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[16]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [16]),
        .I1(\key_mem_reg[6]_6 [16]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [16]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [16]),
        .O(\block_w3_reg[16]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[16]_i_7 
       (.I0(\dec_block/op129_in [5]),
        .I1(\dec_block/op126_in [5]),
        .I2(\dec_block/p_0_in38_in [6]),
        .I3(\dec_block/op127_in [5]),
        .I4(\dec_block/op127_in [6]),
        .I5(\dec_block/p_0_in38_in [7]),
        .O(\block_w3_reg[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[16]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [16]),
        .I1(\key_mem_reg[2]_2 [16]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [16]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [16]),
        .O(\block_w3_reg[16]_i_7__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[16]_i_8 
       (.I0(\dec_block/op129_in [0]),
        .I1(\dec_block/op126_in [0]),
        .O(\block_w3_reg[16]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[16]_i_8__0 
       (.I0(\key_mem_reg[11]_11 [16]),
        .I1(\key_mem_reg[10]_10 [16]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [16]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [16]),
        .O(\block_w3_reg[16]_i_8__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[17]_i_2__0 
       (.I0(\dec_block/op96_in [1]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[17] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[17]_i_3 
       (.I0(\block_w3_reg[17]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[17]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[17]_i_8_n_0 ),
        .O(round_key[17]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[17]_i_4__0 
       (.I0(\block_w3_reg[17]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[17]_i_7_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[17]_i_6__0_n_0 ),
        .I5(dec_new_block[17]),
        .O(\dec_block/op96_in [1]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[17]_i_5 
       (.I0(round_key[17]),
        .I1(core_block[17]),
        .O(addroundkey_return[15]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[17]_i_6 
       (.I0(\block_w2_reg_reg[16] ),
        .I1(\dec_block/p_0_in38_in [2]),
        .I2(\block_w3_reg[20]_i_10_n_0 ),
        .I3(\block_w3_reg[22]_i_14_n_0 ),
        .I4(\dec_block/op126_in [0]),
        .I5(\block_w3_reg[17]_i_9_n_0 ),
        .O(inv_mixcolumns_return0149_out__55[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[17]_i_6__0 
       (.I0(\block_w3_reg[17]_i_9__0_n_0 ),
        .I1(\key_mem_reg[14]_14 [17]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [17]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [17]),
        .O(\block_w3_reg[17]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[17]_i_7 
       (.I0(\key_mem_reg[7]_7 [17]),
        .I1(\key_mem_reg[6]_6 [17]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [17]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [17]),
        .O(\block_w3_reg[17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[17]_i_8 
       (.I0(\key_mem_reg[3]_3 [17]),
        .I1(\key_mem_reg[2]_2 [17]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [17]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [17]),
        .O(\block_w3_reg[17]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[17]_i_9 
       (.I0(\block_w2_reg[7]_i_4_n_0 ),
        .I1(\dec_block/op126_in [7]),
        .O(\block_w3_reg[17]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[17]_i_9__0 
       (.I0(\key_mem_reg[11]_11 [17]),
        .I1(\key_mem_reg[10]_10 [17]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [17]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [17]),
        .O(\block_w3_reg[17]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[18]_i_10 
       (.I0(\dec_block/op126_in [7]),
        .I1(\dec_block/op129_in [7]),
        .O(\block_w3_reg[18]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[18]_i_3 
       (.I0(\block_w3_reg[18]_i_5_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w3_reg[18]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[18]_i_7_n_0 ),
        .O(round_key[18]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[18]_i_4 
       (.I0(round_key[50]),
        .I1(core_block[50]),
        .O(p_0_out[16]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[18]_i_5 
       (.I0(\block_w3_reg[18]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [18]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [18]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [18]),
        .O(\block_w3_reg[18]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[18]_i_6 
       (.I0(\block_w3_reg[18]_i_9_n_0 ),
        .I1(\dec_block/p_0_in38_in [3]),
        .I2(\dec_block/op127_in [1]),
        .I3(\block_w3_reg[18]_i_10_n_0 ),
        .I4(\block_w3_reg[21]_i_10_n_0 ),
        .I5(\block_w2_reg_reg[9] ),
        .O(inv_mixcolumns_return0149_out__55[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[18]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [18]),
        .I1(\key_mem_reg[6]_6 [18]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [18]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [18]),
        .O(\block_w3_reg[18]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[18]_i_7 
       (.I0(\key_mem_reg[3]_3 [18]),
        .I1(\key_mem_reg[2]_2 [18]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [18]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [18]),
        .O(\block_w3_reg[18]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[18]_i_8 
       (.I0(\key_mem_reg[11]_11 [18]),
        .I1(\key_mem_reg[10]_10 [18]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [18]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [18]),
        .O(\block_w3_reg[18]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w3_reg[18]_i_9 
       (.I0(\block_w2_reg_reg[16] ),
        .I1(\block_w2_reg_reg[0] ),
        .I2(\dec_block/op126_in [6]),
        .I3(\dec_block/op129_in [6]),
        .O(\block_w3_reg[18]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[19]_i_10 
       (.I0(\dec_block/op127_in [2]),
        .I1(dec_new_block[43]),
        .I2(round_key[43]),
        .I3(\block_w2_reg[7]_i_4_n_0 ),
        .I4(\dec_block/op129_in [3]),
        .I5(\dec_block/op126_in [2]),
        .O(\block_w3_reg[19]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[19]_i_10__0 
       (.I0(\key_mem_reg[11]_11 [19]),
        .I1(\key_mem_reg[10]_10 [19]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [19]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [19]),
        .O(\block_w3_reg[19]_i_10__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \block_w3_reg[19]_i_11 
       (.I0(dec_new_block[35]),
        .I1(round_key[35]),
        .I2(\dec_block/op129_in [7]),
        .O(\block_w3_reg[19]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[19]_i_12 
       (.I0(\block_w2_reg[18]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[18]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[18]_i_6__0_n_0 ),
        .I5(dec_new_block[50]),
        .O(\dec_block/op127_in [2]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[19]_i_13 
       (.I0(\block_w2_reg[27]_i_10_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w2_reg[27]_i_9_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w2_reg[27]_i_7_n_0 ),
        .I5(dec_new_block[59]),
        .O(\dec_block/op129_in [3]));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[19]_i_2__0 
       (.I0(\dec_block/op96_in [3]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[19] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[19]_i_3 
       (.I0(\block_w3_reg[19]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w3_reg[19]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[19]_i_8_n_0 ),
        .O(round_key[19]));
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[19]_i_4__0 
       (.I0(round_key[19]),
        .I1(dec_new_block[19]),
        .O(\dec_block/op96_in [3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[19]_i_5 
       (.I0(round_key[19]),
        .I1(core_block[19]),
        .O(addroundkey_return[17]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[19]_i_6 
       (.I0(\block_w3_reg[16]_i_7_n_0 ),
        .I1(\block_w3_reg[19]_i_9_n_0 ),
        .I2(\block_w3_reg[19]_i_10_n_0 ),
        .I3(\block_w3_reg[20]_i_11_n_0 ),
        .I4(\block_w3_reg[19]_i_11_n_0 ),
        .O(inv_mixcolumns_return0149_out__55[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[19]_i_6__0 
       (.I0(\block_w3_reg[19]_i_10__0_n_0 ),
        .I1(\key_mem_reg[14]_14 [19]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [19]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [19]),
        .O(\block_w3_reg[19]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[19]_i_7 
       (.I0(\key_mem_reg[7]_7 [19]),
        .I1(\key_mem_reg[6]_6 [19]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [19]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [19]),
        .O(\block_w3_reg[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[19]_i_8 
       (.I0(\key_mem_reg[3]_3 [19]),
        .I1(\key_mem_reg[2]_2 [19]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [19]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [19]),
        .O(\block_w3_reg[19]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w3_reg[19]_i_9 
       (.I0(\block_w2_reg_reg[16] ),
        .I1(\block_w2_reg_reg[0] ),
        .I2(\dec_block/op126_in [0]),
        .I3(\dec_block/op129_in [0]),
        .O(\block_w3_reg[19]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[1]_i_2__0 
       (.I0(\dec_block/p_0_in31_in [2]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[1] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[1]_i_3 
       (.I0(\block_w3_reg[1]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[1]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[1]_i_8_n_0 ),
        .O(round_key[1]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[1]_i_4__0 
       (.I0(\block_w3_reg[1]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[1]_i_7_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[1]_i_6__0_n_0 ),
        .I5(dec_new_block[1]),
        .O(\dec_block/p_0_in31_in [2]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[1]_i_5 
       (.I0(round_key[1]),
        .I1(core_block[1]),
        .O(addroundkey_return[0]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[1]_i_6 
       (.I0(\dec_block/op193_in [0]),
        .I1(\dec_block/op191_in [1]),
        .I2(\block_w3_reg[4]_i_10_n_0 ),
        .I3(\block_w3_reg[6]_i_14_n_0 ),
        .I4(\block_w0_reg_reg[0] ),
        .I5(\block_w3_reg[1]_i_9_n_0 ),
        .O(inv_mixcolumns_return0198_out__63[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[1]_i_6__0 
       (.I0(\block_w3_reg[1]_i_9__0_n_0 ),
        .I1(\key_mem_reg[14]_14 [1]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [1]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [1]),
        .O(\block_w3_reg[1]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[1]_i_7 
       (.I0(\key_mem_reg[7]_7 [1]),
        .I1(\key_mem_reg[6]_6 [1]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [1]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [1]),
        .O(\block_w3_reg[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[1]_i_8 
       (.I0(\key_mem_reg[3]_3 [1]),
        .I1(\key_mem_reg[2]_2 [1]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [1]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [1]),
        .O(\block_w3_reg[1]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[1]_i_9 
       (.I0(\dec_block/op191_in [7]),
        .I1(\dec_block/op193_in [7]),
        .O(\block_w3_reg[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[1]_i_9__0 
       (.I0(\key_mem_reg[11]_11 [1]),
        .I1(\key_mem_reg[10]_10 [1]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [1]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [1]),
        .O(\block_w3_reg[1]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[20]_i_10 
       (.I0(\dec_block/op127_in [5]),
        .I1(\dec_block/p_0_in38_in [6]),
        .I2(\dec_block/op126_in [5]),
        .I3(\dec_block/op129_in [5]),
        .I4(\dec_block/op129_in [1]),
        .I5(\block_w2_reg_reg[9] ),
        .O(\block_w3_reg[20]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[20]_i_10__0 
       (.I0(\key_mem_reg[11]_11 [20]),
        .I1(\key_mem_reg[10]_10 [20]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [20]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [20]),
        .O(\block_w3_reg[20]_i_10__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[20]_i_11 
       (.I0(\dec_block/p_0_in38_in [2]),
        .I1(\dec_block/op127_in [1]),
        .O(\block_w3_reg[20]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[20]_i_2__0 
       (.I0(\dec_block/op96_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[20] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[20]_i_3 
       (.I0(\block_w3_reg[20]_i_7_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[20]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[20]_i_9__0_n_0 ),
        .O(round_key[20]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[20]_i_4 
       (.I0(\block_w3_reg[20]_i_9__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[20]_i_8_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[20]_i_7_n_0 ),
        .I5(dec_new_block[20]),
        .O(\dec_block/op96_in [4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[20]_i_6 
       (.I0(\block_w3_reg[20]_i_9_n_0 ),
        .I1(\dec_block/p_0_in38_in [5]),
        .I2(\block_w3_reg[20]_i_10_n_0 ),
        .I3(\block_w3_reg[20]_i_11_n_0 ),
        .I4(\block_w3_reg[21]_i_11_n_0 ),
        .I5(\block_w3_reg[22]_i_11_n_0 ),
        .O(inv_mixcolumns_return0149_out__55[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[20]_i_6__0 
       (.I0(round_key[20]),
        .I1(core_block[20]),
        .O(addroundkey_return[18]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[20]_i_7 
       (.I0(\block_w3_reg[20]_i_10__0_n_0 ),
        .I1(\key_mem_reg[14]_14 [20]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [20]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [20]),
        .O(\block_w3_reg[20]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[20]_i_8 
       (.I0(\key_mem_reg[7]_7 [20]),
        .I1(\key_mem_reg[6]_6 [20]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [20]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [20]),
        .O(\block_w3_reg[20]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[20]_i_9 
       (.I0(\dec_block/op126_in [4]),
        .I1(\dec_block/op129_in [4]),
        .O(\block_w3_reg[20]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[20]_i_9__0 
       (.I0(\key_mem_reg[3]_3 [20]),
        .I1(\key_mem_reg[2]_2 [20]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [20]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [20]),
        .O(\block_w3_reg[20]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[21]_i_10 
       (.I0(\dec_block/p_0_in38_in [7]),
        .I1(\dec_block/op127_in [6]),
        .I2(round_key[58]),
        .I3(dec_new_block[58]),
        .I4(\dec_block/op126_in [2]),
        .O(\block_w3_reg[21]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[21]_i_11 
       (.I0(\dec_block/op129_in [6]),
        .I1(\dec_block/op126_in [6]),
        .I2(round_key[50]),
        .I3(dec_new_block[50]),
        .I4(\dec_block/p_0_in38_in [3]),
        .O(\block_w3_reg[21]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[21]_i_12 
       (.I0(\dec_block/op126_in [4]),
        .I1(\dec_block/op127_in [4]),
        .O(\block_w3_reg[21]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[21]_i_13 
       (.I0(\dec_block/op129_in [5]),
        .I1(\dec_block/op126_in [5]),
        .O(\block_w3_reg[21]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[21]_i_14 
       (.I0(\dec_block/op129_in [7]),
        .I1(round_key[35]),
        .I2(dec_new_block[35]),
        .I3(\dec_block/op126_in [7]),
        .I4(round_key[51]),
        .I5(dec_new_block[51]),
        .O(\block_w3_reg[21]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[21]_i_2__0 
       (.I0(\dec_block/op96_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[21] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[21]_i_3 
       (.I0(\block_w3_reg[21]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[21]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[21]_i_7__0_n_0 ),
        .O(round_key[21]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[21]_i_4 
       (.I0(\block_w3_reg[21]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[21]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[21]_i_5__0_n_0 ),
        .I5(dec_new_block[21]),
        .O(\dec_block/op96_in [5]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[21]_i_5 
       (.I0(round_key[53]),
        .I1(core_block[53]),
        .O(p_0_out[19]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[21]_i_5__0 
       (.I0(\block_w3_reg[21]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [21]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [21]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [21]),
        .O(\block_w3_reg[21]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[21]_i_6 
       (.I0(\key_mem_reg[7]_7 [21]),
        .I1(\key_mem_reg[6]_6 [21]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [21]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [21]),
        .O(\block_w3_reg[21]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[21]_i_7 
       (.I0(\block_w3_reg[21]_i_10_n_0 ),
        .I1(\block_w3_reg[21]_i_11_n_0 ),
        .I2(\block_w3_reg[21]_i_12_n_0 ),
        .I3(\dec_block/p_0_in38_in [6]),
        .I4(\block_w3_reg[21]_i_13_n_0 ),
        .I5(\block_w3_reg[21]_i_14_n_0 ),
        .O(inv_mixcolumns_return0149_out__55[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[21]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [21]),
        .I1(\key_mem_reg[2]_2 [21]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [21]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [21]),
        .O(\block_w3_reg[21]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[21]_i_8 
       (.I0(\key_mem_reg[11]_11 [21]),
        .I1(\key_mem_reg[10]_10 [21]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [21]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [21]),
        .O(\block_w3_reg[21]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[22]_i_10 
       (.I0(\dec_block/p_0_in38_in [5]),
        .I1(\dec_block/op127_in [4]),
        .O(\block_w3_reg[22]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[22]_i_11 
       (.I0(\dec_block/op126_in [7]),
        .I1(round_key[51]),
        .I2(dec_new_block[51]),
        .I3(\block_w2_reg[7]_i_4_n_0 ),
        .I4(round_key[43]),
        .I5(dec_new_block[43]),
        .O(\block_w3_reg[22]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[22]_i_12 
       (.I0(\dec_block/op129_in [7]),
        .I1(round_key[35]),
        .I2(dec_new_block[35]),
        .I3(\dec_block/op127_in [7]),
        .I4(round_key[59]),
        .I5(dec_new_block[59]),
        .O(\block_w3_reg[22]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[22]_i_13 
       (.I0(\dec_block/op126_in [5]),
        .I1(\dec_block/op127_in [5]),
        .O(\block_w3_reg[22]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[22]_i_14 
       (.I0(\dec_block/op129_in [6]),
        .I1(\dec_block/op126_in [6]),
        .O(\block_w3_reg[22]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[22]_i_2__0 
       (.I0(\dec_block/op96_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[22] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[22]_i_3 
       (.I0(\block_w3_reg[22]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[22]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[22]_i_7__0_n_0 ),
        .O(round_key[22]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[22]_i_4 
       (.I0(\block_w3_reg[22]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[22]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[22]_i_5__0_n_0 ),
        .I5(dec_new_block[22]),
        .O(\dec_block/op96_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[22]_i_5 
       (.I0(round_key[54]),
        .I1(core_block[54]),
        .O(p_0_out[20]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[22]_i_5__0 
       (.I0(\block_w3_reg[22]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [22]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [22]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [22]),
        .O(\block_w3_reg[22]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[22]_i_6 
       (.I0(\key_mem_reg[7]_7 [22]),
        .I1(\key_mem_reg[6]_6 [22]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [22]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [22]),
        .O(\block_w3_reg[22]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[22]_i_7 
       (.I0(\block_w3_reg[22]_i_10_n_0 ),
        .I1(\block_w3_reg[22]_i_11_n_0 ),
        .I2(\block_w3_reg[22]_i_12_n_0 ),
        .I3(\block_w3_reg[22]_i_13_n_0 ),
        .I4(\block_w3_reg[22]_i_14_n_0 ),
        .I5(\dec_block/p_0_in38_in [7]),
        .O(inv_mixcolumns_return0149_out__55[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[22]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [22]),
        .I1(\key_mem_reg[2]_2 [22]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [22]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [22]),
        .O(\block_w3_reg[22]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[22]_i_8 
       (.I0(\key_mem_reg[11]_11 [22]),
        .I1(\key_mem_reg[10]_10 [22]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [22]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [22]),
        .O(\block_w3_reg[22]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[23]_i_11 
       (.I0(\dec_block/p_0_in38_in [5]),
        .I1(\dec_block/op127_in [4]),
        .I2(\dec_block/op126_in [4]),
        .I3(\dec_block/op129_in [4]),
        .I4(\dec_block/op126_in [7]),
        .I5(\block_w2_reg[7]_i_4_n_0 ),
        .O(\block_w3_reg[23]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[23]_i_12 
       (.I0(\dec_block/p_0_in38_in [6]),
        .I1(\dec_block/op127_in [5]),
        .O(\block_w3_reg[23]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[23]_i_2__0 
       (.I0(\dec_block/op96_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[23] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[23]_i_3 
       (.I0(\block_w3_reg[23]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[23]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[23]_i_7__0_n_0 ),
        .O(round_key[23]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[23]_i_4 
       (.I0(\block_w3_reg[23]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[23]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[23]_i_5__0_n_0 ),
        .I5(dec_new_block[23]),
        .O(\dec_block/op96_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[23]_i_5 
       (.I0(round_key[55]),
        .I1(core_block[55]),
        .O(p_0_out[21]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[23]_i_5__0 
       (.I0(\block_w3_reg[23]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [23]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [23]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [23]),
        .O(\block_w3_reg[23]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[23]_i_6 
       (.I0(\key_mem_reg[7]_7 [23]),
        .I1(\key_mem_reg[6]_6 [23]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [23]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [23]),
        .O(\block_w3_reg[23]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[23]_i_7 
       (.I0(\block_w3_reg[23]_i_11_n_0 ),
        .I1(\dec_block/op126_in [6]),
        .I2(\dec_block/op127_in [6]),
        .I3(\dec_block/op129_in [7]),
        .I4(\block_w3_reg[23]_i_12_n_0 ),
        .O(inv_mixcolumns_return0149_out__55[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[23]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [23]),
        .I1(\key_mem_reg[2]_2 [23]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [23]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [23]),
        .O(\block_w3_reg[23]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[23]_i_8 
       (.I0(\key_mem_reg[11]_11 [23]),
        .I1(\key_mem_reg[10]_10 [23]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [23]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [23]),
        .O(\block_w3_reg[23]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w3_reg[24]_i_10 
       (.I0(\dec_block/p_0_in31_in [6]),
        .I1(\dec_block/op96_in [5]),
        .I2(\dec_block/op98_in [5]),
        .I3(\dec_block/op95_in [5]),
        .O(\block_w3_reg[24]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[24]_i_11 
       (.I0(\dec_block/op96_in [7]),
        .I1(\dec_block/op98_in [7]),
        .O(\block_w3_reg[24]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[24]_i_12 
       (.I0(\block_w3_reg_reg[16] ),
        .I1(\block_w3_reg_reg[0] ),
        .O(\block_w3_reg[24]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[24]_i_13 
       (.I0(\dec_block/op95_in [6]),
        .I1(\dec_block/op98_in [6]),
        .O(\block_w3_reg[24]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[24]_i_2__0 
       (.I0(\dec_block/op98_in [0]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[24] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[24]_i_3 
       (.I0(\block_w3_reg[24]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[24]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[24]_i_7__0_n_0 ),
        .O(round_key[24]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[24]_i_4 
       (.I0(\block_w3_reg[24]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[24]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[24]_i_5__0_n_0 ),
        .I5(dec_new_block[24]),
        .O(\dec_block/op98_in [0]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[24]_i_5 
       (.I0(round_key[24]),
        .I1(core_block[24]),
        .O(p_0_out[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[24]_i_5__0 
       (.I0(\block_w3_reg[24]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [24]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [24]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [24]),
        .O(\block_w3_reg[24]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[24]_i_6 
       (.I0(\key_mem_reg[7]_7 [24]),
        .I1(\key_mem_reg[6]_6 [24]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [24]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [24]),
        .O(\block_w3_reg[24]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[24]_i_7 
       (.I0(\block_w3_reg[24]_i_10_n_0 ),
        .I1(\dec_block/op95_in [0]),
        .I2(\block_w3_reg[24]_i_11_n_0 ),
        .I3(\block_w3_reg[24]_i_12_n_0 ),
        .I4(\block_w3_reg[24]_i_13_n_0 ),
        .O(inv_mixcolumns_return0124_out__47[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[24]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [24]),
        .I1(\key_mem_reg[2]_2 [24]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [24]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [24]),
        .O(\block_w3_reg[24]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[24]_i_8 
       (.I0(\key_mem_reg[11]_11 [24]),
        .I1(\key_mem_reg[10]_10 [24]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [24]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [24]),
        .O(\block_w3_reg[24]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[25]_i_10 
       (.I0(\key_mem_reg[3]_3 [25]),
        .I1(\key_mem_reg[2]_2 [25]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [25]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [25]),
        .O(\block_w3_reg[25]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[25]_i_11 
       (.I0(\key_mem_reg[11]_11 [25]),
        .I1(\key_mem_reg[10]_10 [25]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [25]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [25]),
        .O(\block_w3_reg[25]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[25]_i_2__0 
       (.I0(\dec_block/op98_in [1]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[25] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[25]_i_3 
       (.I0(\block_w3_reg[25]_i_7_n_0 ),
        .I1(muxed_round_nr[3]),
        .I2(\block_w3_reg[25]_i_9__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[25]_i_10_n_0 ),
        .O(round_key[25]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[25]_i_4 
       (.I0(\block_w3_reg[25]_i_10_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[25]_i_9__0_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[25]_i_7_n_0 ),
        .I5(dec_new_block[25]),
        .O(\dec_block/op98_in [1]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[25]_i_6 
       (.I0(\block_w1_reg[9]_i_6__0_n_0 ),
        .I1(\block_w3_reg[30]_i_14_n_0 ),
        .I2(\dec_block/op98_in [0]),
        .I3(\block_w0_reg[16]_i_5_n_0 ),
        .I4(\block_w3_reg[25]_i_9_n_0 ),
        .I5(\block_w3_reg_reg[16] ),
        .O(inv_mixcolumns_return0124_out__47[1]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[25]_i_6__0 
       (.I0(round_key[25]),
        .I1(core_block[25]),
        .O(p_0_out[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[25]_i_7 
       (.I0(\block_w3_reg[25]_i_11_n_0 ),
        .I1(\key_mem_reg[14]_14 [25]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [25]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [25]),
        .O(\block_w3_reg[25]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[25]_i_9 
       (.I0(\dec_block/op95_in [1]),
        .I1(\dec_block/op95_in [5]),
        .I2(\dec_block/op98_in [5]),
        .I3(\dec_block/op96_in [5]),
        .I4(\dec_block/p_0_in31_in [6]),
        .O(\block_w3_reg[25]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[25]_i_9__0 
       (.I0(\key_mem_reg[7]_7 [25]),
        .I1(\key_mem_reg[6]_6 [25]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [25]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [25]),
        .O(\block_w3_reg[25]_i_9__0_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[26]_i_3 
       (.I0(\block_w3_reg[26]_i_5_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w3_reg[26]_i_6__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[26]_i_7_n_0 ),
        .O(round_key[26]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[26]_i_4 
       (.I0(round_key[26]),
        .I1(core_block[26]),
        .O(p_0_out[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[26]_i_5 
       (.I0(\block_w3_reg[26]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [26]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [26]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [26]),
        .O(\block_w3_reg[26]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[26]_i_6 
       (.I0(\block_w2_reg[0]_i_6_n_0 ),
        .I1(\block_w3_reg[26]_i_9_n_0 ),
        .I2(\dec_block/op96_in [7]),
        .I3(\block_w3_reg[30]_i_14_n_0 ),
        .I4(\block_w3_reg[29]_i_11_n_0 ),
        .I5(\dec_block/op98_in [1]),
        .O(inv_mixcolumns_return0124_out__47[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[26]_i_6__0 
       (.I0(\key_mem_reg[7]_7 [26]),
        .I1(\key_mem_reg[6]_6 [26]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [26]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [26]),
        .O(\block_w3_reg[26]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[26]_i_7 
       (.I0(\key_mem_reg[3]_3 [26]),
        .I1(\key_mem_reg[2]_2 [26]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [26]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [26]),
        .O(\block_w3_reg[26]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[26]_i_8 
       (.I0(\key_mem_reg[11]_11 [26]),
        .I1(\key_mem_reg[10]_10 [26]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [26]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [26]),
        .O(\block_w3_reg[26]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[26]_i_9 
       (.I0(\dec_block/op95_in [2]),
        .I1(\dec_block/op96_in [1]),
        .O(\block_w3_reg[26]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w3_reg[27]_i_10 
       (.I0(dec_new_block[18]),
        .I1(round_key[18]),
        .I2(\dec_block/op98_in [6]),
        .I3(\dec_block/op95_in [6]),
        .O(\block_w3_reg[27]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[27]_i_10__0 
       (.I0(\key_mem_reg[11]_11 [27]),
        .I1(\key_mem_reg[10]_10 [27]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [27]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [27]),
        .O(\block_w3_reg[27]_i_10__0_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[27]_i_3 
       (.I0(\block_w3_reg[27]_i_6_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[27]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[27]_i_8__0_n_0 ),
        .O(round_key[27]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[27]_i_5 
       (.I0(\block_w3_reg[30]_i_11_n_0 ),
        .I1(\block_w3_reg[27]_i_8_n_0 ),
        .I2(\dec_block/op98_in [2]),
        .I3(\dec_block/p_0_in31_in [4]),
        .I4(\block_w3_reg[28]_i_9_n_0 ),
        .I5(\block_w3_reg[27]_i_10_n_0 ),
        .O(inv_mixcolumns_return0124_out__47[3]));
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[27]_i_5__0 
       (.I0(round_key[27]),
        .I1(core_block[27]),
        .O(p_0_out[3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[27]_i_6 
       (.I0(\block_w3_reg[27]_i_10__0_n_0 ),
        .I1(\key_mem_reg[14]_14 [27]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [27]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [27]),
        .O(\block_w3_reg[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[27]_i_7 
       (.I0(\key_mem_reg[7]_7 [27]),
        .I1(\key_mem_reg[6]_6 [27]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [27]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [27]),
        .O(\block_w3_reg[27]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w3_reg[27]_i_8 
       (.I0(\block_w3_reg_reg[0] ),
        .I1(\block_w3_reg_reg[16] ),
        .I2(\dec_block/op98_in [0]),
        .I3(\dec_block/op95_in [0]),
        .O(\block_w3_reg[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[27]_i_8__0 
       (.I0(\key_mem_reg[3]_3 [27]),
        .I1(\key_mem_reg[2]_2 [27]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [27]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [27]),
        .O(\block_w3_reg[27]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[27]_i_9 
       (.I0(\block_w3_reg[26]_i_7_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[26]_i_6__0_n_0 ),
        .I3(muxed_round_nr[3]),
        .I4(\block_w3_reg[26]_i_5_n_0 ),
        .I5(dec_new_block[26]),
        .O(\dec_block/op98_in [2]));
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w3_reg[28]_i_10 
       (.I0(\dec_block/op95_in [7]),
        .I1(round_key[19]),
        .I2(dec_new_block[19]),
        .I3(\dec_block/op95_in [4]),
        .O(\block_w3_reg[28]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[28]_i_10__0 
       (.I0(\key_mem_reg[11]_11 [28]),
        .I1(\key_mem_reg[10]_10 [28]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [28]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [28]),
        .O(\block_w3_reg[28]_i_10__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[28]_i_11 
       (.I0(\dec_block/op96_in [4]),
        .I1(\dec_block/p_0_in31_in [5]),
        .O(\block_w3_reg[28]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \block_w3_reg[28]_i_12 
       (.I0(dec_new_block[27]),
        .I1(round_key[27]),
        .I2(\dec_block/op96_in [7]),
        .O(\block_w3_reg[28]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[28]_i_2__0 
       (.I0(\dec_block/op98_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[28] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[28]_i_3 
       (.I0(\block_w3_reg[28]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[28]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[28]_i_8_n_0 ),
        .O(round_key[28]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[28]_i_4__0 
       (.I0(\block_w3_reg[28]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[28]_i_7_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w3_reg[28]_i_6__0_n_0 ),
        .I5(dec_new_block[28]),
        .O(\dec_block/op98_in [4]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[28]_i_5 
       (.I0(round_key[28]),
        .I1(core_block[28]),
        .O(p_0_out[4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[28]_i_6 
       (.I0(\block_w3_reg[29]_i_10_n_0 ),
        .I1(\block_w3_reg[28]_i_9_n_0 ),
        .I2(\block_w1_reg[9]_i_6__0_n_0 ),
        .I3(\block_w3_reg[28]_i_10_n_0 ),
        .I4(\block_w3_reg[28]_i_11_n_0 ),
        .I5(\block_w3_reg[28]_i_12_n_0 ),
        .O(inv_mixcolumns_return0124_out__47[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[28]_i_6__0 
       (.I0(\block_w3_reg[28]_i_10__0_n_0 ),
        .I1(\key_mem_reg[14]_14 [28]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [28]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [28]),
        .O(\block_w3_reg[28]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[28]_i_7 
       (.I0(\key_mem_reg[7]_7 [28]),
        .I1(\key_mem_reg[6]_6 [28]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [28]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [28]),
        .O(\block_w3_reg[28]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[28]_i_8 
       (.I0(\key_mem_reg[3]_3 [28]),
        .I1(\key_mem_reg[2]_2 [28]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [28]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [28]),
        .O(\block_w3_reg[28]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[28]_i_9 
       (.I0(\dec_block/p_0_in31_in [6]),
        .I1(\dec_block/op96_in [5]),
        .I2(\dec_block/op98_in [5]),
        .I3(\dec_block/op95_in [5]),
        .I4(\dec_block/op95_in [1]),
        .I5(\dec_block/op98_in [1]),
        .O(\block_w3_reg[28]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[29]_i_10 
       (.I0(\dec_block/op96_in [6]),
        .I1(\dec_block/p_0_in31_in [7]),
        .I2(round_key[26]),
        .I3(dec_new_block[26]),
        .I4(\dec_block/op95_in [2]),
        .O(\block_w3_reg[29]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[29]_i_11 
       (.I0(\dec_block/op95_in [6]),
        .I1(\dec_block/op98_in [6]),
        .I2(round_key[18]),
        .I3(dec_new_block[18]),
        .I4(\dec_block/p_0_in31_in [3]),
        .O(\block_w3_reg[29]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[29]_i_12 
       (.I0(\dec_block/op96_in [4]),
        .I1(\dec_block/op98_in [4]),
        .O(\block_w3_reg[29]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[29]_i_13 
       (.I0(\dec_block/op96_in [5]),
        .I1(\dec_block/p_0_in31_in [6]),
        .O(\block_w3_reg[29]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[29]_i_14 
       (.I0(\dec_block/op96_in [7]),
        .I1(round_key[27]),
        .I2(dec_new_block[27]),
        .I3(\block_w3_reg[7]_i_4_n_0 ),
        .I4(round_key[11]),
        .I5(dec_new_block[11]),
        .O(\block_w3_reg[29]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[29]_i_2__0 
       (.I0(\dec_block/op98_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[29] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[29]_i_3 
       (.I0(\block_w3_reg[29]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[29]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[29]_i_7__0_n_0 ),
        .O(round_key[29]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[29]_i_4 
       (.I0(\block_w3_reg[29]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[29]_i_6_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w3_reg[29]_i_5__0_n_0 ),
        .I5(dec_new_block[29]),
        .O(\dec_block/op98_in [5]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[29]_i_5 
       (.I0(round_key[29]),
        .I1(core_block[29]),
        .O(p_0_out[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[29]_i_5__0 
       (.I0(\block_w3_reg[29]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [29]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [29]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [29]),
        .O(\block_w3_reg[29]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[29]_i_6 
       (.I0(\key_mem_reg[7]_7 [29]),
        .I1(\key_mem_reg[6]_6 [29]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [29]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [29]),
        .O(\block_w3_reg[29]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[29]_i_7 
       (.I0(\block_w3_reg[29]_i_10_n_0 ),
        .I1(\block_w3_reg[29]_i_11_n_0 ),
        .I2(\block_w3_reg[29]_i_12_n_0 ),
        .I3(\dec_block/op95_in [5]),
        .I4(\block_w3_reg[29]_i_13_n_0 ),
        .I5(\block_w3_reg[29]_i_14_n_0 ),
        .O(inv_mixcolumns_return0124_out__47[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[29]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [29]),
        .I1(\key_mem_reg[2]_2 [29]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [29]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [29]),
        .O(\block_w3_reg[29]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[29]_i_8 
       (.I0(\key_mem_reg[11]_11 [29]),
        .I1(\key_mem_reg[10]_10 [29]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [29]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [29]),
        .O(\block_w3_reg[29]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[2]_i_10 
       (.I0(\dec_block/op190_in [7]),
        .I1(\dec_block/op193_in [7]),
        .O(\block_w3_reg[2]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[2]_i_11 
       (.I0(\block_w0_reg_reg[16] ),
        .I1(\block_w0_reg_reg[0] ),
        .O(\block_w3_reg[2]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w3_reg[2]_i_12 
       (.I0(dec_new_block[114]),
        .I1(round_key[114]),
        .I2(\dec_block/op193_in [6]),
        .I3(\dec_block/op190_in [6]),
        .O(\block_w3_reg[2]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[2]_i_2__0 
       (.I0(\dec_block/p_0_in31_in [3]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[2] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[2]_i_3 
       (.I0(\block_w3_reg[2]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[2]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[2]_i_7__0_n_0 ),
        .O(round_key[2]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[2]_i_4 
       (.I0(\block_w3_reg[2]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[2]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[2]_i_5__0_n_0 ),
        .I5(dec_new_block[2]),
        .O(\dec_block/p_0_in31_in [3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[2]_i_5 
       (.I0(round_key[98]),
        .I1(core_block[98]),
        .O(p_0_out[47]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[2]_i_5__0 
       (.I0(\block_w3_reg[2]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [2]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [2]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [2]),
        .O(\block_w3_reg[2]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[2]_i_6 
       (.I0(\key_mem_reg[7]_7 [2]),
        .I1(\key_mem_reg[6]_6 [2]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [2]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [2]),
        .O(\block_w3_reg[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[2]_i_7 
       (.I0(\block_w3_reg[5]_i_10_n_0 ),
        .I1(\dec_block/p_0_in54_in [2]),
        .I2(\dec_block/op193_in [1]),
        .I3(\block_w3_reg[2]_i_10_n_0 ),
        .I4(\block_w3_reg[2]_i_11_n_0 ),
        .I5(\block_w3_reg[2]_i_12_n_0 ),
        .O(inv_mixcolumns_return0198_out__63[1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[2]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [2]),
        .I1(\key_mem_reg[2]_2 [2]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [2]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [2]),
        .O(\block_w3_reg[2]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[2]_i_8 
       (.I0(\key_mem_reg[11]_11 [2]),
        .I1(\key_mem_reg[10]_10 [2]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [2]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [2]),
        .O(\block_w3_reg[2]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[30]_i_10 
       (.I0(\dec_block/op95_in [4]),
        .I1(\dec_block/op98_in [4]),
        .O(\block_w3_reg[30]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[30]_i_11 
       (.I0(\block_w3_reg[7]_i_4_n_0 ),
        .I1(round_key[11]),
        .I2(dec_new_block[11]),
        .I3(\dec_block/op95_in [7]),
        .I4(round_key[19]),
        .I5(dec_new_block[19]),
        .O(\block_w3_reg[30]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[30]_i_12 
       (.I0(\dec_block/op98_in [7]),
        .I1(round_key[3]),
        .I2(dec_new_block[3]),
        .I3(\dec_block/op96_in [7]),
        .I4(round_key[27]),
        .I5(dec_new_block[27]),
        .O(\block_w3_reg[30]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[30]_i_13 
       (.I0(\dec_block/op96_in [5]),
        .I1(\dec_block/op98_in [5]),
        .O(\block_w3_reg[30]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[30]_i_14 
       (.I0(\dec_block/op96_in [6]),
        .I1(\dec_block/p_0_in31_in [7]),
        .O(\block_w3_reg[30]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[30]_i_2__0 
       (.I0(\dec_block/op98_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[30] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[30]_i_3 
       (.I0(\block_w3_reg[30]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[30]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[30]_i_7__0_n_0 ),
        .O(round_key[30]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[30]_i_4 
       (.I0(\block_w3_reg[30]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[30]_i_6_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w3_reg[30]_i_5__0_n_0 ),
        .I5(dec_new_block[30]),
        .O(\dec_block/op98_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[30]_i_5 
       (.I0(round_key[30]),
        .I1(core_block[30]),
        .O(p_0_out[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[30]_i_5__0 
       (.I0(\block_w3_reg[30]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [30]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [30]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [30]),
        .O(\block_w3_reg[30]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[30]_i_6 
       (.I0(\key_mem_reg[7]_7 [30]),
        .I1(\key_mem_reg[6]_6 [30]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [30]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [30]),
        .O(\block_w3_reg[30]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[30]_i_7 
       (.I0(\block_w3_reg[30]_i_10_n_0 ),
        .I1(\block_w3_reg[30]_i_11_n_0 ),
        .I2(\block_w3_reg[30]_i_12_n_0 ),
        .I3(\block_w3_reg[30]_i_13_n_0 ),
        .I4(\block_w3_reg[30]_i_14_n_0 ),
        .I5(\dec_block/op95_in [6]),
        .O(inv_mixcolumns_return0124_out__47[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[30]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [30]),
        .I1(\key_mem_reg[2]_2 [30]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [30]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [30]),
        .O(\block_w3_reg[30]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[30]_i_8 
       (.I0(\key_mem_reg[11]_11 [30]),
        .I1(\key_mem_reg[10]_10 [30]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [30]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [30]),
        .O(\block_w3_reg[30]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[31]_i_13 
       (.I0(\dec_block/op96_in [4]),
        .I1(\dec_block/p_0_in31_in [5]),
        .I2(\dec_block/op95_in [4]),
        .I3(\dec_block/op98_in [4]),
        .I4(\block_w3_reg[7]_i_4_n_0 ),
        .I5(\dec_block/op95_in [7]),
        .O(\block_w3_reg[31]_i_13_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[31]_i_14 
       (.I0(\dec_block/op95_in [5]),
        .I1(\dec_block/op98_in [5]),
        .O(\block_w3_reg[31]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[31]_i_4 
       (.I0(\dec_block/op98_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[31] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[31]_i_4__0 
       (.I0(\block_w3_reg[31]_i_6__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[31]_i_7__0_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[31]_i_8_n_0 ),
        .O(round_key[31]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[31]_i_6 
       (.I0(\block_w3_reg[31]_i_8_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[31]_i_7__0_n_0 ),
        .I3(\block_w0_reg_reg[31]_2 ),
        .I4(\block_w3_reg[31]_i_6__0_n_0 ),
        .I5(dec_new_block[31]),
        .O(\dec_block/op98_in [7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[31]_i_6__0 
       (.I0(\block_w3_reg[31]_i_9__0_n_0 ),
        .I1(\key_mem_reg[14]_14 [31]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [31]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [31]),
        .O(\block_w3_reg[31]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[31]_i_7 
       (.I0(round_key[31]),
        .I1(core_block[31]),
        .O(p_0_out[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[31]_i_7__0 
       (.I0(\key_mem_reg[7]_7 [31]),
        .I1(\key_mem_reg[6]_6 [31]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [31]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [31]),
        .O(\block_w3_reg[31]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[31]_i_8 
       (.I0(\key_mem_reg[3]_3 [31]),
        .I1(\key_mem_reg[2]_2 [31]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [31]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [31]),
        .O(\block_w3_reg[31]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[31]_i_9 
       (.I0(\block_w3_reg[31]_i_13_n_0 ),
        .I1(\dec_block/op98_in [6]),
        .I2(\dec_block/op96_in [6]),
        .I3(\dec_block/op96_in [7]),
        .I4(\block_w3_reg[31]_i_14_n_0 ),
        .O(inv_mixcolumns_return0124_out__47[7]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[31]_i_9__0 
       (.I0(\key_mem_reg[11]_11 [31]),
        .I1(\key_mem_reg[10]_10 [31]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [31]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [31]),
        .O(\block_w3_reg[31]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[3]_i_10 
       (.I0(\dec_block/op190_in [7]),
        .I1(round_key[115]),
        .I2(dec_new_block[115]),
        .I3(dec_new_block[107]),
        .I4(round_key[107]),
        .O(\block_w3_reg[3]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[3]_i_11 
       (.I0(\dec_block/p_0_in54_in [3]),
        .I1(\dec_block/op191_in [5]),
        .I2(\dec_block/p_0_in54_in [6]),
        .I3(\dec_block/op190_in [5]),
        .I4(\dec_block/op193_in [5]),
        .O(\block_w3_reg[3]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w3_reg[3]_i_12 
       (.I0(dec_new_block[122]),
        .I1(round_key[122]),
        .I2(\dec_block/p_0_in54_in [7]),
        .I3(\dec_block/op191_in [6]),
        .O(\block_w3_reg[3]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \block_w3_reg[3]_i_13 
       (.I0(dec_new_block[123]),
        .I1(round_key[123]),
        .I2(\dec_block/op191_in [7]),
        .O(\block_w3_reg[3]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[3]_i_2__0 
       (.I0(\dec_block/p_0_in31_in [4]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[3] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[3]_i_3 
       (.I0(\block_w3_reg[3]_i_6__0_n_0 ),
        .I1(\block_w3_reg_reg[26] ),
        .I2(\block_w3_reg[3]_i_7_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[3]_i_8_n_0 ),
        .O(round_key[3]));
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[3]_i_4__0 
       (.I0(round_key[3]),
        .I1(dec_new_block[3]),
        .O(\dec_block/p_0_in31_in [4]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[3]_i_5 
       (.I0(round_key[3]),
        .I1(core_block[3]),
        .O(addroundkey_return[2]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[3]_i_6 
       (.I0(\block_w3_reg[3]_i_9_n_0 ),
        .I1(\block_w2_reg[9]_i_6_n_0 ),
        .I2(\block_w3_reg[3]_i_10_n_0 ),
        .I3(\block_w3_reg[3]_i_11_n_0 ),
        .I4(\block_w3_reg[3]_i_12_n_0 ),
        .I5(\block_w3_reg[3]_i_13_n_0 ),
        .O(inv_mixcolumns_return0198_out__63[2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[3]_i_6__0 
       (.I0(\block_w3_reg[3]_i_9__0_n_0 ),
        .I1(\key_mem_reg[14]_14 [3]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [3]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [3]),
        .O(\block_w3_reg[3]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[3]_i_7 
       (.I0(\key_mem_reg[7]_7 [3]),
        .I1(\key_mem_reg[6]_6 [3]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [3]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [3]),
        .O(\block_w3_reg[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[3]_i_8 
       (.I0(\key_mem_reg[3]_3 [3]),
        .I1(\key_mem_reg[2]_2 [3]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [3]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [3]),
        .O(\block_w3_reg[3]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w3_reg[3]_i_9 
       (.I0(\dec_block/op193_in [0]),
        .I1(\dec_block/op190_in [0]),
        .I2(\block_w0_reg_reg[0] ),
        .I3(\block_w0_reg_reg[16] ),
        .O(\block_w3_reg[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[3]_i_9__0 
       (.I0(\key_mem_reg[11]_11 [3]),
        .I1(\key_mem_reg[10]_10 [3]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [3]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [3]),
        .O(\block_w3_reg[3]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[4]_i_10 
       (.I0(\dec_block/op193_in [5]),
        .I1(\dec_block/op190_in [5]),
        .I2(\dec_block/p_0_in54_in [6]),
        .I3(\dec_block/op191_in [5]),
        .I4(\dec_block/op190_in [1]),
        .I5(\dec_block/op193_in [1]),
        .O(\block_w3_reg[4]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[4]_i_10__0 
       (.I0(\key_mem_reg[11]_11 [4]),
        .I1(\key_mem_reg[10]_10 [4]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [4]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [4]),
        .O(\block_w3_reg[4]_i_10__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[4]_i_2__0 
       (.I0(\dec_block/p_0_in31_in [5]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[4] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[4]_i_3 
       (.I0(\block_w3_reg[4]_i_7_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[4]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[4]_i_9__0_n_0 ),
        .O(round_key[4]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[4]_i_4 
       (.I0(\block_w3_reg[4]_i_9__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[4]_i_8_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[4]_i_7_n_0 ),
        .I5(dec_new_block[4]),
        .O(\dec_block/p_0_in31_in [5]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[4]_i_6 
       (.I0(\block_w3_reg[4]_i_9_n_0 ),
        .I1(\dec_block/op191_in [4]),
        .I2(\block_w3_reg[4]_i_10_n_0 ),
        .I3(\block_w2_reg[9]_i_6_n_0 ),
        .I4(\block_w3_reg[5]_i_11_n_0 ),
        .I5(\block_w3_reg[6]_i_12_n_0 ),
        .O(inv_mixcolumns_return0198_out__63[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[4]_i_6__0 
       (.I0(round_key[4]),
        .I1(core_block[4]),
        .O(addroundkey_return[3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[4]_i_7 
       (.I0(\block_w3_reg[4]_i_10__0_n_0 ),
        .I1(\key_mem_reg[14]_14 [4]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [4]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [4]),
        .O(\block_w3_reg[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[4]_i_8 
       (.I0(\key_mem_reg[7]_7 [4]),
        .I1(\key_mem_reg[6]_6 [4]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [4]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [4]),
        .O(\block_w3_reg[4]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[4]_i_9 
       (.I0(\dec_block/op190_in [4]),
        .I1(\dec_block/op193_in [4]),
        .O(\block_w3_reg[4]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[4]_i_9__0 
       (.I0(\key_mem_reg[3]_3 [4]),
        .I1(\key_mem_reg[2]_2 [4]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [4]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [4]),
        .O(\block_w3_reg[4]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[5]_i_10 
       (.I0(\dec_block/op191_in [6]),
        .I1(\dec_block/p_0_in54_in [7]),
        .I2(round_key[122]),
        .I3(dec_new_block[122]),
        .I4(\dec_block/op190_in [2]),
        .O(\block_w3_reg[5]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[5]_i_11 
       (.I0(\dec_block/op190_in [6]),
        .I1(\dec_block/op193_in [6]),
        .I2(round_key[114]),
        .I3(dec_new_block[114]),
        .I4(\dec_block/p_0_in54_in [3]),
        .O(\block_w3_reg[5]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[5]_i_12 
       (.I0(\dec_block/p_0_in54_in [5]),
        .I1(\dec_block/op193_in [4]),
        .O(\block_w3_reg[5]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[5]_i_13 
       (.I0(\dec_block/op190_in [5]),
        .I1(\dec_block/op193_in [5]),
        .O(\block_w3_reg[5]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[5]_i_14 
       (.I0(\dec_block/op193_in [7]),
        .I1(round_key[99]),
        .I2(dec_new_block[99]),
        .I3(\dec_block/op190_in [7]),
        .I4(round_key[115]),
        .I5(dec_new_block[115]),
        .O(\block_w3_reg[5]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[5]_i_2__0 
       (.I0(\dec_block/p_0_in31_in [6]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[5] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[5]_i_3 
       (.I0(\block_w3_reg[5]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[5]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[5]_i_7__0_n_0 ),
        .O(round_key[5]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[5]_i_4 
       (.I0(\block_w3_reg[5]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[5]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[5]_i_5__0_n_0 ),
        .I5(dec_new_block[5]),
        .O(\dec_block/p_0_in31_in [6]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[5]_i_5 
       (.I0(round_key[101]),
        .I1(core_block[101]),
        .O(p_0_out[50]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[5]_i_5__0 
       (.I0(\block_w3_reg[5]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [5]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [5]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [5]),
        .O(\block_w3_reg[5]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[5]_i_6 
       (.I0(\key_mem_reg[7]_7 [5]),
        .I1(\key_mem_reg[6]_6 [5]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [5]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [5]),
        .O(\block_w3_reg[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[5]_i_7 
       (.I0(\block_w3_reg[5]_i_10_n_0 ),
        .I1(\block_w3_reg[5]_i_11_n_0 ),
        .I2(\block_w3_reg[5]_i_12_n_0 ),
        .I3(\dec_block/op191_in [5]),
        .I4(\block_w3_reg[5]_i_13_n_0 ),
        .I5(\block_w3_reg[5]_i_14_n_0 ),
        .O(inv_mixcolumns_return0198_out__63[4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[5]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [5]),
        .I1(\key_mem_reg[2]_2 [5]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [5]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [5]),
        .O(\block_w3_reg[5]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[5]_i_8 
       (.I0(\key_mem_reg[11]_11 [5]),
        .I1(\key_mem_reg[10]_10 [5]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [5]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [5]),
        .O(\block_w3_reg[5]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[6]_i_10 
       (.I0(\dec_block/op191_in [4]),
        .I1(\dec_block/p_0_in54_in [5]),
        .O(\block_w3_reg[6]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[6]_i_11 
       (.I0(\block_w0_reg[7]_i_4_n_0 ),
        .I1(round_key[107]),
        .I2(dec_new_block[107]),
        .I3(\dec_block/op190_in [7]),
        .I4(round_key[115]),
        .I5(dec_new_block[115]),
        .O(\block_w3_reg[6]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[6]_i_12 
       (.I0(\dec_block/op193_in [7]),
        .I1(round_key[99]),
        .I2(dec_new_block[99]),
        .I3(\dec_block/op191_in [7]),
        .I4(round_key[123]),
        .I5(dec_new_block[123]),
        .O(\block_w3_reg[6]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[6]_i_13 
       (.I0(\dec_block/p_0_in54_in [6]),
        .I1(\dec_block/op193_in [5]),
        .O(\block_w3_reg[6]_i_13_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[6]_i_14 
       (.I0(\dec_block/op190_in [6]),
        .I1(\dec_block/op193_in [6]),
        .O(\block_w3_reg[6]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[6]_i_2__0 
       (.I0(\dec_block/p_0_in31_in [7]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[6] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[6]_i_3 
       (.I0(\block_w3_reg[6]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[6]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[6]_i_7__0_n_0 ),
        .O(round_key[6]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[6]_i_4 
       (.I0(\block_w3_reg[6]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[6]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[6]_i_5__0_n_0 ),
        .I5(dec_new_block[6]),
        .O(\dec_block/p_0_in31_in [7]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[6]_i_5 
       (.I0(round_key[102]),
        .I1(core_block[102]),
        .O(p_0_out[51]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[6]_i_5__0 
       (.I0(\block_w3_reg[6]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [6]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [6]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [6]),
        .O(\block_w3_reg[6]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[6]_i_6 
       (.I0(\key_mem_reg[7]_7 [6]),
        .I1(\key_mem_reg[6]_6 [6]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [6]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [6]),
        .O(\block_w3_reg[6]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[6]_i_7 
       (.I0(\block_w3_reg[6]_i_10_n_0 ),
        .I1(\block_w3_reg[6]_i_11_n_0 ),
        .I2(\block_w3_reg[6]_i_12_n_0 ),
        .I3(\block_w3_reg[6]_i_13_n_0 ),
        .I4(\block_w3_reg[6]_i_14_n_0 ),
        .I5(\dec_block/op191_in [6]),
        .O(inv_mixcolumns_return0198_out__63[5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[6]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [6]),
        .I1(\key_mem_reg[2]_2 [6]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [6]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [6]),
        .O(\block_w3_reg[6]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[6]_i_8 
       (.I0(\key_mem_reg[11]_11 [6]),
        .I1(\key_mem_reg[10]_10 [6]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [6]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [6]),
        .O(\block_w3_reg[6]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[7]_i_11 
       (.I0(\dec_block/op191_in [4]),
        .I1(\dec_block/p_0_in54_in [5]),
        .I2(\dec_block/op190_in [4]),
        .I3(\dec_block/op193_in [4]),
        .I4(\dec_block/op193_in [7]),
        .I5(\dec_block/op191_in [7]),
        .O(\block_w3_reg[7]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[7]_i_12 
       (.I0(\dec_block/op191_in [5]),
        .I1(\dec_block/p_0_in54_in [6]),
        .O(\block_w3_reg[7]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[7]_i_2__0 
       (.I0(\block_w3_reg[7]_i_4_n_0 ),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[7] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[7]_i_3 
       (.I0(\block_w3_reg[7]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[7]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[7]_i_7__0_n_0 ),
        .O(round_key[7]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[7]_i_4 
       (.I0(\block_w3_reg[7]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[7]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[7]_i_5__0_n_0 ),
        .I5(dec_new_block[7]),
        .O(\block_w3_reg[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[7]_i_5 
       (.I0(round_key[103]),
        .I1(core_block[103]),
        .O(p_0_out[52]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[7]_i_5__0 
       (.I0(\block_w3_reg[7]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [7]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [7]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [7]),
        .O(\block_w3_reg[7]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[7]_i_6 
       (.I0(\key_mem_reg[7]_7 [7]),
        .I1(\key_mem_reg[6]_6 [7]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [7]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [7]),
        .O(\block_w3_reg[7]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[7]_i_7 
       (.I0(\block_w3_reg[7]_i_11_n_0 ),
        .I1(\dec_block/op193_in [6]),
        .I2(\dec_block/p_0_in54_in [7]),
        .I3(\dec_block/op190_in [7]),
        .I4(\block_w3_reg[7]_i_12_n_0 ),
        .O(inv_mixcolumns_return0198_out__63[6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[7]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [7]),
        .I1(\key_mem_reg[2]_2 [7]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [7]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [7]),
        .O(\block_w3_reg[7]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[7]_i_8 
       (.I0(\key_mem_reg[11]_11 [7]),
        .I1(\key_mem_reg[10]_10 [7]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [7]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [7]),
        .O(\block_w3_reg[7]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \block_w3_reg[8]_i_10 
       (.I0(\dec_block/op158_in [5]),
        .I1(\dec_block/op161_in [5]),
        .I2(\dec_block/p_0_in46_in [6]),
        .I3(\dec_block/op159_in [5]),
        .O(\block_w3_reg[8]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[8]_i_11 
       (.I0(\block_w1_reg[7]_i_4_n_0 ),
        .I1(\dec_block/op158_in [7]),
        .O(\block_w3_reg[8]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[8]_i_12 
       (.I0(\block_w1_reg_reg[16] ),
        .I1(\block_w1_reg_reg[0] ),
        .O(\block_w3_reg[8]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[8]_i_2__0 
       (.I0(\dec_block/op95_in [0]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[8] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[8]_i_3 
       (.I0(\block_w3_reg[8]_i_5__0_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[8]_i_6_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[8]_i_7__0_n_0 ),
        .O(round_key[8]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[8]_i_4 
       (.I0(\block_w3_reg[8]_i_7__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[8]_i_6_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[8]_i_5__0_n_0 ),
        .I5(dec_new_block[8]),
        .O(\dec_block/op95_in [0]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[8]_i_5 
       (.I0(round_key[72]),
        .I1(core_block[72]),
        .O(p_0_out[30]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[8]_i_5__0 
       (.I0(\block_w3_reg[8]_i_8_n_0 ),
        .I1(\key_mem_reg[14]_14 [8]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [8]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [8]),
        .O(\block_w3_reg[8]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[8]_i_6 
       (.I0(\key_mem_reg[7]_7 [8]),
        .I1(\key_mem_reg[6]_6 [8]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [8]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [8]),
        .O(\block_w3_reg[8]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[8]_i_7 
       (.I0(\block_w3_reg[8]_i_10_n_0 ),
        .I1(\dec_block/op161_in [0]),
        .I2(\block_w3_reg[8]_i_11_n_0 ),
        .I3(\block_w3_reg[8]_i_12_n_0 ),
        .I4(\block_w3_reg[11]_i_9_n_0 ),
        .O(inv_mixcolumns_return0174_out__63[0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[8]_i_7__0 
       (.I0(\key_mem_reg[3]_3 [8]),
        .I1(\key_mem_reg[2]_2 [8]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [8]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [8]),
        .O(\block_w3_reg[8]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[8]_i_8 
       (.I0(\key_mem_reg[11]_11 [8]),
        .I1(\key_mem_reg[10]_10 [8]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [8]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [8]),
        .O(\block_w3_reg[8]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \block_w3_reg[9]_i_10 
       (.I0(\dec_block/op161_in [1]),
        .I1(\dec_block/op159_in [5]),
        .I2(\dec_block/p_0_in46_in [6]),
        .I3(\dec_block/op161_in [5]),
        .I4(\dec_block/op158_in [5]),
        .O(\block_w3_reg[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[9]_i_10__0 
       (.I0(\key_mem_reg[11]_11 [9]),
        .I1(\key_mem_reg[10]_10 [9]),
        .I2(\block_w0_reg[31]_i_6__0_0 ),
        .I3(\key_mem_reg[9]_9 [9]),
        .I4(\block_w0_reg[31]_i_6__0_1 ),
        .I5(\key_mem_reg[8]_8 [9]),
        .O(\block_w3_reg[9]_i_10__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \block_w3_reg[9]_i_2__0 
       (.I0(\dec_block/op95_in [1]),
        .I1(\block_w0_reg_reg[31]_1 ),
        .O(\block_w3_reg_reg[9] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \block_w3_reg[9]_i_3 
       (.I0(\block_w3_reg[9]_i_7_n_0 ),
        .I1(\block_w0_reg_reg[31]_2 ),
        .I2(\block_w3_reg[9]_i_8_n_0 ),
        .I3(muxed_round_nr[2]),
        .I4(\block_w3_reg[9]_i_9__0_n_0 ),
        .O(round_key[9]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \block_w3_reg[9]_i_4 
       (.I0(\block_w3_reg[9]_i_9__0_n_0 ),
        .I1(muxed_round_nr[2]),
        .I2(\block_w3_reg[9]_i_8_n_0 ),
        .I3(\block_w3_reg_reg[26] ),
        .I4(\block_w3_reg[9]_i_7_n_0 ),
        .I5(dec_new_block[9]),
        .O(\dec_block/op95_in [1]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \block_w3_reg[9]_i_6 
       (.I0(\block_w3_reg[12]_i_10_n_0 ),
        .I1(\block_w3_reg[14]_i_14_n_0 ),
        .I2(\dec_block/op158_in [0]),
        .I3(\block_w3_reg[9]_i_9_n_0 ),
        .I4(\block_w3_reg[9]_i_10_n_0 ),
        .I5(\block_w1_reg_reg[0] ),
        .O(inv_mixcolumns_return0174_out__63[1]));
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[9]_i_6__0 
       (.I0(round_key[9]),
        .I1(core_block[9]),
        .O(addroundkey_return[8]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[9]_i_7 
       (.I0(\block_w3_reg[9]_i_10__0_n_0 ),
        .I1(\key_mem_reg[14]_14 [9]),
        .I2(\block_w3_reg[1]_i_4__0_0 ),
        .I3(\key_mem_reg[13]_13 [9]),
        .I4(\block_w2_reg[31]_i_21_n_0 ),
        .I5(\key_mem_reg[12]_12 [9]),
        .O(\block_w3_reg[9]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[9]_i_8 
       (.I0(\key_mem_reg[7]_7 [9]),
        .I1(\key_mem_reg[6]_6 [9]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[5]_5 [9]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[4]_4 [9]),
        .O(\block_w3_reg[9]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \block_w3_reg[9]_i_9 
       (.I0(\block_w1_reg[7]_i_4_n_0 ),
        .I1(\dec_block/op161_in [7]),
        .O(\block_w3_reg[9]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \block_w3_reg[9]_i_9__0 
       (.I0(\key_mem_reg[3]_3 [9]),
        .I1(\key_mem_reg[2]_2 [9]),
        .I2(\block_w3_reg[30]_i_4_0 ),
        .I3(\key_mem_reg[1]_1 [9]),
        .I4(\block_w3_reg[30]_i_4_1 ),
        .I5(\key_mem_reg[0]_0 [9]),
        .O(\block_w3_reg[9]_i_9__0_n_0 ));
  LUT3 #(
    .INIT(8'h54)) 
    g0_b0_i_8__6
       (.I0(ready_reg_reg_0[1]),
        .I1(p_1_in[0]),
        .I2(ready_reg_reg_0[0]),
        .O(init_state));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][0]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[0]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[0]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[128]),
        .O(key_mem_new[0]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][100]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[100]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[100]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[228]),
        .O(key_mem_new[100]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][101]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[101]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[101]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[229]),
        .O(key_mem_new[101]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][102]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[102]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[102]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[230]),
        .O(key_mem_new[102]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][103]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[103]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[103]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[231]),
        .O(key_mem_new[103]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][104]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[104]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[104]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[232]),
        .O(key_mem_new[104]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][105]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[105]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[105]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[233]),
        .O(key_mem_new[105]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][106]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[106]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[106]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[234]),
        .O(key_mem_new[106]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][107]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[107]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[107]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[235]),
        .O(key_mem_new[107]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][108]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[108]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[108]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[236]),
        .O(key_mem_new[108]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][109]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[109]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[109]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[237]),
        .O(key_mem_new[109]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][10]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[10]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[10]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[138]),
        .O(key_mem_new[10]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][110]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[110]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[110]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[238]),
        .O(key_mem_new[110]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][111]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[111]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[111]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[239]),
        .O(key_mem_new[111]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][112]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[112]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[112]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[240]),
        .O(key_mem_new[112]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][113]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[113]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[113]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[241]),
        .O(key_mem_new[113]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][114]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[114]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[114]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[242]),
        .O(key_mem_new[114]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][115]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[115]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[115]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[243]),
        .O(key_mem_new[115]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][116]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[116]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[116]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[244]),
        .O(key_mem_new[116]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][117]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[117]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[117]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[245]),
        .O(key_mem_new[117]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][118]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[118]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[118]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[246]),
        .O(key_mem_new[118]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][119]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[119]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[119]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[247]),
        .O(key_mem_new[119]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][11]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[11]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[11]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[139]),
        .O(key_mem_new[11]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][120]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[120]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[120]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[248]),
        .O(key_mem_new[120]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][121]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[121]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[121]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[249]),
        .O(key_mem_new[121]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][122]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[122]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[122]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[250]),
        .O(key_mem_new[122]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][123]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[123]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[123]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[251]),
        .O(key_mem_new[123]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][124]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[124]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[124]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[252]),
        .O(key_mem_new[124]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][125]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[125]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[125]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[253]),
        .O(key_mem_new[125]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][126]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[126]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[126]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[254]),
        .O(key_mem_new[126]));
  LUT2 #(
    .INIT(4'h8)) 
    \key_mem[0][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .O(key_mem));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][127]_i_2 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[127]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[127]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[255]),
        .O(key_mem_new[127]));
  LUT4 #(
    .INIT(16'h0001)) 
    \key_mem[0][127]_i_3 
       (.I0(\round_ctr_reg_reg_n_0_[2] ),
        .I1(\round_ctr_reg_reg_n_0_[3] ),
        .I2(p_0_in0),
        .I3(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(\key_mem[0][127]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][12]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[12]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[12]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[140]),
        .O(key_mem_new[12]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][13]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[13]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[13]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[141]),
        .O(key_mem_new[13]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][14]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[14]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[14]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[142]),
        .O(key_mem_new[14]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][15]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[15]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[15]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[143]),
        .O(key_mem_new[15]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][16]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[16]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[16]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[144]),
        .O(key_mem_new[16]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][17]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[17]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[17]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[145]),
        .O(key_mem_new[17]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][18]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[18]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[18]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[146]),
        .O(key_mem_new[18]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][19]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[19]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[19]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[147]),
        .O(key_mem_new[19]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][1]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[1]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[1]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[129]),
        .O(key_mem_new[1]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][20]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[20]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[20]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[148]),
        .O(key_mem_new[20]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][21]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[21]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[21]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[149]),
        .O(key_mem_new[21]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][22]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[22]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[22]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[150]),
        .O(key_mem_new[22]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][23]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[23]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[23]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[151]),
        .O(key_mem_new[23]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][24]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[24]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[24]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[152]),
        .O(key_mem_new[24]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][25]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[25]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[25]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[153]),
        .O(key_mem_new[25]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][26]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[26]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[26]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[154]),
        .O(key_mem_new[26]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][27]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[27]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[27]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[155]),
        .O(key_mem_new[27]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][28]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[28]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[28]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[156]),
        .O(key_mem_new[28]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][29]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[29]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[29]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[157]),
        .O(key_mem_new[29]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][2]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[2]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[2]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[130]),
        .O(key_mem_new[2]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][30]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[30]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[30]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[158]),
        .O(key_mem_new[30]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][31]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[31]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[31]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[159]),
        .O(key_mem_new[31]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][32]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[32]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[32]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[160]),
        .O(key_mem_new[32]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][33]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[33]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[33]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[161]),
        .O(key_mem_new[33]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][34]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[34]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[34]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[162]),
        .O(key_mem_new[34]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][35]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[35]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[35]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[163]),
        .O(key_mem_new[35]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][36]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[36]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[36]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[164]),
        .O(key_mem_new[36]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][37]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[37]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[37]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[165]),
        .O(key_mem_new[37]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][38]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[38]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[38]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[166]),
        .O(key_mem_new[38]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][39]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[39]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[39]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[167]),
        .O(key_mem_new[39]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][3]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[3]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[3]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[131]),
        .O(key_mem_new[3]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][40]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[40]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[40]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[168]),
        .O(key_mem_new[40]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][41]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[41]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[41]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[169]),
        .O(key_mem_new[41]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][42]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[42]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[42]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[170]),
        .O(key_mem_new[42]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][43]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[43]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[43]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[171]),
        .O(key_mem_new[43]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][44]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[44]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[44]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[172]),
        .O(key_mem_new[44]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][45]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[45]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[45]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[173]),
        .O(key_mem_new[45]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][46]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[46]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[46]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[174]),
        .O(key_mem_new[46]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][47]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[47]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[47]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[175]),
        .O(key_mem_new[47]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][48]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[48]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[48]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[176]),
        .O(key_mem_new[48]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][49]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[49]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[49]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[177]),
        .O(key_mem_new[49]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][4]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[4]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[4]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[132]),
        .O(key_mem_new[4]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][50]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[50]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[50]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[178]),
        .O(key_mem_new[50]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][51]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[51]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[51]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[179]),
        .O(key_mem_new[51]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][52]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[52]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[52]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[180]),
        .O(key_mem_new[52]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][53]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[53]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[53]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[181]),
        .O(key_mem_new[53]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][54]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[54]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[54]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[182]),
        .O(key_mem_new[54]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][55]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[55]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[55]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[183]),
        .O(key_mem_new[55]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][56]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[56]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[56]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[184]),
        .O(key_mem_new[56]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][57]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[57]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[57]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[185]),
        .O(key_mem_new[57]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][58]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[58]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[58]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[186]),
        .O(key_mem_new[58]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][59]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[59]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[59]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[187]),
        .O(key_mem_new[59]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][5]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[5]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[5]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[133]),
        .O(key_mem_new[5]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][60]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[60]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[60]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[188]),
        .O(key_mem_new[60]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][61]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[61]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[61]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[189]),
        .O(key_mem_new[61]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][62]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[62]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[62]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[190]),
        .O(key_mem_new[62]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][63]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[63]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[63]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[191]),
        .O(key_mem_new[63]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][64]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[64]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[64]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[192]),
        .O(key_mem_new[64]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][65]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[65]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[65]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[193]),
        .O(key_mem_new[65]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][66]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[66]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[66]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[194]),
        .O(key_mem_new[66]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][67]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[67]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[67]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[195]),
        .O(key_mem_new[67]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][68]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[68]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[68]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[196]),
        .O(key_mem_new[68]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][69]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[69]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[69]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[197]),
        .O(key_mem_new[69]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][6]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[6]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[6]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[134]),
        .O(key_mem_new[6]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][70]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[70]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[70]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[198]),
        .O(key_mem_new[70]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][71]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[71]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[71]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[199]),
        .O(key_mem_new[71]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][72]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[72]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[72]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[200]),
        .O(key_mem_new[72]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][73]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[73]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[73]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[201]),
        .O(key_mem_new[73]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][74]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[74]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[74]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[202]),
        .O(key_mem_new[74]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][75]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[75]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[75]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[203]),
        .O(key_mem_new[75]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][76]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[76]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[76]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[204]),
        .O(key_mem_new[76]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][77]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[77]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[77]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[205]),
        .O(key_mem_new[77]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][78]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[78]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[78]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[206]),
        .O(key_mem_new[78]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][79]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[79]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[79]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[207]),
        .O(key_mem_new[79]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][7]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[7]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[7]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[135]),
        .O(key_mem_new[7]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][80]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[80]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[80]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[208]),
        .O(key_mem_new[80]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][81]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[81]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[81]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[209]),
        .O(key_mem_new[81]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][82]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[82]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[82]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[210]),
        .O(key_mem_new[82]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][83]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[83]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[83]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[211]),
        .O(key_mem_new[83]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][84]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[84]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[84]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[212]),
        .O(key_mem_new[84]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][85]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[85]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[85]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[213]),
        .O(key_mem_new[85]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][86]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[86]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[86]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[214]),
        .O(key_mem_new[86]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][87]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[87]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[87]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[215]),
        .O(key_mem_new[87]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][88]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[88]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[88]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[216]),
        .O(key_mem_new[88]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][89]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[89]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[89]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[217]),
        .O(key_mem_new[89]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][8]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[8]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[8]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[136]),
        .O(key_mem_new[8]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][90]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[90]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[90]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[218]),
        .O(key_mem_new[90]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][91]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[91]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[91]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[219]),
        .O(key_mem_new[91]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][92]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[92]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[92]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[220]),
        .O(key_mem_new[92]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][93]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[93]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[93]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[221]),
        .O(key_mem_new[93]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][94]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[94]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[94]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[222]),
        .O(key_mem_new[94]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][95]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[95]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[95]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[223]),
        .O(key_mem_new[95]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][96]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[96]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[96]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[224]),
        .O(key_mem_new[96]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][97]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[97]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[97]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[225]),
        .O(key_mem_new[97]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][98]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[98]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[98]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[226]),
        .O(key_mem_new[98]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][99]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[99]),
        .I2(\key_mem_reg[14][127]_0 ),
        .I3(prev_key1_new[99]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[227]),
        .O(key_mem_new[99]));
  LUT6 #(
    .INIT(64'hA8A8A8080808A808)) 
    \key_mem[0][9]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(prev_key1_new0_in[9]),
        .I2(\key_mem_reg[14][36]_0 ),
        .I3(prev_key1_new[9]),
        .I4(\key_mem[0][127]_i_3_n_0 ),
        .I5(core_key[137]),
        .O(key_mem_new[9]));
  LUT5 #(
    .INIT(32'h00000080)) 
    \key_mem[10][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(p_0_in0),
        .I2(\round_ctr_reg_reg_n_0_[3] ),
        .I3(\round_ctr_reg_reg_n_0_[0] ),
        .I4(\round_ctr_reg_reg_n_0_[2] ),
        .O(\key_mem[10][127]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00008000)) 
    \key_mem[11][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\round_ctr_reg_reg_n_0_[0] ),
        .I2(p_0_in0),
        .I3(\round_ctr_reg_reg_n_0_[3] ),
        .I4(\round_ctr_reg_reg_n_0_[2] ),
        .O(\key_mem[11][127]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \key_mem[12][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\round_ctr_reg_reg_n_0_[3] ),
        .I2(\round_ctr_reg_reg_n_0_[2] ),
        .I3(\round_ctr_reg_reg_n_0_[0] ),
        .I4(p_0_in0),
        .O(\key_mem[12][127]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00008000)) 
    \key_mem[13][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\round_ctr_reg_reg_n_0_[0] ),
        .I2(\round_ctr_reg_reg_n_0_[3] ),
        .I3(\round_ctr_reg_reg_n_0_[2] ),
        .I4(p_0_in0),
        .O(\key_mem[13][127]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \key_mem[14][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(p_0_in0),
        .I2(\round_ctr_reg_reg_n_0_[3] ),
        .I3(\round_ctr_reg_reg_n_0_[0] ),
        .I4(\round_ctr_reg_reg_n_0_[2] ),
        .O(\key_mem[14][127]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \key_mem[1][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .O(\key_mem[1][127]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \key_mem[2][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I2(p_0_in0),
        .I3(\round_ctr_reg_reg_n_0_[3] ),
        .I4(\round_ctr_reg_reg_n_0_[2] ),
        .O(\key_mem[2][127]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \key_mem[3][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\round_ctr_reg_reg_n_0_[0] ),
        .I2(p_0_in0),
        .I3(\round_ctr_reg_reg_n_0_[3] ),
        .I4(\round_ctr_reg_reg_n_0_[2] ),
        .O(\key_mem[3][127]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \key_mem[4][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\round_ctr_reg_reg_n_0_[0] ),
        .I2(\round_ctr_reg_reg_n_0_[2] ),
        .I3(p_0_in0),
        .I4(\round_ctr_reg_reg_n_0_[3] ),
        .O(\key_mem[4][127]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \key_mem[5][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\round_ctr_reg_reg_n_0_[0] ),
        .I2(\round_ctr_reg_reg_n_0_[2] ),
        .I3(p_0_in0),
        .I4(\round_ctr_reg_reg_n_0_[3] ),
        .O(\key_mem[5][127]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \key_mem[6][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(p_0_in0),
        .I2(\round_ctr_reg_reg_n_0_[2] ),
        .I3(\round_ctr_reg_reg_n_0_[0] ),
        .I4(\round_ctr_reg_reg_n_0_[3] ),
        .O(\key_mem[6][127]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00008000)) 
    \key_mem[7][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\round_ctr_reg_reg_n_0_[0] ),
        .I2(p_0_in0),
        .I3(\round_ctr_reg_reg_n_0_[2] ),
        .I4(\round_ctr_reg_reg_n_0_[3] ),
        .O(\key_mem[7][127]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \key_mem[8][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\round_ctr_reg_reg_n_0_[0] ),
        .I2(\round_ctr_reg_reg_n_0_[3] ),
        .I3(p_0_in0),
        .I4(\round_ctr_reg_reg_n_0_[2] ),
        .O(\key_mem[8][127]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \key_mem[9][127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\round_ctr_reg_reg_n_0_[0] ),
        .I2(\round_ctr_reg_reg_n_0_[3] ),
        .I3(p_0_in0),
        .I4(\round_ctr_reg_reg_n_0_[2] ),
        .O(\key_mem[9][127]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][0] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[0]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][100] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[0]_0 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][101] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[0]_0 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][102] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[0]_0 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][103] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[0]_0 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][104] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[0]_0 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][105] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[0]_0 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][106] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[0]_0 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][107] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[0]_0 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][108] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[0]_0 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][109] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[0]_0 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][10] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[0]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][110] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[0]_0 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][111] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[0]_0 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][112] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[0]_0 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][113] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[0]_0 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][114] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[0]_0 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][115] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[0]_0 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][116] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[0]_0 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][117] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[0]_0 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][118] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[0]_0 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][119] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[0]_0 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][11] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[0]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][120] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[0]_0 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][121] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[0]_0 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][122] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[0]_0 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][123] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[0]_0 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][124] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[0]_0 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][125] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[0]_0 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][126] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[0]_0 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][127] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[0]_0 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][12] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[0]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][13] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[0]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][14] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[0]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][15] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[0]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][16] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[0]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][17] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[0]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][18] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[0]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][19] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[0]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][1] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[0]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][20] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[0]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][21] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[0]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][22] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[0]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][23] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[0]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][24] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[0]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][25] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[0]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][26] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[0]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][27] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[0]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][28] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[0]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][29] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[0]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][2] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[0]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][30] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[0]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][31] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[0]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][32] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[0]_0 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][33] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[0]_0 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][34] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[0]_0 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][35] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[0]_0 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][36] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[0]_0 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][37] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[0]_0 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][38] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[0]_0 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][39] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[0]_0 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][3] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[0]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][40] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[0]_0 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][41] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[0]_0 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][42] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[0]_0 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][43] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[0]_0 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][44] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[0]_0 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][45] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[0]_0 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][46] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[0]_0 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][47] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[0]_0 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][48] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[0]_0 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][49] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[0]_0 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][4] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[0]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][50] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[0]_0 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][51] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[0]_0 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][52] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[0]_0 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][53] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[0]_0 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][54] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[0]_0 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][55] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[0]_0 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][56] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[0]_0 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][57] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[0]_0 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][58] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[0]_0 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][59] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[0]_0 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][5] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[0]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][60] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[0]_0 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][61] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[0]_0 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][62] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[0]_0 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][63] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[0]_0 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][64] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[0]_0 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][65] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[0]_0 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][66] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[0]_0 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][67] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[0]_0 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][68] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[0]_0 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][69] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[0]_0 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][6] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[0]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][70] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[0]_0 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][71] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[0]_0 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][72] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[0]_0 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][73] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[0]_0 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][74] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[0]_0 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][75] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[0]_0 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][76] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[0]_0 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][77] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[0]_0 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][78] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[0]_0 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][79] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[0]_0 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][7] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[0]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][80] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[0]_0 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][81] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[0]_0 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][82] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[0]_0 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][83] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[0]_0 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][84] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[0]_0 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][85] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[0]_0 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][86] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[0]_0 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][87] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[0]_0 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][88] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[0]_0 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][89] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[0]_0 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][8] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[0]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][90] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[0]_0 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][91] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[0]_0 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][92] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[0]_0 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][93] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[0]_0 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][94] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[0]_0 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][95] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[0]_0 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][96] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[0]_0 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][97] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[0]_0 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][98] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[0]_0 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][99] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[0]_0 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[0][9] 
       (.C(clk_i),
        .CE(key_mem),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[0]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][0] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[10]_10 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][100] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[10]_10 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][101] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[10]_10 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][102] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[10]_10 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][103] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[10]_10 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][104] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[10]_10 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][105] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[10]_10 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][106] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[10]_10 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][107] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[10]_10 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][108] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[10]_10 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][109] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[10]_10 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][10] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[10]_10 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][110] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[10]_10 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][111] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[10]_10 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][112] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[10]_10 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][113] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[10]_10 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][114] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[10]_10 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][115] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[10]_10 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][116] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[10]_10 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][117] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[10]_10 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][118] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[10]_10 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][119] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[10]_10 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][11] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[10]_10 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][120] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[10]_10 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][121] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[10]_10 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][122] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[10]_10 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][123] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[10]_10 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][124] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[10]_10 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][125] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[10]_10 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][126] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[10]_10 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][127] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[10]_10 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][12] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[10]_10 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][13] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[10]_10 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][14] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[10]_10 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][15] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[10]_10 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][16] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[10]_10 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][17] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[10]_10 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][18] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[10]_10 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][19] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[10]_10 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][1] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[10]_10 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][20] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[10]_10 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][21] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[10]_10 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][22] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[10]_10 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][23] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[10]_10 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][24] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[10]_10 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][25] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[10]_10 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][26] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[10]_10 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][27] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[10]_10 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][28] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[10]_10 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][29] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[10]_10 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][2] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[10]_10 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][30] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[10]_10 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][31] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[10]_10 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][32] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[10]_10 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][33] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[10]_10 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][34] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[10]_10 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][35] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[10]_10 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][36] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[10]_10 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][37] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[10]_10 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][38] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[10]_10 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][39] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[10]_10 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][3] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[10]_10 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][40] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[10]_10 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][41] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[10]_10 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][42] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[10]_10 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][43] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[10]_10 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][44] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[10]_10 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][45] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[10]_10 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][46] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[10]_10 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][47] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[10]_10 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][48] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[10]_10 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][49] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[10]_10 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][4] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[10]_10 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][50] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[10]_10 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][51] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[10]_10 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][52] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[10]_10 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][53] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[10]_10 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][54] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[10]_10 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][55] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[10]_10 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][56] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[10]_10 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][57] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[10]_10 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][58] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[10]_10 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][59] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[10]_10 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][5] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[10]_10 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][60] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[10]_10 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][61] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[10]_10 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][62] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[10]_10 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][63] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[10]_10 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][64] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[10]_10 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][65] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[10]_10 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][66] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[10]_10 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][67] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[10]_10 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][68] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[10]_10 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][69] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[10]_10 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][6] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[10]_10 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][70] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[10]_10 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][71] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[10]_10 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][72] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[10]_10 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][73] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[10]_10 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][74] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[10]_10 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][75] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[10]_10 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][76] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[10]_10 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][77] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[10]_10 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][78] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[10]_10 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][79] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[10]_10 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][7] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[10]_10 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][80] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[10]_10 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][81] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[10]_10 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][82] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[10]_10 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][83] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[10]_10 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][84] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[10]_10 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][85] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[10]_10 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][86] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[10]_10 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][87] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[10]_10 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][88] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[10]_10 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][89] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[10]_10 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][8] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[10]_10 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][90] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[10]_10 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][91] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[10]_10 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][92] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[10]_10 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][93] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[10]_10 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][94] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[10]_10 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][95] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[10]_10 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][96] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[10]_10 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][97] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[10]_10 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][98] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[10]_10 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][99] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[10]_10 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[10][9] 
       (.C(clk_i),
        .CE(\key_mem[10][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[10]_10 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][0] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[11]_11 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][100] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[11]_11 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][101] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[11]_11 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][102] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[11]_11 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][103] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[11]_11 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][104] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[11]_11 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][105] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[11]_11 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][106] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[11]_11 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][107] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[11]_11 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][108] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[11]_11 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][109] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[11]_11 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][10] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[11]_11 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][110] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[11]_11 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][111] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[11]_11 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][112] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[11]_11 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][113] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[11]_11 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][114] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[11]_11 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][115] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[11]_11 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][116] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[11]_11 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][117] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[11]_11 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][118] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[11]_11 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][119] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[11]_11 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][11] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[11]_11 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][120] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[11]_11 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][121] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[11]_11 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][122] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[11]_11 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][123] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[11]_11 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][124] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[11]_11 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][125] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[11]_11 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][126] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[11]_11 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][127] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[11]_11 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][12] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[11]_11 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][13] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[11]_11 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][14] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[11]_11 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][15] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[11]_11 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][16] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[11]_11 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][17] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[11]_11 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][18] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[11]_11 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][19] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[11]_11 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][1] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[11]_11 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][20] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[11]_11 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][21] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[11]_11 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][22] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[11]_11 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][23] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[11]_11 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][24] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[11]_11 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][25] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[11]_11 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][26] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[11]_11 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][27] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[11]_11 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][28] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[11]_11 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][29] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[11]_11 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][2] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[11]_11 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][30] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[11]_11 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][31] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[11]_11 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][32] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[11]_11 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][33] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[11]_11 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][34] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[11]_11 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][35] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[11]_11 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][36] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[11]_11 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][37] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[11]_11 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][38] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[11]_11 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][39] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[11]_11 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][3] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[11]_11 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][40] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[11]_11 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][41] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[11]_11 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][42] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[11]_11 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][43] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[11]_11 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][44] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[11]_11 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][45] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[11]_11 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][46] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[11]_11 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][47] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[11]_11 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][48] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[11]_11 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][49] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[11]_11 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][4] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[11]_11 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][50] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[11]_11 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][51] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[11]_11 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][52] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[11]_11 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][53] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[11]_11 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][54] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[11]_11 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][55] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[11]_11 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][56] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[11]_11 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][57] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[11]_11 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][58] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[11]_11 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][59] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[11]_11 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][5] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[11]_11 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][60] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[11]_11 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][61] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[11]_11 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][62] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[11]_11 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][63] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[11]_11 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][64] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[11]_11 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][65] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[11]_11 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][66] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[11]_11 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][67] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[11]_11 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][68] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[11]_11 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][69] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[11]_11 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][6] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[11]_11 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][70] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[11]_11 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][71] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[11]_11 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][72] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[11]_11 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][73] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[11]_11 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][74] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[11]_11 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][75] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[11]_11 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][76] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[11]_11 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][77] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[11]_11 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][78] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[11]_11 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][79] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[11]_11 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][7] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[11]_11 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][80] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[11]_11 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][81] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[11]_11 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][82] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[11]_11 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][83] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[11]_11 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][84] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[11]_11 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][85] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[11]_11 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][86] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[11]_11 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][87] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[11]_11 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][88] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[11]_11 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][89] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[11]_11 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][8] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[11]_11 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][90] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[11]_11 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][91] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[11]_11 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][92] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[11]_11 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][93] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[11]_11 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][94] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[11]_11 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][95] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[11]_11 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][96] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[11]_11 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][97] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[11]_11 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][98] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[11]_11 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][99] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[11]_11 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[11][9] 
       (.C(clk_i),
        .CE(\key_mem[11][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[11]_11 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][0] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[12]_12 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][100] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[12]_12 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][101] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[12]_12 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][102] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[12]_12 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][103] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[12]_12 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][104] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[12]_12 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][105] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[12]_12 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][106] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[12]_12 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][107] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[12]_12 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][108] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[12]_12 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][109] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[12]_12 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][10] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[12]_12 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][110] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[12]_12 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][111] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[12]_12 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][112] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[12]_12 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][113] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[12]_12 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][114] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[12]_12 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][115] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[12]_12 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][116] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[12]_12 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][117] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[12]_12 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][118] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[12]_12 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][119] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[12]_12 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][11] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[12]_12 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][120] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[12]_12 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][121] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[12]_12 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][122] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[12]_12 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][123] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[12]_12 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][124] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[12]_12 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][125] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[12]_12 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][126] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[12]_12 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][127] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[12]_12 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][12] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[12]_12 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][13] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[12]_12 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][14] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[12]_12 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][15] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[12]_12 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][16] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[12]_12 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][17] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[12]_12 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][18] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[12]_12 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][19] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[12]_12 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][1] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[12]_12 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][20] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[12]_12 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][21] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[12]_12 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][22] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[12]_12 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][23] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[12]_12 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][24] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[12]_12 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][25] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[12]_12 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][26] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[12]_12 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][27] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[12]_12 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][28] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[12]_12 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][29] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[12]_12 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][2] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[12]_12 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][30] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[12]_12 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][31] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[12]_12 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][32] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[12]_12 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][33] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[12]_12 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][34] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[12]_12 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][35] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[12]_12 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][36] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[12]_12 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][37] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[12]_12 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][38] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[12]_12 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][39] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[12]_12 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][3] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[12]_12 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][40] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[12]_12 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][41] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[12]_12 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][42] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[12]_12 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][43] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[12]_12 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][44] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[12]_12 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][45] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[12]_12 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][46] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[12]_12 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][47] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[12]_12 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][48] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[12]_12 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][49] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[12]_12 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][4] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[12]_12 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][50] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[12]_12 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][51] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[12]_12 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][52] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[12]_12 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][53] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[12]_12 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][54] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[12]_12 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][55] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[12]_12 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][56] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[12]_12 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][57] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[12]_12 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][58] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[12]_12 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][59] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[12]_12 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][5] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[12]_12 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][60] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[12]_12 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][61] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[12]_12 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][62] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[12]_12 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][63] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[12]_12 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][64] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[12]_12 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][65] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[12]_12 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][66] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[12]_12 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][67] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[12]_12 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][68] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[12]_12 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][69] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[12]_12 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][6] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[12]_12 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][70] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[12]_12 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][71] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[12]_12 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][72] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[12]_12 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][73] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[12]_12 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][74] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[12]_12 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][75] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[12]_12 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][76] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[12]_12 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][77] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[12]_12 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][78] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[12]_12 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][79] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[12]_12 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][7] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[12]_12 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][80] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[12]_12 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][81] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[12]_12 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][82] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[12]_12 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][83] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[12]_12 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][84] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[12]_12 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][85] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[12]_12 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][86] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[12]_12 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][87] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[12]_12 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][88] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[12]_12 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][89] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[12]_12 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][8] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[12]_12 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][90] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[12]_12 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][91] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[12]_12 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][92] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[12]_12 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][93] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[12]_12 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][94] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[12]_12 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][95] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[12]_12 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][96] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[12]_12 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][97] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[12]_12 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][98] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[12]_12 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][99] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[12]_12 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[12][9] 
       (.C(clk_i),
        .CE(\key_mem[12][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[12]_12 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][0] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[13]_13 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][100] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[13]_13 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][101] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[13]_13 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][102] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[13]_13 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][103] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[13]_13 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][104] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[13]_13 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][105] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[13]_13 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][106] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[13]_13 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][107] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[13]_13 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][108] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[13]_13 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][109] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[13]_13 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][10] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[13]_13 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][110] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[13]_13 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][111] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[13]_13 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][112] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[13]_13 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][113] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[13]_13 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][114] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[13]_13 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][115] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[13]_13 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][116] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[13]_13 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][117] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[13]_13 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][118] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[13]_13 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][119] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[13]_13 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][11] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[13]_13 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][120] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[13]_13 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][121] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[13]_13 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][122] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[13]_13 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][123] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[13]_13 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][124] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[13]_13 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][125] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[13]_13 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][126] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[13]_13 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][127] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[13]_13 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][12] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[13]_13 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][13] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[13]_13 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][14] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[13]_13 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][15] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[13]_13 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][16] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[13]_13 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][17] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[13]_13 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][18] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[13]_13 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][19] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[13]_13 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][1] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[13]_13 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][20] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[13]_13 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][21] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[13]_13 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][22] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[13]_13 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][23] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[13]_13 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][24] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[13]_13 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][25] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[13]_13 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][26] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[13]_13 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][27] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[13]_13 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][28] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[13]_13 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][29] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[13]_13 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][2] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[13]_13 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][30] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[13]_13 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][31] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[13]_13 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][32] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[13]_13 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][33] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[13]_13 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][34] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[13]_13 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][35] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[13]_13 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][36] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[13]_13 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][37] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[13]_13 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][38] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[13]_13 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][39] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[13]_13 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][3] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[13]_13 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][40] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[13]_13 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][41] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[13]_13 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][42] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[13]_13 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][43] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[13]_13 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][44] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[13]_13 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][45] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[13]_13 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][46] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[13]_13 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][47] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[13]_13 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][48] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[13]_13 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][49] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[13]_13 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][4] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[13]_13 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][50] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[13]_13 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][51] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[13]_13 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][52] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[13]_13 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][53] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[13]_13 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][54] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[13]_13 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][55] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[13]_13 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][56] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[13]_13 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][57] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[13]_13 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][58] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[13]_13 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][59] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[13]_13 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][5] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[13]_13 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][60] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[13]_13 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][61] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[13]_13 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][62] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[13]_13 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][63] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[13]_13 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][64] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[13]_13 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][65] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[13]_13 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][66] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[13]_13 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][67] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[13]_13 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][68] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[13]_13 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][69] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[13]_13 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][6] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[13]_13 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][70] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[13]_13 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][71] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[13]_13 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][72] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[13]_13 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][73] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[13]_13 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][74] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[13]_13 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][75] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[13]_13 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][76] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[13]_13 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][77] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[13]_13 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][78] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[13]_13 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][79] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[13]_13 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][7] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[13]_13 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][80] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[13]_13 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][81] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[13]_13 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][82] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[13]_13 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][83] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[13]_13 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][84] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[13]_13 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][85] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[13]_13 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][86] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[13]_13 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][87] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[13]_13 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][88] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[13]_13 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][89] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[13]_13 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][8] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[13]_13 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][90] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[13]_13 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][91] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[13]_13 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][92] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[13]_13 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][93] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[13]_13 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][94] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[13]_13 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][95] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[13]_13 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][96] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[13]_13 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][97] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[13]_13 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][98] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[13]_13 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][99] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[13]_13 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[13][9] 
       (.C(clk_i),
        .CE(\key_mem[13][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[13]_13 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][0] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[14]_14 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][100] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[14]_14 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][101] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[14]_14 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][102] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[14]_14 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][103] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[14]_14 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][104] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[14]_14 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][105] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[14]_14 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][106] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[14]_14 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][107] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[14]_14 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][108] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[14]_14 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][109] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[14]_14 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][10] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[14]_14 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][110] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[14]_14 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][111] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[14]_14 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][112] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[14]_14 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][113] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[14]_14 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][114] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[14]_14 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][115] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[14]_14 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][116] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[14]_14 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][117] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[14]_14 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][118] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[14]_14 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][119] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[14]_14 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][11] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[14]_14 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][120] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[14]_14 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][121] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[14]_14 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][122] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[14]_14 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][123] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[14]_14 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][124] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[14]_14 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][125] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[14]_14 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][126] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[14]_14 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][127] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[14]_14 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][12] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[14]_14 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][13] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[14]_14 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][14] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[14]_14 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][15] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[14]_14 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][16] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[14]_14 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][17] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[14]_14 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][18] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[14]_14 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][19] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[14]_14 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][1] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[14]_14 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][20] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[14]_14 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][21] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[14]_14 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][22] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[14]_14 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][23] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[14]_14 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][24] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[14]_14 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][25] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[14]_14 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][26] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[14]_14 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][27] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[14]_14 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][28] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[14]_14 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][29] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[14]_14 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][2] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[14]_14 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][30] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[14]_14 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][31] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[14]_14 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][32] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[14]_14 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][33] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[14]_14 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][34] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[14]_14 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][35] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[14]_14 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][36] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[14]_14 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][37] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[14]_14 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][38] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[14]_14 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][39] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[14]_14 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][3] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[14]_14 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][40] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[14]_14 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][41] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[14]_14 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][42] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[14]_14 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][43] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[14]_14 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][44] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[14]_14 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][45] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[14]_14 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][46] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[14]_14 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][47] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[14]_14 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][48] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[14]_14 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][49] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[14]_14 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][4] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[14]_14 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][50] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[14]_14 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][51] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[14]_14 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][52] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[14]_14 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][53] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[14]_14 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][54] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[14]_14 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][55] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[14]_14 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][56] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[14]_14 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][57] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[14]_14 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][58] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[14]_14 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][59] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[14]_14 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][5] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[14]_14 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][60] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[14]_14 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][61] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[14]_14 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][62] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[14]_14 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][63] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[14]_14 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][64] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[14]_14 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][65] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[14]_14 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][66] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[14]_14 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][67] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[14]_14 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][68] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[14]_14 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][69] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[14]_14 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][6] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[14]_14 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][70] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[14]_14 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][71] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[14]_14 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][72] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[14]_14 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][73] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[14]_14 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][74] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[14]_14 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][75] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[14]_14 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][76] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[14]_14 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][77] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[14]_14 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][78] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[14]_14 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][79] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[14]_14 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][7] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[14]_14 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][80] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[14]_14 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][81] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[14]_14 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][82] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[14]_14 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][83] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[14]_14 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][84] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[14]_14 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][85] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[14]_14 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][86] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[14]_14 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][87] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[14]_14 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][88] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[14]_14 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][89] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[14]_14 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][8] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[14]_14 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][90] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[14]_14 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][91] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[14]_14 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][92] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[14]_14 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][93] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[14]_14 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][94] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[14]_14 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][95] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[14]_14 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][96] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[14]_14 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][97] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[14]_14 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][98] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[14]_14 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][99] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[14]_14 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[14][9] 
       (.C(clk_i),
        .CE(\key_mem[14][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[14]_14 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][0] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[1]_1 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][100] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[1]_1 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][101] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[1]_1 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][102] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[1]_1 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][103] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[1]_1 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][104] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[1]_1 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][105] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[1]_1 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][106] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[1]_1 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][107] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[1]_1 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][108] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[1]_1 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][109] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[1]_1 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][10] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[1]_1 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][110] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[1]_1 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][111] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[1]_1 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][112] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[1]_1 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][113] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[1]_1 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][114] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[1]_1 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][115] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[1]_1 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][116] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[1]_1 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][117] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[1]_1 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][118] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[1]_1 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][119] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[1]_1 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][11] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[1]_1 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][120] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[1]_1 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][121] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[1]_1 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][122] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[1]_1 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][123] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[1]_1 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][124] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[1]_1 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][125] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[1]_1 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][126] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[1]_1 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][127] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[1]_1 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][12] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[1]_1 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][13] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[1]_1 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][14] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[1]_1 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][15] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[1]_1 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][16] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[1]_1 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][17] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[1]_1 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][18] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[1]_1 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][19] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[1]_1 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][1] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[1]_1 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][20] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[1]_1 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][21] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[1]_1 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][22] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[1]_1 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][23] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[1]_1 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][24] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[1]_1 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][25] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[1]_1 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][26] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[1]_1 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][27] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[1]_1 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][28] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[1]_1 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][29] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[1]_1 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][2] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[1]_1 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][30] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[1]_1 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][31] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[1]_1 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][32] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[1]_1 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][33] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[1]_1 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][34] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[1]_1 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][35] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[1]_1 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][36] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[1]_1 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][37] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[1]_1 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][38] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[1]_1 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][39] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[1]_1 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][3] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[1]_1 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][40] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[1]_1 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][41] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[1]_1 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][42] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[1]_1 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][43] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[1]_1 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][44] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[1]_1 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][45] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[1]_1 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][46] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[1]_1 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][47] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[1]_1 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][48] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[1]_1 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][49] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[1]_1 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][4] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[1]_1 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][50] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[1]_1 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][51] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[1]_1 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][52] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[1]_1 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][53] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[1]_1 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][54] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[1]_1 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][55] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[1]_1 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][56] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[1]_1 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][57] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[1]_1 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][58] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[1]_1 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][59] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[1]_1 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][5] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[1]_1 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][60] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[1]_1 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][61] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[1]_1 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][62] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[1]_1 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][63] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[1]_1 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][64] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[1]_1 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][65] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[1]_1 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][66] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[1]_1 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][67] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[1]_1 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][68] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[1]_1 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][69] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[1]_1 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][6] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[1]_1 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][70] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[1]_1 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][71] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[1]_1 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][72] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[1]_1 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][73] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[1]_1 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][74] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[1]_1 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][75] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[1]_1 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][76] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[1]_1 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][77] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[1]_1 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][78] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[1]_1 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][79] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[1]_1 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][7] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[1]_1 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][80] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[1]_1 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][81] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[1]_1 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][82] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[1]_1 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][83] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[1]_1 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][84] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[1]_1 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][85] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[1]_1 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][86] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[1]_1 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][87] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[1]_1 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][88] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[1]_1 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][89] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[1]_1 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][8] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[1]_1 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][90] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[1]_1 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][91] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[1]_1 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][92] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[1]_1 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][93] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[1]_1 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][94] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[1]_1 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][95] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[1]_1 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][96] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[1]_1 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][97] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[1]_1 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][98] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[1]_1 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][99] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[1]_1 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[1][9] 
       (.C(clk_i),
        .CE(\key_mem[1][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[1]_1 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][0] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[2]_2 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][100] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[2]_2 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][101] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[2]_2 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][102] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[2]_2 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][103] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[2]_2 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][104] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[2]_2 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][105] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[2]_2 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][106] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[2]_2 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][107] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[2]_2 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][108] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[2]_2 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][109] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[2]_2 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][10] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[2]_2 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][110] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[2]_2 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][111] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[2]_2 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][112] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[2]_2 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][113] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[2]_2 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][114] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[2]_2 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][115] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[2]_2 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][116] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[2]_2 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][117] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[2]_2 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][118] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[2]_2 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][119] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[2]_2 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][11] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[2]_2 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][120] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[2]_2 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][121] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[2]_2 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][122] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[2]_2 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][123] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[2]_2 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][124] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[2]_2 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][125] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[2]_2 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][126] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[2]_2 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][127] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[2]_2 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][12] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[2]_2 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][13] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[2]_2 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][14] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[2]_2 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][15] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[2]_2 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][16] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[2]_2 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][17] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[2]_2 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][18] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[2]_2 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][19] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[2]_2 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][1] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[2]_2 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][20] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[2]_2 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][21] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[2]_2 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][22] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[2]_2 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][23] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[2]_2 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][24] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[2]_2 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][25] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[2]_2 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][26] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[2]_2 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][27] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[2]_2 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][28] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[2]_2 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][29] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[2]_2 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][2] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[2]_2 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][30] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[2]_2 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][31] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[2]_2 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][32] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[2]_2 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][33] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[2]_2 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][34] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[2]_2 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][35] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[2]_2 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][36] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[2]_2 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][37] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[2]_2 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][38] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[2]_2 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][39] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[2]_2 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][3] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[2]_2 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][40] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[2]_2 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][41] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[2]_2 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][42] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[2]_2 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][43] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[2]_2 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][44] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[2]_2 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][45] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[2]_2 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][46] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[2]_2 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][47] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[2]_2 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][48] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[2]_2 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][49] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[2]_2 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][4] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[2]_2 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][50] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[2]_2 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][51] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[2]_2 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][52] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[2]_2 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][53] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[2]_2 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][54] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[2]_2 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][55] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[2]_2 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][56] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[2]_2 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][57] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[2]_2 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][58] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[2]_2 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][59] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[2]_2 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][5] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[2]_2 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][60] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[2]_2 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][61] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[2]_2 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][62] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[2]_2 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][63] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[2]_2 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][64] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[2]_2 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][65] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[2]_2 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][66] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[2]_2 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][67] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[2]_2 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][68] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[2]_2 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][69] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[2]_2 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][6] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[2]_2 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][70] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[2]_2 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][71] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[2]_2 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][72] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[2]_2 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][73] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[2]_2 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][74] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[2]_2 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][75] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[2]_2 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][76] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[2]_2 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][77] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[2]_2 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][78] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[2]_2 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][79] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[2]_2 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][7] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[2]_2 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][80] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[2]_2 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][81] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[2]_2 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][82] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[2]_2 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][83] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[2]_2 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][84] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[2]_2 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][85] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[2]_2 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][86] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[2]_2 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][87] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[2]_2 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][88] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[2]_2 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][89] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[2]_2 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][8] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[2]_2 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][90] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[2]_2 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][91] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[2]_2 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][92] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[2]_2 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][93] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[2]_2 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][94] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[2]_2 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][95] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[2]_2 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][96] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[2]_2 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][97] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[2]_2 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][98] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[2]_2 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][99] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[2]_2 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[2][9] 
       (.C(clk_i),
        .CE(\key_mem[2][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[2]_2 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][0] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[3]_3 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][100] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[3]_3 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][101] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[3]_3 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][102] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[3]_3 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][103] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[3]_3 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][104] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[3]_3 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][105] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[3]_3 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][106] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[3]_3 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][107] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[3]_3 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][108] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[3]_3 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][109] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[3]_3 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][10] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[3]_3 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][110] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[3]_3 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][111] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[3]_3 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][112] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[3]_3 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][113] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[3]_3 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][114] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[3]_3 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][115] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[3]_3 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][116] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[3]_3 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][117] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[3]_3 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][118] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[3]_3 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][119] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[3]_3 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][11] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[3]_3 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][120] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[3]_3 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][121] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[3]_3 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][122] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[3]_3 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][123] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[3]_3 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][124] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[3]_3 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][125] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[3]_3 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][126] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[3]_3 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][127] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[3]_3 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][12] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[3]_3 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][13] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[3]_3 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][14] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[3]_3 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][15] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[3]_3 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][16] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[3]_3 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][17] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[3]_3 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][18] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[3]_3 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][19] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[3]_3 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][1] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[3]_3 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][20] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[3]_3 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][21] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[3]_3 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][22] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[3]_3 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][23] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[3]_3 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][24] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[3]_3 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][25] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[3]_3 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][26] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[3]_3 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][27] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[3]_3 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][28] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[3]_3 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][29] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[3]_3 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][2] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[3]_3 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][30] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[3]_3 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][31] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[3]_3 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][32] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[3]_3 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][33] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[3]_3 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][34] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[3]_3 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][35] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[3]_3 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][36] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[3]_3 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][37] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[3]_3 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][38] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[3]_3 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][39] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[3]_3 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][3] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[3]_3 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][40] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[3]_3 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][41] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[3]_3 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][42] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[3]_3 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][43] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[3]_3 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][44] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[3]_3 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][45] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[3]_3 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][46] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[3]_3 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][47] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[3]_3 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][48] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[3]_3 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][49] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[3]_3 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][4] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[3]_3 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][50] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[3]_3 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][51] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[3]_3 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][52] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[3]_3 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][53] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[3]_3 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][54] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[3]_3 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][55] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[3]_3 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][56] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[3]_3 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][57] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[3]_3 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][58] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[3]_3 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][59] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[3]_3 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][5] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[3]_3 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][60] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[3]_3 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][61] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[3]_3 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][62] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[3]_3 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][63] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[3]_3 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][64] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[3]_3 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][65] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[3]_3 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][66] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[3]_3 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][67] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[3]_3 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][68] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[3]_3 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][69] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[3]_3 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][6] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[3]_3 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][70] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[3]_3 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][71] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[3]_3 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][72] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[3]_3 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][73] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[3]_3 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][74] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[3]_3 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][75] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[3]_3 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][76] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[3]_3 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][77] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[3]_3 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][78] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[3]_3 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][79] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[3]_3 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][7] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[3]_3 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][80] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[3]_3 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][81] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[3]_3 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][82] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[3]_3 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][83] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[3]_3 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][84] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[3]_3 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][85] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[3]_3 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][86] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[3]_3 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][87] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[3]_3 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][88] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[3]_3 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][89] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[3]_3 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][8] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[3]_3 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][90] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[3]_3 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][91] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[3]_3 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][92] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[3]_3 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][93] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[3]_3 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][94] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[3]_3 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][95] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[3]_3 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][96] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[3]_3 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][97] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[3]_3 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][98] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[3]_3 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][99] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[3]_3 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[3][9] 
       (.C(clk_i),
        .CE(\key_mem[3][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[3]_3 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][0] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[4]_4 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][100] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[4]_4 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][101] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[4]_4 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][102] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[4]_4 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][103] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[4]_4 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][104] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[4]_4 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][105] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[4]_4 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][106] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[4]_4 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][107] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[4]_4 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][108] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[4]_4 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][109] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[4]_4 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][10] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[4]_4 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][110] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[4]_4 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][111] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[4]_4 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][112] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[4]_4 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][113] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[4]_4 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][114] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[4]_4 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][115] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[4]_4 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][116] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[4]_4 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][117] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[4]_4 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][118] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[4]_4 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][119] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[4]_4 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][11] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[4]_4 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][120] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[4]_4 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][121] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[4]_4 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][122] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[4]_4 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][123] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[4]_4 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][124] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[4]_4 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][125] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[4]_4 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][126] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[4]_4 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][127] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[4]_4 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][12] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[4]_4 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][13] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[4]_4 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][14] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[4]_4 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][15] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[4]_4 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][16] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[4]_4 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][17] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[4]_4 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][18] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[4]_4 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][19] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[4]_4 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][1] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[4]_4 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][20] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[4]_4 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][21] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[4]_4 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][22] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[4]_4 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][23] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[4]_4 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][24] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[4]_4 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][25] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[4]_4 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][26] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[4]_4 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][27] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[4]_4 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][28] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[4]_4 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][29] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[4]_4 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][2] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[4]_4 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][30] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[4]_4 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][31] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[4]_4 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][32] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[4]_4 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][33] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[4]_4 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][34] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[4]_4 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][35] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[4]_4 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][36] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[4]_4 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][37] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[4]_4 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][38] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[4]_4 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][39] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[4]_4 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][3] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[4]_4 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][40] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[4]_4 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][41] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[4]_4 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][42] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[4]_4 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][43] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[4]_4 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][44] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[4]_4 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][45] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[4]_4 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][46] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[4]_4 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][47] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[4]_4 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][48] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[4]_4 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][49] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[4]_4 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][4] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[4]_4 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][50] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[4]_4 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][51] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[4]_4 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][52] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[4]_4 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][53] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[4]_4 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][54] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[4]_4 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][55] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[4]_4 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][56] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[4]_4 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][57] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[4]_4 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][58] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[4]_4 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][59] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[4]_4 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][5] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[4]_4 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][60] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[4]_4 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][61] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[4]_4 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][62] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[4]_4 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][63] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[4]_4 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][64] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[4]_4 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][65] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[4]_4 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][66] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[4]_4 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][67] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[4]_4 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][68] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[4]_4 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][69] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[4]_4 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][6] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[4]_4 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][70] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[4]_4 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][71] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[4]_4 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][72] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[4]_4 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][73] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[4]_4 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][74] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[4]_4 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][75] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[4]_4 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][76] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[4]_4 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][77] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[4]_4 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][78] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[4]_4 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][79] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[4]_4 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][7] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[4]_4 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][80] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[4]_4 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][81] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[4]_4 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][82] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[4]_4 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][83] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[4]_4 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][84] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[4]_4 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][85] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[4]_4 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][86] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[4]_4 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][87] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[4]_4 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][88] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[4]_4 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][89] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[4]_4 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][8] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[4]_4 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][90] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[4]_4 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][91] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[4]_4 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][92] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[4]_4 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][93] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[4]_4 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][94] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[4]_4 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][95] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[4]_4 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][96] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[4]_4 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][97] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[4]_4 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][98] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[4]_4 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][99] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[4]_4 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[4][9] 
       (.C(clk_i),
        .CE(\key_mem[4][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[4]_4 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][0] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[5]_5 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][100] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[5]_5 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][101] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[5]_5 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][102] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[5]_5 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][103] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[5]_5 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][104] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[5]_5 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][105] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[5]_5 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][106] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[5]_5 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][107] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[5]_5 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][108] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[5]_5 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][109] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[5]_5 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][10] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[5]_5 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][110] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[5]_5 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][111] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[5]_5 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][112] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[5]_5 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][113] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[5]_5 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][114] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[5]_5 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][115] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[5]_5 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][116] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[5]_5 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][117] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[5]_5 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][118] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[5]_5 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][119] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[5]_5 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][11] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[5]_5 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][120] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[5]_5 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][121] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[5]_5 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][122] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[5]_5 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][123] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[5]_5 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][124] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[5]_5 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][125] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[5]_5 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][126] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[5]_5 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][127] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[5]_5 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][12] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[5]_5 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][13] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[5]_5 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][14] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[5]_5 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][15] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[5]_5 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][16] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[5]_5 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][17] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[5]_5 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][18] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[5]_5 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][19] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[5]_5 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][1] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[5]_5 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][20] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[5]_5 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][21] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[5]_5 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][22] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[5]_5 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][23] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[5]_5 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][24] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[5]_5 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][25] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[5]_5 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][26] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[5]_5 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][27] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[5]_5 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][28] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[5]_5 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][29] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[5]_5 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][2] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[5]_5 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][30] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[5]_5 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][31] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[5]_5 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][32] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[5]_5 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][33] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[5]_5 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][34] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[5]_5 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][35] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[5]_5 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][36] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[5]_5 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][37] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[5]_5 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][38] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[5]_5 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][39] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[5]_5 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][3] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[5]_5 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][40] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[5]_5 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][41] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[5]_5 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][42] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[5]_5 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][43] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[5]_5 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][44] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[5]_5 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][45] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[5]_5 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][46] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[5]_5 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][47] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[5]_5 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][48] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[5]_5 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][49] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[5]_5 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][4] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[5]_5 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][50] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[5]_5 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][51] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[5]_5 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][52] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[5]_5 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][53] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[5]_5 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][54] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[5]_5 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][55] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[5]_5 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][56] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[5]_5 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][57] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[5]_5 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][58] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[5]_5 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][59] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[5]_5 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][5] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[5]_5 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][60] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[5]_5 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][61] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[5]_5 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][62] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[5]_5 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][63] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[5]_5 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][64] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[5]_5 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][65] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[5]_5 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][66] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[5]_5 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][67] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[5]_5 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][68] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[5]_5 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][69] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[5]_5 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][6] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[5]_5 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][70] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[5]_5 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][71] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[5]_5 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][72] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[5]_5 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][73] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[5]_5 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][74] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[5]_5 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][75] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[5]_5 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][76] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[5]_5 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][77] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[5]_5 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][78] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[5]_5 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][79] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[5]_5 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][7] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[5]_5 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][80] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[5]_5 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][81] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[5]_5 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][82] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[5]_5 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][83] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[5]_5 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][84] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[5]_5 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][85] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[5]_5 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][86] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[5]_5 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][87] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[5]_5 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][88] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[5]_5 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][89] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[5]_5 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][8] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[5]_5 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][90] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[5]_5 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][91] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[5]_5 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][92] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[5]_5 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][93] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[5]_5 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][94] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[5]_5 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][95] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[5]_5 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][96] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[5]_5 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][97] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[5]_5 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][98] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[5]_5 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][99] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[5]_5 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[5][9] 
       (.C(clk_i),
        .CE(\key_mem[5][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[5]_5 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][0] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[6]_6 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][100] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[6]_6 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][101] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[6]_6 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][102] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[6]_6 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][103] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[6]_6 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][104] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[6]_6 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][105] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[6]_6 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][106] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[6]_6 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][107] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[6]_6 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][108] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[6]_6 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][109] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[6]_6 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][10] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[6]_6 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][110] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[6]_6 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][111] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[6]_6 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][112] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[6]_6 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][113] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[6]_6 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][114] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[6]_6 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][115] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[6]_6 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][116] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[6]_6 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][117] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[6]_6 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][118] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[6]_6 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][119] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[6]_6 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][11] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[6]_6 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][120] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[6]_6 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][121] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[6]_6 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][122] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[6]_6 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][123] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[6]_6 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][124] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[6]_6 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][125] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[6]_6 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][126] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[6]_6 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][127] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[6]_6 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][12] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[6]_6 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][13] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[6]_6 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][14] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[6]_6 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][15] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[6]_6 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][16] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[6]_6 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][17] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[6]_6 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][18] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[6]_6 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][19] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[6]_6 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][1] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[6]_6 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][20] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[6]_6 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][21] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[6]_6 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][22] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[6]_6 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][23] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[6]_6 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][24] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[6]_6 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][25] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[6]_6 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][26] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[6]_6 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][27] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[6]_6 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][28] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[6]_6 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][29] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[6]_6 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][2] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[6]_6 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][30] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[6]_6 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][31] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[6]_6 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][32] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[6]_6 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][33] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[6]_6 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][34] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[6]_6 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][35] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[6]_6 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][36] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[6]_6 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][37] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[6]_6 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][38] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[6]_6 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][39] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[6]_6 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][3] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[6]_6 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][40] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[6]_6 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][41] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[6]_6 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][42] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[6]_6 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][43] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[6]_6 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][44] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[6]_6 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][45] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[6]_6 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][46] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[6]_6 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][47] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[6]_6 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][48] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[6]_6 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][49] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[6]_6 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][4] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[6]_6 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][50] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[6]_6 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][51] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[6]_6 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][52] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[6]_6 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][53] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[6]_6 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][54] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[6]_6 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][55] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[6]_6 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][56] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[6]_6 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][57] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[6]_6 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][58] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[6]_6 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][59] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[6]_6 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][5] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[6]_6 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][60] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[6]_6 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][61] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[6]_6 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][62] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[6]_6 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][63] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[6]_6 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][64] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[6]_6 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][65] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[6]_6 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][66] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[6]_6 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][67] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[6]_6 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][68] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[6]_6 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][69] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[6]_6 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][6] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[6]_6 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][70] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[6]_6 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][71] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[6]_6 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][72] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[6]_6 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][73] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[6]_6 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][74] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[6]_6 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][75] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[6]_6 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][76] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[6]_6 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][77] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[6]_6 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][78] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[6]_6 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][79] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[6]_6 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][7] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[6]_6 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][80] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[6]_6 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][81] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[6]_6 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][82] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[6]_6 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][83] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[6]_6 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][84] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[6]_6 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][85] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[6]_6 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][86] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[6]_6 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][87] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[6]_6 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][88] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[6]_6 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][89] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[6]_6 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][8] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[6]_6 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][90] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[6]_6 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][91] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[6]_6 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][92] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[6]_6 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][93] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[6]_6 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][94] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[6]_6 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][95] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[6]_6 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][96] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[6]_6 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][97] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[6]_6 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][98] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[6]_6 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][99] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[6]_6 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[6][9] 
       (.C(clk_i),
        .CE(\key_mem[6][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[6]_6 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][0] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[7]_7 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][100] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[7]_7 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][101] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[7]_7 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][102] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[7]_7 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][103] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[7]_7 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][104] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[7]_7 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][105] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[7]_7 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][106] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[7]_7 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][107] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[7]_7 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][108] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[7]_7 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][109] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[7]_7 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][10] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[7]_7 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][110] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[7]_7 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][111] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[7]_7 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][112] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[7]_7 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][113] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[7]_7 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][114] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[7]_7 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][115] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[7]_7 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][116] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[7]_7 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][117] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[7]_7 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][118] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[7]_7 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][119] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[7]_7 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][11] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[7]_7 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][120] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[7]_7 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][121] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[7]_7 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][122] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[7]_7 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][123] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[7]_7 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][124] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[7]_7 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][125] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[7]_7 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][126] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[7]_7 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][127] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[7]_7 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][12] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[7]_7 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][13] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[7]_7 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][14] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[7]_7 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][15] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[7]_7 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][16] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[7]_7 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][17] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[7]_7 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][18] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[7]_7 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][19] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[7]_7 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][1] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[7]_7 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][20] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[7]_7 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][21] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[7]_7 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][22] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[7]_7 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][23] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[7]_7 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][24] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[7]_7 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][25] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[7]_7 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][26] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[7]_7 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][27] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[7]_7 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][28] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[7]_7 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][29] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[7]_7 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][2] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[7]_7 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][30] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[7]_7 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][31] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[7]_7 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][32] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[7]_7 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][33] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[7]_7 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][34] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[7]_7 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][35] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[7]_7 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][36] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[7]_7 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][37] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[7]_7 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][38] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[7]_7 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][39] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[7]_7 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][3] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[7]_7 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][40] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[7]_7 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][41] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[7]_7 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][42] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[7]_7 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][43] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[7]_7 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][44] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[7]_7 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][45] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[7]_7 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][46] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[7]_7 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][47] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[7]_7 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][48] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[7]_7 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][49] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[7]_7 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][4] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[7]_7 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][50] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[7]_7 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][51] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[7]_7 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][52] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[7]_7 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][53] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[7]_7 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][54] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[7]_7 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][55] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[7]_7 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][56] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[7]_7 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][57] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[7]_7 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][58] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[7]_7 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][59] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[7]_7 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][5] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[7]_7 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][60] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[7]_7 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][61] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[7]_7 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][62] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[7]_7 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][63] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[7]_7 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][64] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[7]_7 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][65] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[7]_7 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][66] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[7]_7 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][67] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[7]_7 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][68] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[7]_7 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][69] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[7]_7 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][6] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[7]_7 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][70] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[7]_7 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][71] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[7]_7 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][72] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[7]_7 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][73] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[7]_7 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][74] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[7]_7 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][75] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[7]_7 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][76] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[7]_7 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][77] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[7]_7 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][78] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[7]_7 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][79] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[7]_7 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][7] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[7]_7 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][80] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[7]_7 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][81] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[7]_7 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][82] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[7]_7 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][83] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[7]_7 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][84] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[7]_7 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][85] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[7]_7 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][86] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[7]_7 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][87] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[7]_7 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][88] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[7]_7 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][89] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[7]_7 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][8] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[7]_7 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][90] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[7]_7 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][91] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[7]_7 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][92] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[7]_7 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][93] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[7]_7 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][94] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[7]_7 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][95] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[7]_7 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][96] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[7]_7 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][97] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[7]_7 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][98] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[7]_7 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][99] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[7]_7 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[7][9] 
       (.C(clk_i),
        .CE(\key_mem[7][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[7]_7 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][0] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[8]_8 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][100] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[8]_8 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][101] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[8]_8 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][102] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[8]_8 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][103] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[8]_8 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][104] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[8]_8 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][105] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[8]_8 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][106] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[8]_8 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][107] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[8]_8 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][108] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[8]_8 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][109] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[8]_8 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][10] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[8]_8 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][110] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[8]_8 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][111] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[8]_8 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][112] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[8]_8 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][113] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[8]_8 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][114] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[8]_8 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][115] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[8]_8 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][116] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[8]_8 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][117] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[8]_8 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][118] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[8]_8 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][119] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[8]_8 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][11] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[8]_8 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][120] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[8]_8 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][121] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[8]_8 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][122] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[8]_8 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][123] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[8]_8 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][124] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[8]_8 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][125] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[8]_8 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][126] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[8]_8 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][127] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[8]_8 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][12] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[8]_8 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][13] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[8]_8 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][14] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[8]_8 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][15] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[8]_8 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][16] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[8]_8 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][17] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[8]_8 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][18] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[8]_8 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][19] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[8]_8 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][1] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[8]_8 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][20] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[8]_8 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][21] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[8]_8 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][22] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[8]_8 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][23] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[8]_8 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][24] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[8]_8 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][25] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[8]_8 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][26] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[8]_8 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][27] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[8]_8 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][28] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[8]_8 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][29] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[8]_8 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][2] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[8]_8 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][30] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[8]_8 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][31] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[8]_8 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][32] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[8]_8 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][33] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[8]_8 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][34] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[8]_8 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][35] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[8]_8 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][36] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[8]_8 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][37] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[8]_8 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][38] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[8]_8 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][39] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[8]_8 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][3] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[8]_8 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][40] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[8]_8 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][41] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[8]_8 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][42] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[8]_8 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][43] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[8]_8 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][44] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[8]_8 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][45] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[8]_8 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][46] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[8]_8 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][47] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[8]_8 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][48] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[8]_8 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][49] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[8]_8 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][4] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[8]_8 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][50] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[8]_8 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][51] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[8]_8 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][52] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[8]_8 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][53] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[8]_8 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][54] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[8]_8 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][55] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[8]_8 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][56] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[8]_8 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][57] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[8]_8 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][58] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[8]_8 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][59] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[8]_8 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][5] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[8]_8 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][60] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[8]_8 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][61] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[8]_8 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][62] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[8]_8 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][63] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[8]_8 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][64] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[8]_8 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][65] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[8]_8 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][66] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[8]_8 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][67] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[8]_8 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][68] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[8]_8 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][69] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[8]_8 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][6] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[8]_8 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][70] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[8]_8 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][71] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[8]_8 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][72] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[8]_8 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][73] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[8]_8 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][74] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[8]_8 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][75] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[8]_8 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][76] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[8]_8 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][77] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[8]_8 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][78] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[8]_8 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][79] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[8]_8 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][7] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[8]_8 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][80] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[8]_8 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][81] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[8]_8 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][82] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[8]_8 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][83] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[8]_8 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][84] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[8]_8 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][85] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[8]_8 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][86] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[8]_8 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][87] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[8]_8 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][88] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[8]_8 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][89] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[8]_8 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][8] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[8]_8 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][90] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[8]_8 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][91] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[8]_8 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][92] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[8]_8 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][93] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[8]_8 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][94] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[8]_8 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][95] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[8]_8 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][96] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[8]_8 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][97] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[8]_8 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][98] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[8]_8 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][99] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[8]_8 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[8][9] 
       (.C(clk_i),
        .CE(\key_mem[8][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[8]_8 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][0] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[0]),
        .Q(\key_mem_reg[9]_9 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][100] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[100]),
        .Q(\key_mem_reg[9]_9 [100]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][101] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[101]),
        .Q(\key_mem_reg[9]_9 [101]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][102] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[102]),
        .Q(\key_mem_reg[9]_9 [102]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][103] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[103]),
        .Q(\key_mem_reg[9]_9 [103]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][104] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[104]),
        .Q(\key_mem_reg[9]_9 [104]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][105] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[105]),
        .Q(\key_mem_reg[9]_9 [105]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][106] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[106]),
        .Q(\key_mem_reg[9]_9 [106]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][107] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[107]),
        .Q(\key_mem_reg[9]_9 [107]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][108] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[108]),
        .Q(\key_mem_reg[9]_9 [108]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][109] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[109]),
        .Q(\key_mem_reg[9]_9 [109]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][10] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[10]),
        .Q(\key_mem_reg[9]_9 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][110] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[110]),
        .Q(\key_mem_reg[9]_9 [110]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][111] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[111]),
        .Q(\key_mem_reg[9]_9 [111]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][112] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[112]),
        .Q(\key_mem_reg[9]_9 [112]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][113] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[113]),
        .Q(\key_mem_reg[9]_9 [113]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][114] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[114]),
        .Q(\key_mem_reg[9]_9 [114]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][115] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[115]),
        .Q(\key_mem_reg[9]_9 [115]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][116] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[116]),
        .Q(\key_mem_reg[9]_9 [116]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][117] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[117]),
        .Q(\key_mem_reg[9]_9 [117]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][118] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[118]),
        .Q(\key_mem_reg[9]_9 [118]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][119] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[119]),
        .Q(\key_mem_reg[9]_9 [119]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][11] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[11]),
        .Q(\key_mem_reg[9]_9 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][120] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[120]),
        .Q(\key_mem_reg[9]_9 [120]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][121] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[121]),
        .Q(\key_mem_reg[9]_9 [121]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][122] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[122]),
        .Q(\key_mem_reg[9]_9 [122]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][123] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[123]),
        .Q(\key_mem_reg[9]_9 [123]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][124] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[124]),
        .Q(\key_mem_reg[9]_9 [124]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][125] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[125]),
        .Q(\key_mem_reg[9]_9 [125]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][126] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[126]),
        .Q(\key_mem_reg[9]_9 [126]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][127] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[127]),
        .Q(\key_mem_reg[9]_9 [127]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][12] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[12]),
        .Q(\key_mem_reg[9]_9 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][13] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[13]),
        .Q(\key_mem_reg[9]_9 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][14] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[14]),
        .Q(\key_mem_reg[9]_9 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][15] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[15]),
        .Q(\key_mem_reg[9]_9 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][16] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[16]),
        .Q(\key_mem_reg[9]_9 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][17] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[17]),
        .Q(\key_mem_reg[9]_9 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][18] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[18]),
        .Q(\key_mem_reg[9]_9 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][19] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[19]),
        .Q(\key_mem_reg[9]_9 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][1] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[1]),
        .Q(\key_mem_reg[9]_9 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][20] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[20]),
        .Q(\key_mem_reg[9]_9 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][21] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[21]),
        .Q(\key_mem_reg[9]_9 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][22] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[22]),
        .Q(\key_mem_reg[9]_9 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][23] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[23]),
        .Q(\key_mem_reg[9]_9 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][24] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[24]),
        .Q(\key_mem_reg[9]_9 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][25] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[25]),
        .Q(\key_mem_reg[9]_9 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][26] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[26]),
        .Q(\key_mem_reg[9]_9 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][27] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[27]),
        .Q(\key_mem_reg[9]_9 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][28] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[28]),
        .Q(\key_mem_reg[9]_9 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][29] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[29]),
        .Q(\key_mem_reg[9]_9 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][2] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[2]),
        .Q(\key_mem_reg[9]_9 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][30] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[30]),
        .Q(\key_mem_reg[9]_9 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][31] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[31]),
        .Q(\key_mem_reg[9]_9 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][32] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[32]),
        .Q(\key_mem_reg[9]_9 [32]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][33] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[33]),
        .Q(\key_mem_reg[9]_9 [33]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][34] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[34]),
        .Q(\key_mem_reg[9]_9 [34]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][35] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[35]),
        .Q(\key_mem_reg[9]_9 [35]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][36] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[36]),
        .Q(\key_mem_reg[9]_9 [36]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][37] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[37]),
        .Q(\key_mem_reg[9]_9 [37]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][38] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[38]),
        .Q(\key_mem_reg[9]_9 [38]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][39] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[39]),
        .Q(\key_mem_reg[9]_9 [39]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][3] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[3]),
        .Q(\key_mem_reg[9]_9 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][40] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[40]),
        .Q(\key_mem_reg[9]_9 [40]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][41] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[41]),
        .Q(\key_mem_reg[9]_9 [41]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][42] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[42]),
        .Q(\key_mem_reg[9]_9 [42]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][43] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[43]),
        .Q(\key_mem_reg[9]_9 [43]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][44] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[44]),
        .Q(\key_mem_reg[9]_9 [44]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][45] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[45]),
        .Q(\key_mem_reg[9]_9 [45]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][46] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[46]),
        .Q(\key_mem_reg[9]_9 [46]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][47] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[47]),
        .Q(\key_mem_reg[9]_9 [47]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][48] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[48]),
        .Q(\key_mem_reg[9]_9 [48]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][49] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[49]),
        .Q(\key_mem_reg[9]_9 [49]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][4] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[4]),
        .Q(\key_mem_reg[9]_9 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][50] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[50]),
        .Q(\key_mem_reg[9]_9 [50]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][51] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[51]),
        .Q(\key_mem_reg[9]_9 [51]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][52] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[52]),
        .Q(\key_mem_reg[9]_9 [52]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][53] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[53]),
        .Q(\key_mem_reg[9]_9 [53]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][54] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[54]),
        .Q(\key_mem_reg[9]_9 [54]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][55] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[55]),
        .Q(\key_mem_reg[9]_9 [55]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][56] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[56]),
        .Q(\key_mem_reg[9]_9 [56]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][57] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[57]),
        .Q(\key_mem_reg[9]_9 [57]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][58] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[58]),
        .Q(\key_mem_reg[9]_9 [58]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][59] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[59]),
        .Q(\key_mem_reg[9]_9 [59]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][5] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[5]),
        .Q(\key_mem_reg[9]_9 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][60] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[60]),
        .Q(\key_mem_reg[9]_9 [60]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][61] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[61]),
        .Q(\key_mem_reg[9]_9 [61]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][62] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[62]),
        .Q(\key_mem_reg[9]_9 [62]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][63] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[63]),
        .Q(\key_mem_reg[9]_9 [63]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][64] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[64]),
        .Q(\key_mem_reg[9]_9 [64]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][65] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[65]),
        .Q(\key_mem_reg[9]_9 [65]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][66] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[66]),
        .Q(\key_mem_reg[9]_9 [66]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][67] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[67]),
        .Q(\key_mem_reg[9]_9 [67]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][68] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[68]),
        .Q(\key_mem_reg[9]_9 [68]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][69] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[69]),
        .Q(\key_mem_reg[9]_9 [69]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][6] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[6]),
        .Q(\key_mem_reg[9]_9 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][70] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[70]),
        .Q(\key_mem_reg[9]_9 [70]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][71] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[71]),
        .Q(\key_mem_reg[9]_9 [71]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][72] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[72]),
        .Q(\key_mem_reg[9]_9 [72]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][73] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[73]),
        .Q(\key_mem_reg[9]_9 [73]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][74] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[74]),
        .Q(\key_mem_reg[9]_9 [74]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][75] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[75]),
        .Q(\key_mem_reg[9]_9 [75]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][76] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[76]),
        .Q(\key_mem_reg[9]_9 [76]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][77] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[77]),
        .Q(\key_mem_reg[9]_9 [77]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][78] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[78]),
        .Q(\key_mem_reg[9]_9 [78]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][79] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[79]),
        .Q(\key_mem_reg[9]_9 [79]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][7] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[7]),
        .Q(\key_mem_reg[9]_9 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][80] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[80]),
        .Q(\key_mem_reg[9]_9 [80]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][81] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[81]),
        .Q(\key_mem_reg[9]_9 [81]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][82] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[82]),
        .Q(\key_mem_reg[9]_9 [82]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][83] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[83]),
        .Q(\key_mem_reg[9]_9 [83]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][84] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[84]),
        .Q(\key_mem_reg[9]_9 [84]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][85] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[85]),
        .Q(\key_mem_reg[9]_9 [85]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][86] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[86]),
        .Q(\key_mem_reg[9]_9 [86]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][87] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[87]),
        .Q(\key_mem_reg[9]_9 [87]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][88] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[88]),
        .Q(\key_mem_reg[9]_9 [88]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][89] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[89]),
        .Q(\key_mem_reg[9]_9 [89]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][8] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[8]),
        .Q(\key_mem_reg[9]_9 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][90] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[90]),
        .Q(\key_mem_reg[9]_9 [90]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][91] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[91]),
        .Q(\key_mem_reg[9]_9 [91]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][92] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[92]),
        .Q(\key_mem_reg[9]_9 [92]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][93] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[93]),
        .Q(\key_mem_reg[9]_9 [93]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][94] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[94]),
        .Q(\key_mem_reg[9]_9 [94]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][95] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[95]),
        .Q(\key_mem_reg[9]_9 [95]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][96] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[96]),
        .Q(\key_mem_reg[9]_9 [96]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][97] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[97]),
        .Q(\key_mem_reg[9]_9 [97]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][98] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[98]),
        .Q(\key_mem_reg[9]_9 [98]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][99] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[99]),
        .Q(\key_mem_reg[9]_9 [99]));
  FDCE #(
    .INIT(1'b0)) 
    \key_mem_reg[9][9] 
       (.C(clk_i),
        .CE(\key_mem[9][127]_i_1_n_0 ),
        .CLR(rst_i),
        .D(key_mem_new[9]),
        .Q(\key_mem_reg[9]_9 [9]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[0]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[0]),
        .I4(core_key[128]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[0]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[100]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[4]),
        .I4(core_key[228]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[100]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[101]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[5]),
        .I4(core_key[229]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[101]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[102]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[6]),
        .I4(core_key[230]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[102]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[103]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[7]),
        .I4(core_key[231]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[103]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[104]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[8]),
        .I4(core_key[232]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[104]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[105]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[9]),
        .I4(core_key[233]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[105]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[106]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[10]),
        .I4(core_key[234]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[106]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[107]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[11]),
        .I4(core_key[235]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[107]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[108]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[12]),
        .I4(core_key[236]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[108]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[109]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[13]),
        .I4(core_key[237]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[109]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[10]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[10]),
        .I4(core_key[138]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[10]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[110]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[14]),
        .I4(core_key[238]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[110]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[111]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[15]),
        .I4(core_key[239]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[111]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[112]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[16]),
        .I4(core_key[240]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[112]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[113]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[17]),
        .I4(core_key[241]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[113]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[114]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[18]),
        .I4(core_key[242]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[114]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[115]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[19]),
        .I4(core_key[243]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[115]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[116]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[20]),
        .I4(core_key[244]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[116]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[117]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[21]),
        .I4(core_key[245]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[117]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[118]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[22]),
        .I4(core_key[246]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[118]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[119]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[23]),
        .I4(core_key[247]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[119]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[11]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[11]),
        .I4(core_key[139]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[11]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[120]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[24]),
        .I4(core_key[248]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[120]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[121]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[25]),
        .I4(core_key[249]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[121]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[122]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[26]),
        .I4(core_key[250]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[122]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[123]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[27]),
        .I4(core_key[251]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[123]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[124]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[28]),
        .I4(core_key[252]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[124]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[125]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[29]),
        .I4(core_key[253]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[125]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[126]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[30]),
        .I4(core_key[254]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[126]));
  LUT3 #(
    .INIT(8'h20)) 
    \prev_key0_reg[127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(p_1_in[2]),
        .O(prev_key0_we2_out));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[127]_i_2 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[31]),
        .I4(core_key[255]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[127]));
  LUT4 #(
    .INIT(16'h0010)) 
    \prev_key0_reg[127]_i_3 
       (.I0(\round_ctr_reg_reg_n_0_[2] ),
        .I1(\round_ctr_reg_reg_n_0_[3] ),
        .I2(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I3(p_0_in0),
        .O(\prev_key0_reg[127]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[12]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[12]),
        .I4(core_key[140]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[12]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[13]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[13]),
        .I4(core_key[141]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[13]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[14]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[14]),
        .I4(core_key[142]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[14]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[15]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[15]),
        .I4(core_key[143]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[15]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[16]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[16]),
        .I4(core_key[144]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[16]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[17]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[17]),
        .I4(core_key[145]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[17]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[18]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[18]),
        .I4(core_key[146]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[18]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[19]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[19]),
        .I4(core_key[147]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[19]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[1]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[1]),
        .I4(core_key[129]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[1]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[20]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[20]),
        .I4(core_key[148]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[20]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[21]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[21]),
        .I4(core_key[149]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[21]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[22]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[22]),
        .I4(core_key[150]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[22]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[23]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[23]),
        .I4(core_key[151]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[23]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[24]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[24]),
        .I4(core_key[152]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[24]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[25]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[25]),
        .I4(core_key[153]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[25]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[26]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[26]),
        .I4(core_key[154]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[26]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[27]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[27]),
        .I4(core_key[155]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[27]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[28]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[28]),
        .I4(core_key[156]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[28]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[29]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[29]),
        .I4(core_key[157]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[29]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[2]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[2]),
        .I4(core_key[130]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[2]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[30]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[30]),
        .I4(core_key[158]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[30]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[31]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[31]),
        .I4(core_key[159]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[31]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[32]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[0]),
        .I4(core_key[160]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[32]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[33]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[1]),
        .I4(core_key[161]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[33]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[34]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[2]),
        .I4(core_key[162]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[34]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[35]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[3]),
        .I4(core_key[163]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[35]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[36]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[4]),
        .I4(core_key[164]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[36]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[37]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[5]),
        .I4(core_key[165]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[37]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[38]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[6]),
        .I4(core_key[166]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[38]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[39]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[7]),
        .I4(core_key[167]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[39]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[3]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[3]),
        .I4(core_key[131]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[3]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[40]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[8]),
        .I4(core_key[168]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[40]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[41]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[9]),
        .I4(core_key[169]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[41]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[42]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[10]),
        .I4(core_key[170]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[42]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[43]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[11]),
        .I4(core_key[171]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[43]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[44]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[12]),
        .I4(core_key[172]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[44]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[45]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[13]),
        .I4(core_key[173]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[45]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[46]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[14]),
        .I4(core_key[174]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[46]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[47]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[15]),
        .I4(core_key[175]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[47]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[48]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[16]),
        .I4(core_key[176]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[48]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[49]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[17]),
        .I4(core_key[177]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[49]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[4]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[4]),
        .I4(core_key[132]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[4]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[50]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[18]),
        .I4(core_key[178]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[50]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[51]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[19]),
        .I4(core_key[179]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[51]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[52]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[20]),
        .I4(core_key[180]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[52]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[53]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[21]),
        .I4(core_key[181]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[53]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[54]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[22]),
        .I4(core_key[182]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[54]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[55]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[23]),
        .I4(core_key[183]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[55]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[56]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[24]),
        .I4(core_key[184]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[56]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[57]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[25]),
        .I4(core_key[185]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[57]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[58]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[26]),
        .I4(core_key[186]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[58]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[59]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[27]),
        .I4(core_key[187]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[59]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[5]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[5]),
        .I4(core_key[133]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[5]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[60]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[28]),
        .I4(core_key[188]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[60]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[61]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[29]),
        .I4(core_key[189]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[61]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[62]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[30]),
        .I4(core_key[190]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[62]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[63]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w6[31]),
        .I4(core_key[191]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[63]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[64]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[0]),
        .I4(core_key[192]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[64]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[65]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[1]),
        .I4(core_key[193]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[65]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[66]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[2]),
        .I4(core_key[194]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[66]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[67]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[3]),
        .I4(core_key[195]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[67]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[68]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[4]),
        .I4(core_key[196]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[68]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[69]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[5]),
        .I4(core_key[197]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[69]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[6]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[6]),
        .I4(core_key[134]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[6]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[70]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[6]),
        .I4(core_key[198]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[70]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[71]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[7]),
        .I4(core_key[199]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[71]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[72]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[8]),
        .I4(core_key[200]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[72]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[73]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[9]),
        .I4(core_key[201]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[73]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[74]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[10]),
        .I4(core_key[202]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[74]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[75]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[11]),
        .I4(core_key[203]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[75]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[76]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[12]),
        .I4(core_key[204]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[76]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[77]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[13]),
        .I4(core_key[205]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[77]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[78]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[14]),
        .I4(core_key[206]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[78]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[79]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[15]),
        .I4(core_key[207]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[79]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[7]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[7]),
        .I4(core_key[135]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[7]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[80]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[16]),
        .I4(core_key[208]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[80]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[81]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[17]),
        .I4(core_key[209]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[81]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[82]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[18]),
        .I4(core_key[210]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[82]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[83]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[19]),
        .I4(core_key[211]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[83]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[84]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[20]),
        .I4(core_key[212]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[84]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[85]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[21]),
        .I4(core_key[213]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[85]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[86]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[22]),
        .I4(core_key[214]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[86]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[87]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[23]),
        .I4(core_key[215]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[87]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[88]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[24]),
        .I4(core_key[216]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[88]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[89]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[25]),
        .I4(core_key[217]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[89]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[8]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[8]),
        .I4(core_key[136]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[8]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[90]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[26]),
        .I4(core_key[218]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[90]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[91]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[27]),
        .I4(core_key[219]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[91]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[92]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[28]),
        .I4(core_key[220]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[92]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[93]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[29]),
        .I4(core_key[221]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[93]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[94]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[30]),
        .I4(core_key[222]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[94]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[95]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w5[31]),
        .I4(core_key[223]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[95]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[96]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[0]),
        .I4(core_key[224]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[96]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[97]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[1]),
        .I4(core_key[225]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[97]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[98]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[2]),
        .I4(core_key[226]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[98]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[99]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(w4[3]),
        .I4(core_key[227]),
        .I5(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .O(prev_key0_new[99]));
  LUT6 #(
    .INIT(64'hFE00FE00FF01FE00)) 
    \prev_key0_reg[9]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[3] ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(p_0_in0),
        .I3(Q[9]),
        .I4(core_key[137]),
        .I5(\round_ctr_reg_reg[0]_rep_n_0 ),
        .O(prev_key0_new[9]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[0] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[0]),
        .Q(\prev_key0_reg_reg_n_0_[0] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[100] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[100]),
        .Q(w0[4]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[101] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[101]),
        .Q(w0[5]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[102] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[102]),
        .Q(w0[6]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[103] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[103]),
        .Q(w0[7]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[104] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[104]),
        .Q(w0[8]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[105] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[105]),
        .Q(w0[9]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[106] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[106]),
        .Q(w0[10]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[107] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[107]),
        .Q(w0[11]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[108] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[108]),
        .Q(w0[12]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[109] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[109]),
        .Q(w0[13]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[10] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[10]),
        .Q(\prev_key0_reg_reg_n_0_[10] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[110] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[110]),
        .Q(w0[14]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[111] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[111]),
        .Q(w0[15]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[112] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[112]),
        .Q(w0[16]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[113] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[113]),
        .Q(w0[17]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[114] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[114]),
        .Q(w0[18]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[115] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[115]),
        .Q(w0[19]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[116] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[116]),
        .Q(w0[20]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[117] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[117]),
        .Q(w0[21]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[118] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[118]),
        .Q(w0[22]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[119] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[119]),
        .Q(w0[23]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[11] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[11]),
        .Q(\prev_key0_reg_reg_n_0_[11] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[120] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[120]),
        .Q(w0[24]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[121] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[121]),
        .Q(w0[25]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[122] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[122]),
        .Q(w0[26]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[123] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[123]),
        .Q(w0[27]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[124] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[124]),
        .Q(w0[28]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[125] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[125]),
        .Q(w0[29]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[126] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[126]),
        .Q(w0[30]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[127] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[127]),
        .Q(w0[31]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[12] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[12]),
        .Q(\prev_key0_reg_reg_n_0_[12] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[13] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[13]),
        .Q(\prev_key0_reg_reg_n_0_[13] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[14] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[14]),
        .Q(\prev_key0_reg_reg_n_0_[14] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[15] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[15]),
        .Q(\prev_key0_reg_reg_n_0_[15] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[16] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[16]),
        .Q(\prev_key0_reg_reg_n_0_[16] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[17] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[17]),
        .Q(\prev_key0_reg_reg_n_0_[17] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[18] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[18]),
        .Q(\prev_key0_reg_reg_n_0_[18] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[19] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[19]),
        .Q(\prev_key0_reg_reg_n_0_[19] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[1] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[1]),
        .Q(\prev_key0_reg_reg_n_0_[1] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[20] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[20]),
        .Q(\prev_key0_reg_reg_n_0_[20] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[21] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[21]),
        .Q(\prev_key0_reg_reg_n_0_[21] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[22] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[22]),
        .Q(\prev_key0_reg_reg_n_0_[22] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[23] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[23]),
        .Q(\prev_key0_reg_reg_n_0_[23] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[24] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[24]),
        .Q(\prev_key0_reg_reg_n_0_[24] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[25] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[25]),
        .Q(\prev_key0_reg_reg_n_0_[25] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[26] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[26]),
        .Q(\prev_key0_reg_reg_n_0_[26] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[27] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[27]),
        .Q(\prev_key0_reg_reg_n_0_[27] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[28] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[28]),
        .Q(\prev_key0_reg_reg_n_0_[28] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[29] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[29]),
        .Q(\prev_key0_reg_reg_n_0_[29] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[2] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[2]),
        .Q(\prev_key0_reg_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[30] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[30]),
        .Q(\prev_key0_reg_reg_n_0_[30] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[31] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[31]),
        .Q(\prev_key0_reg_reg_n_0_[31] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[32] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[32]),
        .Q(w2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[33] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[33]),
        .Q(w2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[34] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[34]),
        .Q(w2[2]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[35] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[35]),
        .Q(w2[3]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[36] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[36]),
        .Q(w2[4]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[37] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[37]),
        .Q(w2[5]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[38] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[38]),
        .Q(w2[6]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[39] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[39]),
        .Q(w2[7]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[3] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[3]),
        .Q(\prev_key0_reg_reg_n_0_[3] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[40] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[40]),
        .Q(w2[8]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[41] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[41]),
        .Q(w2[9]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[42] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[42]),
        .Q(w2[10]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[43] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[43]),
        .Q(w2[11]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[44] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[44]),
        .Q(w2[12]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[45] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[45]),
        .Q(w2[13]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[46] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[46]),
        .Q(w2[14]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[47] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[47]),
        .Q(w2[15]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[48] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[48]),
        .Q(w2[16]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[49] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[49]),
        .Q(w2[17]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[4] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[4]),
        .Q(\prev_key0_reg_reg_n_0_[4] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[50] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[50]),
        .Q(w2[18]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[51] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[51]),
        .Q(w2[19]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[52] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[52]),
        .Q(w2[20]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[53] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[53]),
        .Q(w2[21]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[54] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[54]),
        .Q(w2[22]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[55] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[55]),
        .Q(w2[23]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[56] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[56]),
        .Q(w2[24]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[57] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[57]),
        .Q(w2[25]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[58] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[58]),
        .Q(w2[26]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[59] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[59]),
        .Q(w2[27]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[5] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[5]),
        .Q(\prev_key0_reg_reg_n_0_[5] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[60] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[60]),
        .Q(w2[28]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[61] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[61]),
        .Q(w2[29]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[62] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[62]),
        .Q(w2[30]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[63] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[63]),
        .Q(w2[31]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[64] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[64]),
        .Q(w1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[65] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[65]),
        .Q(w1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[66] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[66]),
        .Q(w1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[67] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[67]),
        .Q(w1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[68] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[68]),
        .Q(w1[4]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[69] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[69]),
        .Q(w1[5]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[6] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[6]),
        .Q(\prev_key0_reg_reg_n_0_[6] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[70] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[70]),
        .Q(w1[6]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[71] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[71]),
        .Q(w1[7]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[72] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[72]),
        .Q(w1[8]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[73] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[73]),
        .Q(w1[9]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[74] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[74]),
        .Q(w1[10]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[75] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[75]),
        .Q(w1[11]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[76] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[76]),
        .Q(w1[12]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[77] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[77]),
        .Q(w1[13]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[78] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[78]),
        .Q(w1[14]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[79] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[79]),
        .Q(w1[15]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[7] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[7]),
        .Q(\prev_key0_reg_reg_n_0_[7] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[80] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[80]),
        .Q(w1[16]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[81] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[81]),
        .Q(w1[17]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[82] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[82]),
        .Q(w1[18]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[83] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[83]),
        .Q(w1[19]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[84] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[84]),
        .Q(w1[20]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[85] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[85]),
        .Q(w1[21]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[86] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[86]),
        .Q(w1[22]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[87] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[87]),
        .Q(w1[23]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[88] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[88]),
        .Q(w1[24]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[89] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[89]),
        .Q(w1[25]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[8] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[8]),
        .Q(\prev_key0_reg_reg_n_0_[8] ));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[90] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[90]),
        .Q(w1[26]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[91] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[91]),
        .Q(w1[27]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[92] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[92]),
        .Q(w1[28]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[93] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[93]),
        .Q(w1[29]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[94] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[94]),
        .Q(w1[30]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[95] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[95]),
        .Q(w1[31]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[96] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[96]),
        .Q(w0[0]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[97] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[97]),
        .Q(w0[1]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[98] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[98]),
        .Q(w0[2]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[99] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[99]),
        .Q(w0[3]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key0_reg_reg[9] 
       (.C(clk_i),
        .CE(prev_key0_we2_out),
        .CLR(rst_i),
        .D(prev_key0_new[9]),
        .Q(\prev_key0_reg_reg_n_0_[9] ));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[0]_i_1 
       (.I0(prev_key1_new0_in[0]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[0]),
        .O(\prev_key1_reg[0]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[0]_i_2 
       (.I0(core_key[128]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[24]),
        .I3(Q[0]),
        .I4(\prev_key1_reg[0]_i_4_n_0 ),
        .O(prev_key1_new0_in[0]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[0]_i_3 
       (.I0(core_key[0]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[0]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[0]),
        .I5(new_sboxw[24]),
        .O(prev_key1_new[0]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[0]_i_4 
       (.I0(w5[0]),
        .I1(w4[0]),
        .I2(w6[0]),
        .O(\prev_key1_reg[0]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[0]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[0] ),
        .I1(w1[0]),
        .I2(w2[0]),
        .I3(w0[0]),
        .O(p_2_in[0]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[100]_i_1 
       (.I0(prev_key1_new0_in[100]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[100]),
        .O(\prev_key1_reg[100]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[100]_i_2 
       (.I0(core_key[228]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[28]),
        .I3(w4[4]),
        .O(prev_key1_new0_in[100]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[100]_i_3 
       (.I0(core_key[100]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[4]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[4]),
        .I5(new_sboxw[28]),
        .O(prev_key1_new[100]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[101]_i_1 
       (.I0(prev_key1_new0_in[101]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[101]),
        .O(\prev_key1_reg[101]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[101]_i_2 
       (.I0(core_key[229]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[29]),
        .I3(w4[5]),
        .O(prev_key1_new0_in[101]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[101]_i_3 
       (.I0(core_key[101]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[5]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[5]),
        .I5(new_sboxw[29]),
        .O(prev_key1_new[101]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[102]_i_1 
       (.I0(prev_key1_new0_in[102]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[102]),
        .O(\prev_key1_reg[102]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[102]_i_2 
       (.I0(core_key[230]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[30]),
        .I3(w4[6]),
        .O(prev_key1_new0_in[102]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[102]_i_3 
       (.I0(core_key[102]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[6]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[6]),
        .I5(new_sboxw[30]),
        .O(prev_key1_new[102]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[103]_i_1 
       (.I0(prev_key1_new0_in[103]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[103]),
        .O(\prev_key1_reg[103]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[103]_i_2 
       (.I0(core_key[231]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[31]),
        .I3(w4[7]),
        .O(prev_key1_new0_in[103]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[103]_i_3 
       (.I0(core_key[103]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[7]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[7]),
        .I5(new_sboxw[31]),
        .O(prev_key1_new[103]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[104]_i_1 
       (.I0(prev_key1_new0_in[104]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[104]),
        .O(\prev_key1_reg[104]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[104]_i_2 
       (.I0(core_key[232]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[0]),
        .I3(w4[8]),
        .O(prev_key1_new0_in[104]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[104]_i_3 
       (.I0(core_key[104]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[8]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[8]),
        .I5(new_sboxw[0]),
        .O(prev_key1_new[104]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[105]_i_1 
       (.I0(prev_key1_new0_in[105]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[105]),
        .O(\prev_key1_reg[105]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[105]_i_2 
       (.I0(core_key[233]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[1]),
        .I3(w4[9]),
        .O(prev_key1_new0_in[105]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[105]_i_3 
       (.I0(core_key[105]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[9]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[9]),
        .I5(new_sboxw[1]),
        .O(prev_key1_new[105]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[106]_i_1 
       (.I0(prev_key1_new0_in[106]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[106]),
        .O(\prev_key1_reg[106]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[106]_i_2 
       (.I0(core_key[234]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[2]),
        .I3(w4[10]),
        .O(prev_key1_new0_in[106]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[106]_i_3 
       (.I0(core_key[106]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[10]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[10]),
        .I5(new_sboxw[2]),
        .O(prev_key1_new[106]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[107]_i_1 
       (.I0(prev_key1_new0_in[107]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[107]),
        .O(\prev_key1_reg[107]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[107]_i_2 
       (.I0(core_key[235]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[3]),
        .I3(w4[11]),
        .O(prev_key1_new0_in[107]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[107]_i_3 
       (.I0(core_key[107]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[11]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[11]),
        .I5(new_sboxw[3]),
        .O(prev_key1_new[107]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[108]_i_1 
       (.I0(prev_key1_new0_in[108]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[108]),
        .O(\prev_key1_reg[108]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[108]_i_2 
       (.I0(core_key[236]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[4]),
        .I3(w4[12]),
        .O(prev_key1_new0_in[108]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[108]_i_3 
       (.I0(core_key[108]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[12]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[12]),
        .I5(new_sboxw[4]),
        .O(prev_key1_new[108]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[109]_i_1 
       (.I0(prev_key1_new0_in[109]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[109]),
        .O(\prev_key1_reg[109]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[109]_i_2 
       (.I0(core_key[237]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[5]),
        .I3(w4[13]),
        .O(prev_key1_new0_in[109]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[109]_i_3 
       (.I0(core_key[109]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[13]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[13]),
        .I5(new_sboxw[5]),
        .O(prev_key1_new[109]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[10]_i_1 
       (.I0(prev_key1_new0_in[10]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[10]),
        .O(\prev_key1_reg[10]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[10]_i_2 
       (.I0(core_key[138]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[2]),
        .I3(Q[10]),
        .I4(\prev_key1_reg[10]_i_4_n_0 ),
        .O(prev_key1_new0_in[10]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[10]_i_3 
       (.I0(core_key[10]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[10]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[10]),
        .I5(new_sboxw[2]),
        .O(prev_key1_new[10]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[10]_i_4 
       (.I0(w5[10]),
        .I1(w4[10]),
        .I2(w6[10]),
        .O(\prev_key1_reg[10]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[10]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[10] ),
        .I1(w1[10]),
        .I2(w2[10]),
        .I3(w0[10]),
        .O(p_2_in[10]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[110]_i_1 
       (.I0(prev_key1_new0_in[110]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[110]),
        .O(\prev_key1_reg[110]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[110]_i_2 
       (.I0(core_key[238]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[6]),
        .I3(w4[14]),
        .O(prev_key1_new0_in[110]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[110]_i_3 
       (.I0(core_key[110]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[14]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[14]),
        .I5(new_sboxw[6]),
        .O(prev_key1_new[110]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[111]_i_1 
       (.I0(prev_key1_new0_in[111]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[111]),
        .O(\prev_key1_reg[111]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[111]_i_2 
       (.I0(core_key[239]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[7]),
        .I3(w4[15]),
        .O(prev_key1_new0_in[111]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[111]_i_3 
       (.I0(core_key[111]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[15]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[15]),
        .I5(new_sboxw[7]),
        .O(prev_key1_new[111]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[112]_i_1 
       (.I0(prev_key1_new0_in[112]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[112]),
        .O(\prev_key1_reg[112]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[112]_i_2 
       (.I0(core_key[240]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[8]),
        .I3(w4[16]),
        .O(prev_key1_new0_in[112]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[112]_i_3 
       (.I0(core_key[112]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[16]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[16]),
        .I5(new_sboxw[8]),
        .O(prev_key1_new[112]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[113]_i_1 
       (.I0(prev_key1_new0_in[113]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[113]),
        .O(\prev_key1_reg[113]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[113]_i_2 
       (.I0(core_key[241]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[9]),
        .I3(w4[17]),
        .O(prev_key1_new0_in[113]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[113]_i_3 
       (.I0(core_key[113]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[17]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[17]),
        .I5(new_sboxw[9]),
        .O(prev_key1_new[113]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[114]_i_1 
       (.I0(prev_key1_new0_in[114]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[114]),
        .O(\prev_key1_reg[114]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[114]_i_2 
       (.I0(core_key[242]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[10]),
        .I3(w4[18]),
        .O(prev_key1_new0_in[114]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[114]_i_3 
       (.I0(core_key[114]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[18]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[18]),
        .I5(new_sboxw[10]),
        .O(prev_key1_new[114]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[115]_i_1 
       (.I0(prev_key1_new0_in[115]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[115]),
        .O(\prev_key1_reg[115]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[115]_i_2 
       (.I0(core_key[243]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[11]),
        .I3(w4[19]),
        .O(prev_key1_new0_in[115]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[115]_i_3 
       (.I0(core_key[115]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[19]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[19]),
        .I5(new_sboxw[11]),
        .O(prev_key1_new[115]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[116]_i_1 
       (.I0(prev_key1_new0_in[116]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[116]),
        .O(\prev_key1_reg[116]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[116]_i_2 
       (.I0(core_key[244]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[12]),
        .I3(w4[20]),
        .O(prev_key1_new0_in[116]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[116]_i_3 
       (.I0(core_key[116]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[20]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[20]),
        .I5(new_sboxw[12]),
        .O(prev_key1_new[116]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[117]_i_1 
       (.I0(prev_key1_new0_in[117]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[117]),
        .O(\prev_key1_reg[117]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[117]_i_2 
       (.I0(core_key[245]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[13]),
        .I3(w4[21]),
        .O(prev_key1_new0_in[117]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[117]_i_3 
       (.I0(core_key[117]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[21]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[21]),
        .I5(new_sboxw[13]),
        .O(prev_key1_new[117]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[118]_i_1 
       (.I0(prev_key1_new0_in[118]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[118]),
        .O(\prev_key1_reg[118]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[118]_i_2 
       (.I0(core_key[246]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[14]),
        .I3(w4[22]),
        .O(prev_key1_new0_in[118]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[118]_i_3 
       (.I0(core_key[118]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[22]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[22]),
        .I5(new_sboxw[14]),
        .O(prev_key1_new[118]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[119]_i_1 
       (.I0(prev_key1_new0_in[119]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[119]),
        .O(\prev_key1_reg[119]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[119]_i_2 
       (.I0(core_key[247]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[15]),
        .I3(w4[23]),
        .O(prev_key1_new0_in[119]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[119]_i_3 
       (.I0(core_key[119]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[23]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[23]),
        .I5(new_sboxw[15]),
        .O(prev_key1_new[119]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[11]_i_1 
       (.I0(prev_key1_new0_in[11]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[11]),
        .O(\prev_key1_reg[11]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[11]_i_2 
       (.I0(core_key[139]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[3]),
        .I3(Q[11]),
        .I4(\prev_key1_reg[11]_i_4_n_0 ),
        .O(prev_key1_new0_in[11]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[11]_i_3 
       (.I0(core_key[11]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[11]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[11]),
        .I5(new_sboxw[3]),
        .O(prev_key1_new[11]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[11]_i_4 
       (.I0(w5[11]),
        .I1(w4[11]),
        .I2(w6[11]),
        .O(\prev_key1_reg[11]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[11]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[11] ),
        .I1(w1[11]),
        .I2(w2[11]),
        .I3(w0[11]),
        .O(p_2_in[11]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[120]_i_1 
       (.I0(prev_key1_new0_in[120]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[120]),
        .O(\prev_key1_reg[120]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[120]_i_2 
       (.I0(core_key[248]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [0]),
        .I3(new_sboxw[16]),
        .I4(w4[24]),
        .O(prev_key1_new0_in[120]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[120]_i_3 
       (.I0(core_key[120]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[24]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[24]),
        .I5(p_19_in[0]),
        .O(prev_key1_new[120]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[121]_i_1 
       (.I0(prev_key1_new0_in[121]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[121]),
        .O(\prev_key1_reg[121]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[121]_i_2 
       (.I0(core_key[249]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [1]),
        .I3(new_sboxw[17]),
        .I4(w4[25]),
        .O(prev_key1_new0_in[121]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[121]_i_3 
       (.I0(core_key[121]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[25]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[25]),
        .I5(p_19_in[1]),
        .O(prev_key1_new[121]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[122]_i_1 
       (.I0(prev_key1_new0_in[122]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[122]),
        .O(\prev_key1_reg[122]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[122]_i_2 
       (.I0(core_key[250]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [2]),
        .I3(new_sboxw[18]),
        .I4(w4[26]),
        .O(prev_key1_new0_in[122]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[122]_i_3 
       (.I0(core_key[122]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[26]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[26]),
        .I5(p_19_in[2]),
        .O(prev_key1_new[122]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[123]_i_1 
       (.I0(prev_key1_new0_in[123]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[123]),
        .O(\prev_key1_reg[123]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[123]_i_2 
       (.I0(core_key[251]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [3]),
        .I3(new_sboxw[19]),
        .I4(w4[27]),
        .O(prev_key1_new0_in[123]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[123]_i_3 
       (.I0(core_key[123]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[27]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[27]),
        .I5(p_19_in[3]),
        .O(prev_key1_new[123]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[124]_i_1 
       (.I0(prev_key1_new0_in[124]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[124]),
        .O(\prev_key1_reg[124]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[124]_i_2 
       (.I0(core_key[252]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [4]),
        .I3(new_sboxw[20]),
        .I4(w4[28]),
        .O(prev_key1_new0_in[124]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[124]_i_3 
       (.I0(core_key[124]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[28]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[28]),
        .I5(p_19_in[4]),
        .O(prev_key1_new[124]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[125]_i_1 
       (.I0(prev_key1_new0_in[125]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[125]),
        .O(\prev_key1_reg[125]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[125]_i_2 
       (.I0(core_key[253]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [5]),
        .I3(new_sboxw[21]),
        .I4(w4[29]),
        .O(prev_key1_new0_in[125]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[125]_i_3 
       (.I0(core_key[125]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[29]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[29]),
        .I5(p_19_in[5]),
        .O(prev_key1_new[125]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[126]_i_1 
       (.I0(prev_key1_new0_in[126]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[126]),
        .O(\prev_key1_reg[126]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[126]_i_2 
       (.I0(core_key[254]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [6]),
        .I3(new_sboxw[22]),
        .I4(w4[30]),
        .O(prev_key1_new0_in[126]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[126]_i_3 
       (.I0(core_key[126]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[30]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[30]),
        .I5(p_19_in[6]),
        .O(prev_key1_new[126]));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \prev_key1_reg[127]_i_1 
       (.I0(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I1(\round_ctr_reg_reg_n_0_[2] ),
        .I2(\round_ctr_reg_reg_n_0_[3] ),
        .I3(\round_ctr_reg_reg[0]_rep_n_0 ),
        .I4(p_1_in[2]),
        .I5(p_0_in0),
        .O(prev_key1_we1_out));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[127]_i_2 
       (.I0(prev_key1_new0_in[127]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[127]),
        .O(\prev_key1_reg[127]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[127]_i_3 
       (.I0(core_key[255]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [7]),
        .I3(new_sboxw[23]),
        .I4(w4[31]),
        .O(prev_key1_new0_in[127]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \prev_key1_reg[127]_i_4 
       (.I0(\round_ctr_reg_reg[0]_rep_n_0 ),
        .I1(p_0_in0),
        .I2(\round_ctr_reg_reg_n_0_[2] ),
        .I3(\round_ctr_reg_reg_n_0_[3] ),
        .O(\prev_key1_reg[127]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[127]_i_5 
       (.I0(core_key[127]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[31]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[31]),
        .I5(p_19_in[7]),
        .O(prev_key1_new[127]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[12]_i_1 
       (.I0(prev_key1_new0_in[12]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[12]),
        .O(\prev_key1_reg[12]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[12]_i_2 
       (.I0(core_key[140]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[4]),
        .I3(Q[12]),
        .I4(\prev_key1_reg[12]_i_4_n_0 ),
        .O(prev_key1_new0_in[12]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[12]_i_3 
       (.I0(core_key[12]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[12]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[12]),
        .I5(new_sboxw[4]),
        .O(prev_key1_new[12]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[12]_i_4 
       (.I0(w5[12]),
        .I1(w4[12]),
        .I2(w6[12]),
        .O(\prev_key1_reg[12]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[12]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[12] ),
        .I1(w1[12]),
        .I2(w2[12]),
        .I3(w0[12]),
        .O(p_2_in[12]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[13]_i_1 
       (.I0(prev_key1_new0_in[13]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[13]),
        .O(\prev_key1_reg[13]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[13]_i_2 
       (.I0(core_key[141]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[5]),
        .I3(Q[13]),
        .I4(\prev_key1_reg[13]_i_4_n_0 ),
        .O(prev_key1_new0_in[13]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[13]_i_3 
       (.I0(core_key[13]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[13]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[13]),
        .I5(new_sboxw[5]),
        .O(prev_key1_new[13]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[13]_i_4 
       (.I0(w5[13]),
        .I1(w4[13]),
        .I2(w6[13]),
        .O(\prev_key1_reg[13]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[13]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[13] ),
        .I1(w1[13]),
        .I2(w2[13]),
        .I3(w0[13]),
        .O(p_2_in[13]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[14]_i_1 
       (.I0(prev_key1_new0_in[14]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[14]),
        .O(\prev_key1_reg[14]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[14]_i_2 
       (.I0(core_key[142]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[6]),
        .I3(Q[14]),
        .I4(\prev_key1_reg[14]_i_4_n_0 ),
        .O(prev_key1_new0_in[14]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[14]_i_3 
       (.I0(core_key[14]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[14]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[14]),
        .I5(new_sboxw[6]),
        .O(prev_key1_new[14]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[14]_i_4 
       (.I0(w5[14]),
        .I1(w4[14]),
        .I2(w6[14]),
        .O(\prev_key1_reg[14]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[14]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[14] ),
        .I1(w1[14]),
        .I2(w2[14]),
        .I3(w0[14]),
        .O(p_2_in[14]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[15]_i_1 
       (.I0(prev_key1_new0_in[15]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[15]),
        .O(\prev_key1_reg[15]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[15]_i_2 
       (.I0(core_key[143]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[7]),
        .I3(Q[15]),
        .I4(\prev_key1_reg[15]_i_4_n_0 ),
        .O(prev_key1_new0_in[15]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[15]_i_3 
       (.I0(core_key[15]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[15]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[15]),
        .I5(new_sboxw[7]),
        .O(prev_key1_new[15]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[15]_i_4 
       (.I0(w5[15]),
        .I1(w4[15]),
        .I2(w6[15]),
        .O(\prev_key1_reg[15]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[15]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[15] ),
        .I1(w1[15]),
        .I2(w2[15]),
        .I3(w0[15]),
        .O(p_2_in[15]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[16]_i_1 
       (.I0(prev_key1_new0_in[16]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[16]),
        .O(\prev_key1_reg[16]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[16]_i_2 
       (.I0(core_key[144]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[8]),
        .I3(Q[16]),
        .I4(\prev_key1_reg[16]_i_4_n_0 ),
        .O(prev_key1_new0_in[16]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[16]_i_3 
       (.I0(core_key[16]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[16]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[16]),
        .I5(new_sboxw[8]),
        .O(prev_key1_new[16]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[16]_i_4 
       (.I0(w5[16]),
        .I1(w4[16]),
        .I2(w6[16]),
        .O(\prev_key1_reg[16]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[16]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[16] ),
        .I1(w1[16]),
        .I2(w2[16]),
        .I3(w0[16]),
        .O(p_2_in[16]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[17]_i_1 
       (.I0(prev_key1_new0_in[17]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[17]),
        .O(\prev_key1_reg[17]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[17]_i_2 
       (.I0(core_key[145]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[9]),
        .I3(Q[17]),
        .I4(\prev_key1_reg[17]_i_4_n_0 ),
        .O(prev_key1_new0_in[17]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[17]_i_3 
       (.I0(core_key[17]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[17]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[17]),
        .I5(new_sboxw[9]),
        .O(prev_key1_new[17]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[17]_i_4 
       (.I0(w5[17]),
        .I1(w4[17]),
        .I2(w6[17]),
        .O(\prev_key1_reg[17]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[17]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[17] ),
        .I1(w1[17]),
        .I2(w2[17]),
        .I3(w0[17]),
        .O(p_2_in[17]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[18]_i_1 
       (.I0(prev_key1_new0_in[18]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[18]),
        .O(\prev_key1_reg[18]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[18]_i_2 
       (.I0(core_key[146]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[10]),
        .I3(Q[18]),
        .I4(\prev_key1_reg[18]_i_4_n_0 ),
        .O(prev_key1_new0_in[18]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[18]_i_3 
       (.I0(core_key[18]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[18]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[18]),
        .I5(new_sboxw[10]),
        .O(prev_key1_new[18]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[18]_i_4 
       (.I0(w5[18]),
        .I1(w4[18]),
        .I2(w6[18]),
        .O(\prev_key1_reg[18]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[18]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[18] ),
        .I1(w1[18]),
        .I2(w2[18]),
        .I3(w0[18]),
        .O(p_2_in[18]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[19]_i_1 
       (.I0(prev_key1_new0_in[19]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[19]),
        .O(\prev_key1_reg[19]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[19]_i_2 
       (.I0(core_key[147]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[11]),
        .I3(Q[19]),
        .I4(\prev_key1_reg[19]_i_4_n_0 ),
        .O(prev_key1_new0_in[19]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[19]_i_3 
       (.I0(core_key[19]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[19]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[19]),
        .I5(new_sboxw[11]),
        .O(prev_key1_new[19]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[19]_i_4 
       (.I0(w5[19]),
        .I1(w4[19]),
        .I2(w6[19]),
        .O(\prev_key1_reg[19]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[19]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[19] ),
        .I1(w1[19]),
        .I2(w2[19]),
        .I3(w0[19]),
        .O(p_2_in[19]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[1]_i_1 
       (.I0(prev_key1_new0_in[1]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[1]),
        .O(\prev_key1_reg[1]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[1]_i_2 
       (.I0(core_key[129]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[25]),
        .I3(Q[1]),
        .I4(\prev_key1_reg[1]_i_4_n_0 ),
        .O(prev_key1_new0_in[1]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[1]_i_3 
       (.I0(core_key[1]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[1]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[1]),
        .I5(new_sboxw[25]),
        .O(prev_key1_new[1]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[1]_i_4 
       (.I0(w5[1]),
        .I1(w4[1]),
        .I2(w6[1]),
        .O(\prev_key1_reg[1]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[1]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[1] ),
        .I1(w1[1]),
        .I2(w2[1]),
        .I3(w0[1]),
        .O(p_2_in[1]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[20]_i_1 
       (.I0(prev_key1_new0_in[20]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[20]),
        .O(\prev_key1_reg[20]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[20]_i_2 
       (.I0(core_key[148]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[12]),
        .I3(Q[20]),
        .I4(\prev_key1_reg[20]_i_4_n_0 ),
        .O(prev_key1_new0_in[20]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[20]_i_3 
       (.I0(core_key[20]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[20]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[20]),
        .I5(new_sboxw[12]),
        .O(prev_key1_new[20]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[20]_i_4 
       (.I0(w5[20]),
        .I1(w4[20]),
        .I2(w6[20]),
        .O(\prev_key1_reg[20]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[20]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[20] ),
        .I1(w1[20]),
        .I2(w2[20]),
        .I3(w0[20]),
        .O(p_2_in[20]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[21]_i_1 
       (.I0(prev_key1_new0_in[21]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[21]),
        .O(\prev_key1_reg[21]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[21]_i_2 
       (.I0(core_key[149]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[13]),
        .I3(Q[21]),
        .I4(\prev_key1_reg[21]_i_4_n_0 ),
        .O(prev_key1_new0_in[21]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[21]_i_3 
       (.I0(core_key[21]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[21]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[21]),
        .I5(new_sboxw[13]),
        .O(prev_key1_new[21]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[21]_i_4 
       (.I0(w5[21]),
        .I1(w4[21]),
        .I2(w6[21]),
        .O(\prev_key1_reg[21]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[21]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[21] ),
        .I1(w1[21]),
        .I2(w2[21]),
        .I3(w0[21]),
        .O(p_2_in[21]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[22]_i_1 
       (.I0(prev_key1_new0_in[22]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[22]),
        .O(\prev_key1_reg[22]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[22]_i_2 
       (.I0(core_key[150]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[14]),
        .I3(Q[22]),
        .I4(\prev_key1_reg[22]_i_4_n_0 ),
        .O(prev_key1_new0_in[22]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[22]_i_3 
       (.I0(core_key[22]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[22]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[22]),
        .I5(new_sboxw[14]),
        .O(prev_key1_new[22]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[22]_i_4 
       (.I0(w5[22]),
        .I1(w4[22]),
        .I2(w6[22]),
        .O(\prev_key1_reg[22]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[22]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[22] ),
        .I1(w1[22]),
        .I2(w2[22]),
        .I3(w0[22]),
        .O(p_2_in[22]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[23]_i_1 
       (.I0(prev_key1_new0_in[23]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[23]),
        .O(\prev_key1_reg[23]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[23]_i_2 
       (.I0(core_key[151]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[15]),
        .I3(Q[23]),
        .I4(\prev_key1_reg[23]_i_4_n_0 ),
        .O(prev_key1_new0_in[23]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[23]_i_3 
       (.I0(core_key[23]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[23]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[23]),
        .I5(new_sboxw[15]),
        .O(prev_key1_new[23]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[23]_i_4 
       (.I0(w5[23]),
        .I1(w4[23]),
        .I2(w6[23]),
        .O(\prev_key1_reg[23]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[23]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[23] ),
        .I1(w1[23]),
        .I2(w2[23]),
        .I3(w0[23]),
        .O(p_2_in[23]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[24]_i_1 
       (.I0(prev_key1_new0_in[24]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[24]),
        .O(\prev_key1_reg[24]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[24]_i_2 
       (.I0(core_key[152]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[16]),
        .I3(\rcon_reg_reg[7]_0 [0]),
        .I4(Q[24]),
        .I5(\prev_key1_reg[24]_i_4_n_0 ),
        .O(prev_key1_new0_in[24]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[24]_i_3 
       (.I0(core_key[24]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[24]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[24]),
        .I5(p_19_in[0]),
        .O(prev_key1_new[24]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[24]_i_4 
       (.I0(w5[24]),
        .I1(w4[24]),
        .I2(w6[24]),
        .O(\prev_key1_reg[24]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[24]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[24] ),
        .I1(w1[24]),
        .I2(w2[24]),
        .I3(w0[24]),
        .O(p_2_in[24]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[25]_i_1 
       (.I0(prev_key1_new0_in[25]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[25]),
        .O(\prev_key1_reg[25]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[25]_i_2 
       (.I0(core_key[153]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[17]),
        .I3(\rcon_reg_reg[7]_0 [1]),
        .I4(Q[25]),
        .I5(\prev_key1_reg[25]_i_4_n_0 ),
        .O(prev_key1_new0_in[25]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[25]_i_3 
       (.I0(core_key[25]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[25]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[25]),
        .I5(p_19_in[1]),
        .O(prev_key1_new[25]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[25]_i_4 
       (.I0(w5[25]),
        .I1(w4[25]),
        .I2(w6[25]),
        .O(\prev_key1_reg[25]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[25]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[25] ),
        .I1(w1[25]),
        .I2(w2[25]),
        .I3(w0[25]),
        .O(p_2_in[25]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[26]_i_1 
       (.I0(prev_key1_new0_in[26]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[26]),
        .O(\prev_key1_reg[26]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[26]_i_2 
       (.I0(core_key[154]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[18]),
        .I3(\rcon_reg_reg[7]_0 [2]),
        .I4(Q[26]),
        .I5(\prev_key1_reg[26]_i_4_n_0 ),
        .O(prev_key1_new0_in[26]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[26]_i_3 
       (.I0(core_key[26]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[26]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[26]),
        .I5(p_19_in[2]),
        .O(prev_key1_new[26]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[26]_i_4 
       (.I0(w5[26]),
        .I1(w4[26]),
        .I2(w6[26]),
        .O(\prev_key1_reg[26]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[26]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[26] ),
        .I1(w1[26]),
        .I2(w2[26]),
        .I3(w0[26]),
        .O(p_2_in[26]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[27]_i_1 
       (.I0(prev_key1_new0_in[27]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[27]),
        .O(\prev_key1_reg[27]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[27]_i_2 
       (.I0(core_key[155]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[19]),
        .I3(\rcon_reg_reg[7]_0 [3]),
        .I4(Q[27]),
        .I5(\prev_key1_reg[27]_i_4_n_0 ),
        .O(prev_key1_new0_in[27]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[27]_i_3 
       (.I0(core_key[27]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[27]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[27]),
        .I5(p_19_in[3]),
        .O(prev_key1_new[27]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[27]_i_4 
       (.I0(w5[27]),
        .I1(w4[27]),
        .I2(w6[27]),
        .O(\prev_key1_reg[27]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[27]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[27] ),
        .I1(w1[27]),
        .I2(w2[27]),
        .I3(w0[27]),
        .O(p_2_in[27]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[28]_i_1 
       (.I0(prev_key1_new0_in[28]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[28]),
        .O(\prev_key1_reg[28]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[28]_i_2 
       (.I0(core_key[156]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[20]),
        .I3(\rcon_reg_reg[7]_0 [4]),
        .I4(Q[28]),
        .I5(\prev_key1_reg[28]_i_4_n_0 ),
        .O(prev_key1_new0_in[28]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[28]_i_3 
       (.I0(core_key[28]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[28]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[28]),
        .I5(p_19_in[4]),
        .O(prev_key1_new[28]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[28]_i_4 
       (.I0(w5[28]),
        .I1(w4[28]),
        .I2(w6[28]),
        .O(\prev_key1_reg[28]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[28]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[28] ),
        .I1(w1[28]),
        .I2(w2[28]),
        .I3(w0[28]),
        .O(p_2_in[28]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[29]_i_1 
       (.I0(prev_key1_new0_in[29]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[29]),
        .O(\prev_key1_reg[29]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[29]_i_2 
       (.I0(core_key[157]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[21]),
        .I3(\rcon_reg_reg[7]_0 [5]),
        .I4(Q[29]),
        .I5(\prev_key1_reg[29]_i_4_n_0 ),
        .O(prev_key1_new0_in[29]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[29]_i_3 
       (.I0(core_key[29]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[29]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[29]),
        .I5(p_19_in[5]),
        .O(prev_key1_new[29]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[29]_i_4 
       (.I0(w5[29]),
        .I1(w4[29]),
        .I2(w6[29]),
        .O(\prev_key1_reg[29]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[29]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[29] ),
        .I1(w1[29]),
        .I2(w2[29]),
        .I3(w0[29]),
        .O(p_2_in[29]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[2]_i_1 
       (.I0(prev_key1_new0_in[2]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[2]),
        .O(\prev_key1_reg[2]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[2]_i_2 
       (.I0(core_key[130]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[26]),
        .I3(Q[2]),
        .I4(\prev_key1_reg[2]_i_4_n_0 ),
        .O(prev_key1_new0_in[2]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[2]_i_3 
       (.I0(core_key[2]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[2]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[2]),
        .I5(new_sboxw[26]),
        .O(prev_key1_new[2]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[2]_i_4 
       (.I0(w5[2]),
        .I1(w4[2]),
        .I2(w6[2]),
        .O(\prev_key1_reg[2]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[2]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[2] ),
        .I1(w1[2]),
        .I2(w2[2]),
        .I3(w0[2]),
        .O(p_2_in[2]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[30]_i_1 
       (.I0(prev_key1_new0_in[30]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[30]),
        .O(\prev_key1_reg[30]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[30]_i_2 
       (.I0(core_key[158]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[22]),
        .I3(\rcon_reg_reg[7]_0 [6]),
        .I4(Q[30]),
        .I5(\prev_key1_reg[30]_i_4_n_0 ),
        .O(prev_key1_new0_in[30]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[30]_i_3 
       (.I0(core_key[30]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[30]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[30]),
        .I5(p_19_in[6]),
        .O(prev_key1_new[30]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[30]_i_4 
       (.I0(w5[30]),
        .I1(w4[30]),
        .I2(w6[30]),
        .O(\prev_key1_reg[30]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[30]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[30] ),
        .I1(w1[30]),
        .I2(w2[30]),
        .I3(w0[30]),
        .O(p_2_in[30]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[31]_i_1 
       (.I0(prev_key1_new0_in[31]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[31]),
        .O(\prev_key1_reg[31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[31]_i_2 
       (.I0(core_key[159]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[23]),
        .I3(\rcon_reg_reg[7]_0 [7]),
        .I4(Q[31]),
        .I5(\prev_key1_reg[31]_i_4_n_0 ),
        .O(prev_key1_new0_in[31]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[31]_i_3 
       (.I0(core_key[31]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[31]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[31]),
        .I5(p_19_in[7]),
        .O(prev_key1_new[31]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[31]_i_4 
       (.I0(w5[31]),
        .I1(w4[31]),
        .I2(w6[31]),
        .O(\prev_key1_reg[31]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[31]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[31] ),
        .I1(w1[31]),
        .I2(w2[31]),
        .I3(w0[31]),
        .O(p_2_in[31]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[32]_i_1 
       (.I0(prev_key1_new0_in[32]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[32]),
        .O(\prev_key1_reg[32]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[32]_i_2 
       (.I0(core_key[160]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[24]),
        .I3(w6[0]),
        .I4(w4[0]),
        .I5(w5[0]),
        .O(prev_key1_new0_in[32]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[32]_i_3 
       (.I0(core_key[32]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[0]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[0]),
        .I5(new_sboxw[24]),
        .O(prev_key1_new[32]));
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[32]_i_4 
       (.I0(w0[0]),
        .I1(w2[0]),
        .I2(w1[0]),
        .O(p_6_in[0]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[33]_i_1 
       (.I0(prev_key1_new0_in[33]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[33]),
        .O(\prev_key1_reg[33]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[33]_i_2 
       (.I0(core_key[161]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[25]),
        .I3(w6[1]),
        .I4(w4[1]),
        .I5(w5[1]),
        .O(prev_key1_new0_in[33]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[33]_i_3 
       (.I0(core_key[33]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[1]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[1]),
        .I5(new_sboxw[25]),
        .O(prev_key1_new[33]));
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[33]_i_4 
       (.I0(w0[1]),
        .I1(w2[1]),
        .I2(w1[1]),
        .O(p_6_in[1]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[34]_i_1 
       (.I0(prev_key1_new0_in[34]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[34]),
        .O(\prev_key1_reg[34]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[34]_i_2 
       (.I0(core_key[162]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[26]),
        .I3(w6[2]),
        .I4(w4[2]),
        .I5(w5[2]),
        .O(prev_key1_new0_in[34]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[34]_i_3 
       (.I0(core_key[34]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[2]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[2]),
        .I5(new_sboxw[26]),
        .O(prev_key1_new[34]));
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[34]_i_4 
       (.I0(w0[2]),
        .I1(w2[2]),
        .I2(w1[2]),
        .O(p_6_in[2]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[35]_i_1 
       (.I0(prev_key1_new0_in[35]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[35]),
        .O(\prev_key1_reg[35]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[35]_i_2 
       (.I0(core_key[163]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[27]),
        .I3(w6[3]),
        .I4(w4[3]),
        .I5(w5[3]),
        .O(prev_key1_new0_in[35]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[35]_i_3 
       (.I0(core_key[35]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[3]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[3]),
        .I5(new_sboxw[27]),
        .O(prev_key1_new[35]));
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[35]_i_4 
       (.I0(w0[3]),
        .I1(w2[3]),
        .I2(w1[3]),
        .O(p_6_in[3]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[36]_i_1 
       (.I0(prev_key1_new0_in[36]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[36]),
        .O(\prev_key1_reg[36]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[36]_i_2 
       (.I0(core_key[164]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[28]),
        .I3(w6[4]),
        .I4(w4[4]),
        .I5(w5[4]),
        .O(prev_key1_new0_in[36]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[36]_i_3 
       (.I0(core_key[36]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[4]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[4]),
        .I5(new_sboxw[28]),
        .O(prev_key1_new[36]));
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[36]_i_4 
       (.I0(w0[4]),
        .I1(w2[4]),
        .I2(w1[4]),
        .O(p_6_in[4]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[37]_i_1 
       (.I0(prev_key1_new0_in[37]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[37]),
        .O(\prev_key1_reg[37]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[37]_i_2 
       (.I0(core_key[165]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[29]),
        .I3(w6[5]),
        .I4(w4[5]),
        .I5(w5[5]),
        .O(prev_key1_new0_in[37]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[37]_i_3 
       (.I0(core_key[37]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[5]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[5]),
        .I5(new_sboxw[29]),
        .O(prev_key1_new[37]));
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[37]_i_4 
       (.I0(w0[5]),
        .I1(w2[5]),
        .I2(w1[5]),
        .O(p_6_in[5]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[38]_i_1 
       (.I0(prev_key1_new0_in[38]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[38]),
        .O(\prev_key1_reg[38]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[38]_i_2 
       (.I0(core_key[166]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[30]),
        .I3(w6[6]),
        .I4(w4[6]),
        .I5(w5[6]),
        .O(prev_key1_new0_in[38]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[38]_i_3 
       (.I0(core_key[38]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[6]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[6]),
        .I5(new_sboxw[30]),
        .O(prev_key1_new[38]));
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[38]_i_4 
       (.I0(w0[6]),
        .I1(w2[6]),
        .I2(w1[6]),
        .O(p_6_in[6]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[39]_i_1 
       (.I0(prev_key1_new0_in[39]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[39]),
        .O(\prev_key1_reg[39]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[39]_i_2 
       (.I0(core_key[167]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[31]),
        .I3(w6[7]),
        .I4(w4[7]),
        .I5(w5[7]),
        .O(prev_key1_new0_in[39]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[39]_i_3 
       (.I0(core_key[39]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[7]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[7]),
        .I5(new_sboxw[31]),
        .O(prev_key1_new[39]));
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[39]_i_4 
       (.I0(w0[7]),
        .I1(w2[7]),
        .I2(w1[7]),
        .O(p_6_in[7]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[3]_i_1 
       (.I0(prev_key1_new0_in[3]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[3]),
        .O(\prev_key1_reg[3]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[3]_i_2 
       (.I0(core_key[131]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[27]),
        .I3(Q[3]),
        .I4(\prev_key1_reg[3]_i_4_n_0 ),
        .O(prev_key1_new0_in[3]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[3]_i_3 
       (.I0(core_key[3]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[3]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[3]),
        .I5(new_sboxw[27]),
        .O(prev_key1_new[3]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[3]_i_4 
       (.I0(w5[3]),
        .I1(w4[3]),
        .I2(w6[3]),
        .O(\prev_key1_reg[3]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[3]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[3] ),
        .I1(w1[3]),
        .I2(w2[3]),
        .I3(w0[3]),
        .O(p_2_in[3]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[40]_i_1 
       (.I0(prev_key1_new0_in[40]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[40]),
        .O(\prev_key1_reg[40]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[40]_i_2 
       (.I0(core_key[168]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[0]),
        .I3(w6[8]),
        .I4(w4[8]),
        .I5(w5[8]),
        .O(prev_key1_new0_in[40]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[40]_i_3 
       (.I0(core_key[40]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[8]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[8]),
        .I5(new_sboxw[0]),
        .O(prev_key1_new[40]));
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[40]_i_4 
       (.I0(w0[8]),
        .I1(w2[8]),
        .I2(w1[8]),
        .O(p_6_in[8]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[41]_i_1 
       (.I0(prev_key1_new0_in[41]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[41]),
        .O(\prev_key1_reg[41]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[41]_i_2 
       (.I0(core_key[169]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[1]),
        .I3(w6[9]),
        .I4(w4[9]),
        .I5(w5[9]),
        .O(prev_key1_new0_in[41]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[41]_i_3 
       (.I0(core_key[41]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[9]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[9]),
        .I5(new_sboxw[1]),
        .O(prev_key1_new[41]));
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[41]_i_4 
       (.I0(w0[9]),
        .I1(w2[9]),
        .I2(w1[9]),
        .O(p_6_in[9]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[42]_i_1 
       (.I0(prev_key1_new0_in[42]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[42]),
        .O(\prev_key1_reg[42]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[42]_i_2 
       (.I0(core_key[170]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[2]),
        .I3(w6[10]),
        .I4(w4[10]),
        .I5(w5[10]),
        .O(prev_key1_new0_in[42]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[42]_i_3 
       (.I0(core_key[42]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[10]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[10]),
        .I5(new_sboxw[2]),
        .O(prev_key1_new[42]));
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[42]_i_4 
       (.I0(w0[10]),
        .I1(w2[10]),
        .I2(w1[10]),
        .O(p_6_in[10]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[43]_i_1 
       (.I0(prev_key1_new0_in[43]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[43]),
        .O(\prev_key1_reg[43]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[43]_i_2 
       (.I0(core_key[171]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[3]),
        .I3(w6[11]),
        .I4(w4[11]),
        .I5(w5[11]),
        .O(prev_key1_new0_in[43]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[43]_i_3 
       (.I0(core_key[43]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[11]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[11]),
        .I5(new_sboxw[3]),
        .O(prev_key1_new[43]));
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[43]_i_4 
       (.I0(w0[11]),
        .I1(w2[11]),
        .I2(w1[11]),
        .O(p_6_in[11]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[44]_i_1 
       (.I0(prev_key1_new0_in[44]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[44]),
        .O(\prev_key1_reg[44]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[44]_i_2 
       (.I0(core_key[172]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[4]),
        .I3(w6[12]),
        .I4(w4[12]),
        .I5(w5[12]),
        .O(prev_key1_new0_in[44]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[44]_i_3 
       (.I0(core_key[44]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[12]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[12]),
        .I5(new_sboxw[4]),
        .O(prev_key1_new[44]));
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[44]_i_4 
       (.I0(w0[12]),
        .I1(w2[12]),
        .I2(w1[12]),
        .O(p_6_in[12]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[45]_i_1 
       (.I0(prev_key1_new0_in[45]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[45]),
        .O(\prev_key1_reg[45]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[45]_i_2 
       (.I0(core_key[173]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[5]),
        .I3(w6[13]),
        .I4(w4[13]),
        .I5(w5[13]),
        .O(prev_key1_new0_in[45]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[45]_i_3 
       (.I0(core_key[45]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[13]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[13]),
        .I5(new_sboxw[5]),
        .O(prev_key1_new[45]));
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[45]_i_4 
       (.I0(w0[13]),
        .I1(w2[13]),
        .I2(w1[13]),
        .O(p_6_in[13]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[46]_i_1 
       (.I0(prev_key1_new0_in[46]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[46]),
        .O(\prev_key1_reg[46]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[46]_i_2 
       (.I0(core_key[174]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[6]),
        .I3(w6[14]),
        .I4(w4[14]),
        .I5(w5[14]),
        .O(prev_key1_new0_in[46]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[46]_i_3 
       (.I0(core_key[46]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[14]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[14]),
        .I5(new_sboxw[6]),
        .O(prev_key1_new[46]));
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[46]_i_4 
       (.I0(w0[14]),
        .I1(w2[14]),
        .I2(w1[14]),
        .O(p_6_in[14]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[47]_i_1 
       (.I0(prev_key1_new0_in[47]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[47]),
        .O(\prev_key1_reg[47]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[47]_i_2 
       (.I0(core_key[175]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[7]),
        .I3(w6[15]),
        .I4(w4[15]),
        .I5(w5[15]),
        .O(prev_key1_new0_in[47]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[47]_i_3 
       (.I0(core_key[47]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[15]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[15]),
        .I5(new_sboxw[7]),
        .O(prev_key1_new[47]));
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[47]_i_4 
       (.I0(w0[15]),
        .I1(w2[15]),
        .I2(w1[15]),
        .O(p_6_in[15]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[48]_i_1 
       (.I0(prev_key1_new0_in[48]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[48]),
        .O(\prev_key1_reg[48]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[48]_i_2 
       (.I0(core_key[176]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[8]),
        .I3(w6[16]),
        .I4(w4[16]),
        .I5(w5[16]),
        .O(prev_key1_new0_in[48]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[48]_i_3 
       (.I0(core_key[48]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[16]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[16]),
        .I5(new_sboxw[8]),
        .O(prev_key1_new[48]));
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[48]_i_4 
       (.I0(w0[16]),
        .I1(w2[16]),
        .I2(w1[16]),
        .O(p_6_in[16]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[49]_i_1 
       (.I0(prev_key1_new0_in[49]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[49]),
        .O(\prev_key1_reg[49]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[49]_i_2 
       (.I0(core_key[177]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[9]),
        .I3(w6[17]),
        .I4(w4[17]),
        .I5(w5[17]),
        .O(prev_key1_new0_in[49]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[49]_i_3 
       (.I0(core_key[49]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[17]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[17]),
        .I5(new_sboxw[9]),
        .O(prev_key1_new[49]));
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[49]_i_4 
       (.I0(w0[17]),
        .I1(w2[17]),
        .I2(w1[17]),
        .O(p_6_in[17]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[4]_i_1 
       (.I0(prev_key1_new0_in[4]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[4]),
        .O(\prev_key1_reg[4]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[4]_i_2 
       (.I0(core_key[132]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[28]),
        .I3(Q[4]),
        .I4(\prev_key1_reg[4]_i_4_n_0 ),
        .O(prev_key1_new0_in[4]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[4]_i_3 
       (.I0(core_key[4]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[4]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[4]),
        .I5(new_sboxw[28]),
        .O(prev_key1_new[4]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[4]_i_4 
       (.I0(w5[4]),
        .I1(w4[4]),
        .I2(w6[4]),
        .O(\prev_key1_reg[4]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[4]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[4] ),
        .I1(w1[4]),
        .I2(w2[4]),
        .I3(w0[4]),
        .O(p_2_in[4]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[50]_i_1 
       (.I0(prev_key1_new0_in[50]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[50]),
        .O(\prev_key1_reg[50]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[50]_i_2 
       (.I0(core_key[178]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[10]),
        .I3(w6[18]),
        .I4(w4[18]),
        .I5(w5[18]),
        .O(prev_key1_new0_in[50]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[50]_i_3 
       (.I0(core_key[50]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[18]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[18]),
        .I5(new_sboxw[10]),
        .O(prev_key1_new[50]));
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[50]_i_4 
       (.I0(w0[18]),
        .I1(w2[18]),
        .I2(w1[18]),
        .O(p_6_in[18]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[51]_i_1 
       (.I0(prev_key1_new0_in[51]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[51]),
        .O(\prev_key1_reg[51]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[51]_i_2 
       (.I0(core_key[179]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[11]),
        .I3(w6[19]),
        .I4(w4[19]),
        .I5(w5[19]),
        .O(prev_key1_new0_in[51]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[51]_i_3 
       (.I0(core_key[51]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[19]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[19]),
        .I5(new_sboxw[11]),
        .O(prev_key1_new[51]));
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[51]_i_4 
       (.I0(w0[19]),
        .I1(w2[19]),
        .I2(w1[19]),
        .O(p_6_in[19]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[52]_i_1 
       (.I0(prev_key1_new0_in[52]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[52]),
        .O(\prev_key1_reg[52]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[52]_i_2 
       (.I0(core_key[180]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[12]),
        .I3(w6[20]),
        .I4(w4[20]),
        .I5(w5[20]),
        .O(prev_key1_new0_in[52]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[52]_i_3 
       (.I0(core_key[52]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[20]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[20]),
        .I5(new_sboxw[12]),
        .O(prev_key1_new[52]));
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[52]_i_4 
       (.I0(w0[20]),
        .I1(w2[20]),
        .I2(w1[20]),
        .O(p_6_in[20]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[53]_i_1 
       (.I0(prev_key1_new0_in[53]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[53]),
        .O(\prev_key1_reg[53]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[53]_i_2 
       (.I0(core_key[181]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[13]),
        .I3(w6[21]),
        .I4(w4[21]),
        .I5(w5[21]),
        .O(prev_key1_new0_in[53]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[53]_i_3 
       (.I0(core_key[53]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[21]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[21]),
        .I5(new_sboxw[13]),
        .O(prev_key1_new[53]));
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[53]_i_4 
       (.I0(w0[21]),
        .I1(w2[21]),
        .I2(w1[21]),
        .O(p_6_in[21]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[54]_i_1 
       (.I0(prev_key1_new0_in[54]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[54]),
        .O(\prev_key1_reg[54]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[54]_i_2 
       (.I0(core_key[182]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[14]),
        .I3(w6[22]),
        .I4(w4[22]),
        .I5(w5[22]),
        .O(prev_key1_new0_in[54]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[54]_i_3 
       (.I0(core_key[54]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[22]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[22]),
        .I5(new_sboxw[14]),
        .O(prev_key1_new[54]));
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[54]_i_4 
       (.I0(w0[22]),
        .I1(w2[22]),
        .I2(w1[22]),
        .O(p_6_in[22]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[55]_i_1 
       (.I0(prev_key1_new0_in[55]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[55]),
        .O(\prev_key1_reg[55]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[55]_i_2 
       (.I0(core_key[183]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[15]),
        .I3(w6[23]),
        .I4(w4[23]),
        .I5(w5[23]),
        .O(prev_key1_new0_in[55]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[55]_i_3 
       (.I0(core_key[55]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[23]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[23]),
        .I5(new_sboxw[15]),
        .O(prev_key1_new[55]));
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[55]_i_4 
       (.I0(w0[23]),
        .I1(w2[23]),
        .I2(w1[23]),
        .O(p_6_in[23]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[56]_i_1 
       (.I0(prev_key1_new0_in[56]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[56]),
        .O(\prev_key1_reg[56]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[56]_i_2 
       (.I0(core_key[184]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(p_19_in[0]),
        .I3(w6[24]),
        .I4(w4[24]),
        .I5(w5[24]),
        .O(prev_key1_new0_in[56]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[56]_i_3 
       (.I0(core_key[56]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[24]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[24]),
        .I5(p_19_in[0]),
        .O(prev_key1_new[56]));
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[56]_i_4 
       (.I0(w0[24]),
        .I1(w2[24]),
        .I2(w1[24]),
        .O(p_6_in[24]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[57]_i_1 
       (.I0(prev_key1_new0_in[57]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[57]),
        .O(\prev_key1_reg[57]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[57]_i_2 
       (.I0(core_key[185]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(p_19_in[1]),
        .I3(w6[25]),
        .I4(w4[25]),
        .I5(w5[25]),
        .O(prev_key1_new0_in[57]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[57]_i_3 
       (.I0(core_key[57]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[25]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[25]),
        .I5(p_19_in[1]),
        .O(prev_key1_new[57]));
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[57]_i_4 
       (.I0(w0[25]),
        .I1(w2[25]),
        .I2(w1[25]),
        .O(p_6_in[25]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[58]_i_1 
       (.I0(prev_key1_new0_in[58]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[58]),
        .O(\prev_key1_reg[58]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[58]_i_2 
       (.I0(core_key[186]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(p_19_in[2]),
        .I3(w6[26]),
        .I4(w4[26]),
        .I5(w5[26]),
        .O(prev_key1_new0_in[58]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[58]_i_3 
       (.I0(core_key[58]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[26]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[26]),
        .I5(p_19_in[2]),
        .O(prev_key1_new[58]));
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[58]_i_4 
       (.I0(w0[26]),
        .I1(w2[26]),
        .I2(w1[26]),
        .O(p_6_in[26]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[59]_i_1 
       (.I0(prev_key1_new0_in[59]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[59]),
        .O(\prev_key1_reg[59]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[59]_i_2 
       (.I0(core_key[187]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(p_19_in[3]),
        .I3(w6[27]),
        .I4(w4[27]),
        .I5(w5[27]),
        .O(prev_key1_new0_in[59]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[59]_i_3 
       (.I0(core_key[59]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[27]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[27]),
        .I5(p_19_in[3]),
        .O(prev_key1_new[59]));
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[59]_i_4 
       (.I0(w0[27]),
        .I1(w2[27]),
        .I2(w1[27]),
        .O(p_6_in[27]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[5]_i_1 
       (.I0(prev_key1_new0_in[5]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[5]),
        .O(\prev_key1_reg[5]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[5]_i_2 
       (.I0(core_key[133]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[29]),
        .I3(Q[5]),
        .I4(\prev_key1_reg[5]_i_4_n_0 ),
        .O(prev_key1_new0_in[5]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[5]_i_3 
       (.I0(core_key[5]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[5]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[5]),
        .I5(new_sboxw[29]),
        .O(prev_key1_new[5]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[5]_i_4 
       (.I0(w5[5]),
        .I1(w4[5]),
        .I2(w6[5]),
        .O(\prev_key1_reg[5]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[5]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[5] ),
        .I1(w1[5]),
        .I2(w2[5]),
        .I3(w0[5]),
        .O(p_2_in[5]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[60]_i_1 
       (.I0(prev_key1_new0_in[60]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[60]),
        .O(\prev_key1_reg[60]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[60]_i_2 
       (.I0(core_key[188]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(p_19_in[4]),
        .I3(w6[28]),
        .I4(w4[28]),
        .I5(w5[28]),
        .O(prev_key1_new0_in[60]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[60]_i_3 
       (.I0(core_key[60]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[28]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[28]),
        .I5(p_19_in[4]),
        .O(prev_key1_new[60]));
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[60]_i_4 
       (.I0(w0[28]),
        .I1(w2[28]),
        .I2(w1[28]),
        .O(p_6_in[28]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[61]_i_1 
       (.I0(prev_key1_new0_in[61]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[61]),
        .O(\prev_key1_reg[61]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[61]_i_2 
       (.I0(core_key[189]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(p_19_in[5]),
        .I3(w6[29]),
        .I4(w4[29]),
        .I5(w5[29]),
        .O(prev_key1_new0_in[61]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[61]_i_3 
       (.I0(core_key[61]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[29]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[29]),
        .I5(p_19_in[5]),
        .O(prev_key1_new[61]));
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[61]_i_4 
       (.I0(w0[29]),
        .I1(w2[29]),
        .I2(w1[29]),
        .O(p_6_in[29]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[62]_i_1 
       (.I0(prev_key1_new0_in[62]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[62]),
        .O(\prev_key1_reg[62]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[62]_i_2 
       (.I0(core_key[190]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(p_19_in[6]),
        .I3(w6[30]),
        .I4(w4[30]),
        .I5(w5[30]),
        .O(prev_key1_new0_in[62]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[62]_i_3 
       (.I0(core_key[62]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[30]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[30]),
        .I5(p_19_in[6]),
        .O(prev_key1_new[62]));
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[62]_i_4 
       (.I0(w0[30]),
        .I1(w2[30]),
        .I2(w1[30]),
        .O(p_6_in[30]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[63]_i_1 
       (.I0(prev_key1_new0_in[63]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[63]),
        .O(\prev_key1_reg[63]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[63]_i_2 
       (.I0(core_key[191]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(p_19_in[7]),
        .I3(w6[31]),
        .I4(w4[31]),
        .I5(w5[31]),
        .O(prev_key1_new0_in[63]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[63]_i_3 
       (.I0(core_key[63]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[31]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_6_in[31]),
        .I5(p_19_in[7]),
        .O(prev_key1_new[63]));
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[63]_i_4 
       (.I0(w0[31]),
        .I1(w2[31]),
        .I2(w1[31]),
        .O(p_6_in[31]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[64]_i_1 
       (.I0(prev_key1_new0_in[64]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[64]),
        .O(\prev_key1_reg[64]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[64]_i_2 
       (.I0(core_key[192]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[24]),
        .I3(w5[0]),
        .I4(w4[0]),
        .O(prev_key1_new0_in[64]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[64]_i_3 
       (.I0(core_key[64]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[0]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[0]),
        .I5(new_sboxw[24]),
        .O(prev_key1_new[64]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[64]_i_4 
       (.I0(w0[0]),
        .I1(w1[0]),
        .O(p_10_in[0]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[65]_i_1 
       (.I0(prev_key1_new0_in[65]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[65]),
        .O(\prev_key1_reg[65]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[65]_i_2 
       (.I0(core_key[193]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[25]),
        .I3(w5[1]),
        .I4(w4[1]),
        .O(prev_key1_new0_in[65]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[65]_i_3 
       (.I0(core_key[65]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[1]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[1]),
        .I5(new_sboxw[25]),
        .O(prev_key1_new[65]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[65]_i_4 
       (.I0(w0[1]),
        .I1(w1[1]),
        .O(p_10_in[1]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[66]_i_1 
       (.I0(prev_key1_new0_in[66]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[66]),
        .O(\prev_key1_reg[66]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[66]_i_2 
       (.I0(core_key[194]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[26]),
        .I3(w5[2]),
        .I4(w4[2]),
        .O(prev_key1_new0_in[66]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[66]_i_3 
       (.I0(core_key[66]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[2]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[2]),
        .I5(new_sboxw[26]),
        .O(prev_key1_new[66]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[66]_i_4 
       (.I0(w0[2]),
        .I1(w1[2]),
        .O(p_10_in[2]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[67]_i_1 
       (.I0(prev_key1_new0_in[67]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[67]),
        .O(\prev_key1_reg[67]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[67]_i_2 
       (.I0(core_key[195]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[27]),
        .I3(w5[3]),
        .I4(w4[3]),
        .O(prev_key1_new0_in[67]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[67]_i_3 
       (.I0(core_key[67]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[3]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[3]),
        .I5(new_sboxw[27]),
        .O(prev_key1_new[67]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[67]_i_4 
       (.I0(w0[3]),
        .I1(w1[3]),
        .O(p_10_in[3]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[68]_i_1 
       (.I0(prev_key1_new0_in[68]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[68]),
        .O(\prev_key1_reg[68]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[68]_i_2 
       (.I0(core_key[196]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[28]),
        .I3(w5[4]),
        .I4(w4[4]),
        .O(prev_key1_new0_in[68]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[68]_i_3 
       (.I0(core_key[68]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[4]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[4]),
        .I5(new_sboxw[28]),
        .O(prev_key1_new[68]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[68]_i_4 
       (.I0(w0[4]),
        .I1(w1[4]),
        .O(p_10_in[4]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[69]_i_1 
       (.I0(prev_key1_new0_in[69]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[69]),
        .O(\prev_key1_reg[69]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[69]_i_2 
       (.I0(core_key[197]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[29]),
        .I3(w5[5]),
        .I4(w4[5]),
        .O(prev_key1_new0_in[69]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[69]_i_3 
       (.I0(core_key[69]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[5]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[5]),
        .I5(new_sboxw[29]),
        .O(prev_key1_new[69]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[69]_i_4 
       (.I0(w0[5]),
        .I1(w1[5]),
        .O(p_10_in[5]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[6]_i_1 
       (.I0(prev_key1_new0_in[6]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[6]),
        .O(\prev_key1_reg[6]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[6]_i_2 
       (.I0(core_key[134]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[30]),
        .I3(Q[6]),
        .I4(\prev_key1_reg[6]_i_4_n_0 ),
        .O(prev_key1_new0_in[6]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[6]_i_3 
       (.I0(core_key[6]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[6]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[6]),
        .I5(new_sboxw[30]),
        .O(prev_key1_new[6]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[6]_i_4 
       (.I0(w5[6]),
        .I1(w4[6]),
        .I2(w6[6]),
        .O(\prev_key1_reg[6]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[6]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[6] ),
        .I1(w1[6]),
        .I2(w2[6]),
        .I3(w0[6]),
        .O(p_2_in[6]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[70]_i_1 
       (.I0(prev_key1_new0_in[70]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[70]),
        .O(\prev_key1_reg[70]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[70]_i_2 
       (.I0(core_key[198]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[30]),
        .I3(w5[6]),
        .I4(w4[6]),
        .O(prev_key1_new0_in[70]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[70]_i_3 
       (.I0(core_key[70]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[6]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[6]),
        .I5(new_sboxw[30]),
        .O(prev_key1_new[70]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[70]_i_4 
       (.I0(w0[6]),
        .I1(w1[6]),
        .O(p_10_in[6]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[71]_i_1 
       (.I0(prev_key1_new0_in[71]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[71]),
        .O(\prev_key1_reg[71]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[71]_i_2 
       (.I0(core_key[199]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[31]),
        .I3(w5[7]),
        .I4(w4[7]),
        .O(prev_key1_new0_in[71]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[71]_i_3 
       (.I0(core_key[71]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[7]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[7]),
        .I5(new_sboxw[31]),
        .O(prev_key1_new[71]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[71]_i_4 
       (.I0(w0[7]),
        .I1(w1[7]),
        .O(p_10_in[7]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[72]_i_1 
       (.I0(prev_key1_new0_in[72]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[72]),
        .O(\prev_key1_reg[72]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[72]_i_2 
       (.I0(core_key[200]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[0]),
        .I3(w5[8]),
        .I4(w4[8]),
        .O(prev_key1_new0_in[72]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[72]_i_3 
       (.I0(core_key[72]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[8]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[8]),
        .I5(new_sboxw[0]),
        .O(prev_key1_new[72]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[72]_i_4 
       (.I0(w0[8]),
        .I1(w1[8]),
        .O(p_10_in[8]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[73]_i_1 
       (.I0(prev_key1_new0_in[73]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[73]),
        .O(\prev_key1_reg[73]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[73]_i_2 
       (.I0(core_key[201]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[1]),
        .I3(w5[9]),
        .I4(w4[9]),
        .O(prev_key1_new0_in[73]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[73]_i_3 
       (.I0(core_key[73]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[9]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[9]),
        .I5(new_sboxw[1]),
        .O(prev_key1_new[73]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[73]_i_4 
       (.I0(w0[9]),
        .I1(w1[9]),
        .O(p_10_in[9]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[74]_i_1 
       (.I0(prev_key1_new0_in[74]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[74]),
        .O(\prev_key1_reg[74]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[74]_i_2 
       (.I0(core_key[202]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[2]),
        .I3(w5[10]),
        .I4(w4[10]),
        .O(prev_key1_new0_in[74]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[74]_i_3 
       (.I0(core_key[74]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[10]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[10]),
        .I5(new_sboxw[2]),
        .O(prev_key1_new[74]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[74]_i_4 
       (.I0(w0[10]),
        .I1(w1[10]),
        .O(p_10_in[10]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[75]_i_1 
       (.I0(prev_key1_new0_in[75]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[75]),
        .O(\prev_key1_reg[75]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[75]_i_2 
       (.I0(core_key[203]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[3]),
        .I3(w5[11]),
        .I4(w4[11]),
        .O(prev_key1_new0_in[75]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[75]_i_3 
       (.I0(core_key[75]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[11]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[11]),
        .I5(new_sboxw[3]),
        .O(prev_key1_new[75]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[75]_i_4 
       (.I0(w0[11]),
        .I1(w1[11]),
        .O(p_10_in[11]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[76]_i_1 
       (.I0(prev_key1_new0_in[76]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[76]),
        .O(\prev_key1_reg[76]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[76]_i_2 
       (.I0(core_key[204]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[4]),
        .I3(w5[12]),
        .I4(w4[12]),
        .O(prev_key1_new0_in[76]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[76]_i_3 
       (.I0(core_key[76]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[12]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[12]),
        .I5(new_sboxw[4]),
        .O(prev_key1_new[76]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[76]_i_4 
       (.I0(w0[12]),
        .I1(w1[12]),
        .O(p_10_in[12]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[77]_i_1 
       (.I0(prev_key1_new0_in[77]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[77]),
        .O(\prev_key1_reg[77]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[77]_i_2 
       (.I0(core_key[205]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[5]),
        .I3(w5[13]),
        .I4(w4[13]),
        .O(prev_key1_new0_in[77]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[77]_i_3 
       (.I0(core_key[77]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[13]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[13]),
        .I5(new_sboxw[5]),
        .O(prev_key1_new[77]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[77]_i_4 
       (.I0(w0[13]),
        .I1(w1[13]),
        .O(p_10_in[13]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[78]_i_1 
       (.I0(prev_key1_new0_in[78]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[78]),
        .O(\prev_key1_reg[78]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[78]_i_2 
       (.I0(core_key[206]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[6]),
        .I3(w5[14]),
        .I4(w4[14]),
        .O(prev_key1_new0_in[78]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[78]_i_3 
       (.I0(core_key[78]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[14]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[14]),
        .I5(new_sboxw[6]),
        .O(prev_key1_new[78]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[78]_i_4 
       (.I0(w0[14]),
        .I1(w1[14]),
        .O(p_10_in[14]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[79]_i_1 
       (.I0(prev_key1_new0_in[79]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[79]),
        .O(\prev_key1_reg[79]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[79]_i_2 
       (.I0(core_key[207]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[7]),
        .I3(w5[15]),
        .I4(w4[15]),
        .O(prev_key1_new0_in[79]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[79]_i_3 
       (.I0(core_key[79]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[15]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[15]),
        .I5(new_sboxw[7]),
        .O(prev_key1_new[79]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[79]_i_4 
       (.I0(w0[15]),
        .I1(w1[15]),
        .O(p_10_in[15]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[7]_i_1 
       (.I0(prev_key1_new0_in[7]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[7]),
        .O(\prev_key1_reg[7]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[7]_i_2 
       (.I0(core_key[135]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[31]),
        .I3(Q[7]),
        .I4(\prev_key1_reg[7]_i_4_n_0 ),
        .O(prev_key1_new0_in[7]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[7]_i_3 
       (.I0(core_key[7]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[7]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[7]),
        .I5(new_sboxw[31]),
        .O(prev_key1_new[7]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[7]_i_4 
       (.I0(w5[7]),
        .I1(w4[7]),
        .I2(w6[7]),
        .O(\prev_key1_reg[7]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[7]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[7] ),
        .I1(w1[7]),
        .I2(w2[7]),
        .I3(w0[7]),
        .O(p_2_in[7]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[80]_i_1 
       (.I0(prev_key1_new0_in[80]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[80]),
        .O(\prev_key1_reg[80]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[80]_i_2 
       (.I0(core_key[208]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[8]),
        .I3(w5[16]),
        .I4(w4[16]),
        .O(prev_key1_new0_in[80]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[80]_i_3 
       (.I0(core_key[80]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[16]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[16]),
        .I5(new_sboxw[8]),
        .O(prev_key1_new[80]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[80]_i_4 
       (.I0(w0[16]),
        .I1(w1[16]),
        .O(p_10_in[16]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[81]_i_1 
       (.I0(prev_key1_new0_in[81]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[81]),
        .O(\prev_key1_reg[81]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[81]_i_2 
       (.I0(core_key[209]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[9]),
        .I3(w5[17]),
        .I4(w4[17]),
        .O(prev_key1_new0_in[81]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[81]_i_3 
       (.I0(core_key[81]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[17]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[17]),
        .I5(new_sboxw[9]),
        .O(prev_key1_new[81]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[81]_i_4 
       (.I0(w0[17]),
        .I1(w1[17]),
        .O(p_10_in[17]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[82]_i_1 
       (.I0(prev_key1_new0_in[82]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[82]),
        .O(\prev_key1_reg[82]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[82]_i_2 
       (.I0(core_key[210]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[10]),
        .I3(w5[18]),
        .I4(w4[18]),
        .O(prev_key1_new0_in[82]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[82]_i_3 
       (.I0(core_key[82]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[18]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[18]),
        .I5(new_sboxw[10]),
        .O(prev_key1_new[82]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[82]_i_4 
       (.I0(w0[18]),
        .I1(w1[18]),
        .O(p_10_in[18]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[83]_i_1 
       (.I0(prev_key1_new0_in[83]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[83]),
        .O(\prev_key1_reg[83]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[83]_i_2 
       (.I0(core_key[211]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[11]),
        .I3(w5[19]),
        .I4(w4[19]),
        .O(prev_key1_new0_in[83]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[83]_i_3 
       (.I0(core_key[83]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[19]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[19]),
        .I5(new_sboxw[11]),
        .O(prev_key1_new[83]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[83]_i_4 
       (.I0(w0[19]),
        .I1(w1[19]),
        .O(p_10_in[19]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[84]_i_1 
       (.I0(prev_key1_new0_in[84]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[84]),
        .O(\prev_key1_reg[84]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[84]_i_2 
       (.I0(core_key[212]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[12]),
        .I3(w5[20]),
        .I4(w4[20]),
        .O(prev_key1_new0_in[84]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[84]_i_3 
       (.I0(core_key[84]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[20]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[20]),
        .I5(new_sboxw[12]),
        .O(prev_key1_new[84]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[84]_i_4 
       (.I0(w0[20]),
        .I1(w1[20]),
        .O(p_10_in[20]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[85]_i_1 
       (.I0(prev_key1_new0_in[85]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[85]),
        .O(\prev_key1_reg[85]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[85]_i_2 
       (.I0(core_key[213]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[13]),
        .I3(w5[21]),
        .I4(w4[21]),
        .O(prev_key1_new0_in[85]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[85]_i_3 
       (.I0(core_key[85]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[21]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[21]),
        .I5(new_sboxw[13]),
        .O(prev_key1_new[85]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[85]_i_4 
       (.I0(w0[21]),
        .I1(w1[21]),
        .O(p_10_in[21]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[86]_i_1 
       (.I0(prev_key1_new0_in[86]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[86]),
        .O(\prev_key1_reg[86]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[86]_i_2 
       (.I0(core_key[214]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[14]),
        .I3(w5[22]),
        .I4(w4[22]),
        .O(prev_key1_new0_in[86]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[86]_i_3 
       (.I0(core_key[86]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[22]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[22]),
        .I5(new_sboxw[14]),
        .O(prev_key1_new[86]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[86]_i_4 
       (.I0(w0[22]),
        .I1(w1[22]),
        .O(p_10_in[22]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[87]_i_1 
       (.I0(prev_key1_new0_in[87]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[87]),
        .O(\prev_key1_reg[87]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[87]_i_2 
       (.I0(core_key[215]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[15]),
        .I3(w5[23]),
        .I4(w4[23]),
        .O(prev_key1_new0_in[87]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[87]_i_3 
       (.I0(core_key[87]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[23]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[23]),
        .I5(new_sboxw[15]),
        .O(prev_key1_new[87]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[87]_i_4 
       (.I0(w0[23]),
        .I1(w1[23]),
        .O(p_10_in[23]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[88]_i_1 
       (.I0(prev_key1_new0_in[88]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[88]),
        .O(\prev_key1_reg[88]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[88]_i_2 
       (.I0(core_key[216]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [0]),
        .I3(new_sboxw[16]),
        .I4(w5[24]),
        .I5(w4[24]),
        .O(prev_key1_new0_in[88]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[88]_i_3 
       (.I0(core_key[88]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[24]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_10_in[24]),
        .I5(p_19_in[0]),
        .O(prev_key1_new[88]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[88]_i_4 
       (.I0(w0[24]),
        .I1(w1[24]),
        .O(p_10_in[24]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[89]_i_1 
       (.I0(prev_key1_new0_in[89]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[89]),
        .O(\prev_key1_reg[89]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[89]_i_2 
       (.I0(core_key[217]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [1]),
        .I3(new_sboxw[17]),
        .I4(w5[25]),
        .I5(w4[25]),
        .O(prev_key1_new0_in[89]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[89]_i_3 
       (.I0(core_key[89]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[25]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(p_10_in[25]),
        .I5(p_19_in[1]),
        .O(prev_key1_new[89]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[89]_i_4 
       (.I0(w0[25]),
        .I1(w1[25]),
        .O(p_10_in[25]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[8]_i_1 
       (.I0(prev_key1_new0_in[8]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[8]),
        .O(\prev_key1_reg[8]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[8]_i_2 
       (.I0(core_key[136]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[0]),
        .I3(Q[8]),
        .I4(\prev_key1_reg[8]_i_4_n_0 ),
        .O(prev_key1_new0_in[8]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[8]_i_3 
       (.I0(core_key[8]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[8]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[8]),
        .I5(new_sboxw[0]),
        .O(prev_key1_new[8]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[8]_i_4 
       (.I0(w5[8]),
        .I1(w4[8]),
        .I2(w6[8]),
        .O(\prev_key1_reg[8]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[8]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[8] ),
        .I1(w1[8]),
        .I2(w2[8]),
        .I3(w0[8]),
        .O(p_2_in[8]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[90]_i_1 
       (.I0(prev_key1_new0_in[90]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[90]),
        .O(\prev_key1_reg[90]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[90]_i_2 
       (.I0(core_key[218]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [2]),
        .I3(new_sboxw[18]),
        .I4(w5[26]),
        .I5(w4[26]),
        .O(prev_key1_new0_in[90]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[90]_i_3 
       (.I0(core_key[90]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[26]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(p_10_in[26]),
        .I5(p_19_in[2]),
        .O(prev_key1_new[90]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[90]_i_4 
       (.I0(w0[26]),
        .I1(w1[26]),
        .O(p_10_in[26]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[91]_i_1 
       (.I0(prev_key1_new0_in[91]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[91]),
        .O(\prev_key1_reg[91]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[91]_i_2 
       (.I0(core_key[219]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [3]),
        .I3(new_sboxw[19]),
        .I4(w5[27]),
        .I5(w4[27]),
        .O(prev_key1_new0_in[91]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[91]_i_3 
       (.I0(core_key[91]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[27]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(p_10_in[27]),
        .I5(p_19_in[3]),
        .O(prev_key1_new[91]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[91]_i_4 
       (.I0(w0[27]),
        .I1(w1[27]),
        .O(p_10_in[27]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[92]_i_1 
       (.I0(prev_key1_new0_in[92]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[92]),
        .O(\prev_key1_reg[92]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[92]_i_2 
       (.I0(core_key[220]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [4]),
        .I3(new_sboxw[20]),
        .I4(w5[28]),
        .I5(w4[28]),
        .O(prev_key1_new0_in[92]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[92]_i_3 
       (.I0(core_key[92]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[28]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(p_10_in[28]),
        .I5(p_19_in[4]),
        .O(prev_key1_new[92]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[92]_i_4 
       (.I0(w0[28]),
        .I1(w1[28]),
        .O(p_10_in[28]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[93]_i_1 
       (.I0(prev_key1_new0_in[93]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[93]),
        .O(\prev_key1_reg[93]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[93]_i_2 
       (.I0(core_key[221]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [5]),
        .I3(new_sboxw[21]),
        .I4(w5[29]),
        .I5(w4[29]),
        .O(prev_key1_new0_in[93]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[93]_i_3 
       (.I0(core_key[93]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[29]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(p_10_in[29]),
        .I5(p_19_in[5]),
        .O(prev_key1_new[93]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[93]_i_4 
       (.I0(w0[29]),
        .I1(w1[29]),
        .O(p_10_in[29]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[94]_i_1 
       (.I0(prev_key1_new0_in[94]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[94]),
        .O(\prev_key1_reg[94]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[94]_i_2 
       (.I0(core_key[222]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [6]),
        .I3(new_sboxw[22]),
        .I4(w5[30]),
        .I5(w4[30]),
        .O(prev_key1_new0_in[94]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[94]_i_3 
       (.I0(core_key[94]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[30]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(p_10_in[30]),
        .I5(p_19_in[6]),
        .O(prev_key1_new[94]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[94]_i_4 
       (.I0(w0[30]),
        .I1(w1[30]),
        .O(p_10_in[30]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[95]_i_1 
       (.I0(prev_key1_new0_in[95]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[95]),
        .O(\prev_key1_reg[95]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \prev_key1_reg[95]_i_2 
       (.I0(core_key[223]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(\rcon_reg_reg[7]_0 [7]),
        .I3(new_sboxw[23]),
        .I4(w5[31]),
        .I5(w4[31]),
        .O(prev_key1_new0_in[95]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[95]_i_3 
       (.I0(core_key[95]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[31]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(p_10_in[31]),
        .I5(p_19_in[7]),
        .O(prev_key1_new[95]));
  LUT2 #(
    .INIT(4'h6)) 
    \prev_key1_reg[95]_i_4 
       (.I0(w0[31]),
        .I1(w1[31]),
        .O(p_10_in[31]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[96]_i_1 
       (.I0(prev_key1_new0_in[96]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[96]),
        .O(\prev_key1_reg[96]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[96]_i_2 
       (.I0(core_key[224]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[24]),
        .I3(w4[0]),
        .O(prev_key1_new0_in[96]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[96]_i_3 
       (.I0(core_key[96]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[0]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[0]),
        .I5(new_sboxw[24]),
        .O(prev_key1_new[96]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[97]_i_1 
       (.I0(prev_key1_new0_in[97]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[97]),
        .O(\prev_key1_reg[97]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[97]_i_2 
       (.I0(core_key[225]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[25]),
        .I3(w4[1]),
        .O(prev_key1_new0_in[97]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[97]_i_3 
       (.I0(core_key[97]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[1]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[1]),
        .I5(new_sboxw[25]),
        .O(prev_key1_new[97]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[98]_i_1 
       (.I0(prev_key1_new0_in[98]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[98]),
        .O(\prev_key1_reg[98]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[98]_i_2 
       (.I0(core_key[226]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[26]),
        .I3(w4[2]),
        .O(prev_key1_new0_in[98]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[98]_i_3 
       (.I0(core_key[98]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[2]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[2]),
        .I5(new_sboxw[26]),
        .O(prev_key1_new[98]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[99]_i_1 
       (.I0(prev_key1_new0_in[99]),
        .I1(\key_mem_reg[14][36]_0 ),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[99]),
        .O(\prev_key1_reg[99]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8BB8)) 
    \prev_key1_reg[99]_i_2 
       (.I0(core_key[227]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[27]),
        .I3(w4[3]),
        .O(prev_key1_new0_in[99]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[99]_i_3 
       (.I0(core_key[99]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[3]),
        .I3(\round_ctr_reg_reg[0]_rep__0_n_0 ),
        .I4(w0[3]),
        .I5(new_sboxw[27]),
        .O(prev_key1_new[99]));
  LUT4 #(
    .INIT(16'hE222)) 
    \prev_key1_reg[9]_i_1 
       (.I0(prev_key1_new0_in[9]),
        .I1(p_1_in[2]),
        .I2(\prev_key1_reg[127]_i_4_n_0 ),
        .I3(prev_key1_new[9]),
        .O(\prev_key1_reg[9]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB88B8BB8)) 
    \prev_key1_reg[9]_i_2 
       (.I0(core_key[137]),
        .I1(\key_mem[0][127]_i_3_n_0 ),
        .I2(new_sboxw[1]),
        .I3(Q[9]),
        .I4(\prev_key1_reg[9]_i_4_n_0 ),
        .O(prev_key1_new0_in[9]));
  LUT6 #(
    .INIT(64'h8B88B8BB8BBBB888)) 
    \prev_key1_reg[9]_i_3 
       (.I0(core_key[9]),
        .I1(\prev_key0_reg[127]_i_3_n_0 ),
        .I2(new_sboxw[9]),
        .I3(\round_ctr_reg_reg[0]_rep__1_n_0 ),
        .I4(p_2_in[9]),
        .I5(new_sboxw[1]),
        .O(prev_key1_new[9]));
  LUT3 #(
    .INIT(8'h96)) 
    \prev_key1_reg[9]_i_4 
       (.I0(w5[9]),
        .I1(w4[9]),
        .I2(w6[9]),
        .O(\prev_key1_reg[9]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \prev_key1_reg[9]_i_5 
       (.I0(\prev_key0_reg_reg_n_0_[9] ),
        .I1(w1[9]),
        .I2(w2[9]),
        .I3(w0[9]),
        .O(p_2_in[9]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[0] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[0]_i_1_n_0 ),
        .Q(Q[0]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[100] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[100]_i_1_n_0 ),
        .Q(w4[4]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[101] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[101]_i_1_n_0 ),
        .Q(w4[5]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[102] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[102]_i_1_n_0 ),
        .Q(w4[6]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[103] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[103]_i_1_n_0 ),
        .Q(w4[7]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[104] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[104]_i_1_n_0 ),
        .Q(w4[8]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[105] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[105]_i_1_n_0 ),
        .Q(w4[9]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[106] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[106]_i_1_n_0 ),
        .Q(w4[10]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[107] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[107]_i_1_n_0 ),
        .Q(w4[11]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[108] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[108]_i_1_n_0 ),
        .Q(w4[12]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[109] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[109]_i_1_n_0 ),
        .Q(w4[13]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[10] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[10]_i_1_n_0 ),
        .Q(Q[10]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[110] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[110]_i_1_n_0 ),
        .Q(w4[14]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[111] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[111]_i_1_n_0 ),
        .Q(w4[15]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[112] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[112]_i_1_n_0 ),
        .Q(w4[16]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[113] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[113]_i_1_n_0 ),
        .Q(w4[17]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[114] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[114]_i_1_n_0 ),
        .Q(w4[18]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[115] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[115]_i_1_n_0 ),
        .Q(w4[19]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[116] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[116]_i_1_n_0 ),
        .Q(w4[20]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[117] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[117]_i_1_n_0 ),
        .Q(w4[21]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[118] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[118]_i_1_n_0 ),
        .Q(w4[22]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[119] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[119]_i_1_n_0 ),
        .Q(w4[23]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[11] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[11]_i_1_n_0 ),
        .Q(Q[11]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[120] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[120]_i_1_n_0 ),
        .Q(w4[24]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[121] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[121]_i_1_n_0 ),
        .Q(w4[25]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[122] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[122]_i_1_n_0 ),
        .Q(w4[26]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[123] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[123]_i_1_n_0 ),
        .Q(w4[27]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[124] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[124]_i_1_n_0 ),
        .Q(w4[28]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[125] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[125]_i_1_n_0 ),
        .Q(w4[29]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[126] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[126]_i_1_n_0 ),
        .Q(w4[30]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[127] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[127]_i_2_n_0 ),
        .Q(w4[31]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[12] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[12]_i_1_n_0 ),
        .Q(Q[12]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[13] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[13]_i_1_n_0 ),
        .Q(Q[13]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[14] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[14]_i_1_n_0 ),
        .Q(Q[14]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[15] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[15]_i_1_n_0 ),
        .Q(Q[15]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[16] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[16]_i_1_n_0 ),
        .Q(Q[16]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[17] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[17]_i_1_n_0 ),
        .Q(Q[17]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[18] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[18]_i_1_n_0 ),
        .Q(Q[18]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[19] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[19]_i_1_n_0 ),
        .Q(Q[19]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[1] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[1]_i_1_n_0 ),
        .Q(Q[1]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[20] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[20]_i_1_n_0 ),
        .Q(Q[20]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[21] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[21]_i_1_n_0 ),
        .Q(Q[21]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[22] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[22]_i_1_n_0 ),
        .Q(Q[22]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[23] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[23]_i_1_n_0 ),
        .Q(Q[23]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[24] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[24]_i_1_n_0 ),
        .Q(Q[24]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[25] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[25]_i_1_n_0 ),
        .Q(Q[25]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[26] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[26]_i_1_n_0 ),
        .Q(Q[26]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[27] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[27]_i_1_n_0 ),
        .Q(Q[27]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[28] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[28]_i_1_n_0 ),
        .Q(Q[28]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[29] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[29]_i_1_n_0 ),
        .Q(Q[29]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[2] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[2]_i_1_n_0 ),
        .Q(Q[2]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[30] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[30]_i_1_n_0 ),
        .Q(Q[30]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[31] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[31]_i_1_n_0 ),
        .Q(Q[31]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[32] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[32]_i_1_n_0 ),
        .Q(w6[0]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[33] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[33]_i_1_n_0 ),
        .Q(w6[1]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[34] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[34]_i_1_n_0 ),
        .Q(w6[2]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[35] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[35]_i_1_n_0 ),
        .Q(w6[3]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[36] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[36]_i_1_n_0 ),
        .Q(w6[4]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[37] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[37]_i_1_n_0 ),
        .Q(w6[5]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[38] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[38]_i_1_n_0 ),
        .Q(w6[6]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[39] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[39]_i_1_n_0 ),
        .Q(w6[7]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[3] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[3]_i_1_n_0 ),
        .Q(Q[3]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[40] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[40]_i_1_n_0 ),
        .Q(w6[8]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[41] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[41]_i_1_n_0 ),
        .Q(w6[9]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[42] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[42]_i_1_n_0 ),
        .Q(w6[10]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[43] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[43]_i_1_n_0 ),
        .Q(w6[11]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[44] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[44]_i_1_n_0 ),
        .Q(w6[12]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[45] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[45]_i_1_n_0 ),
        .Q(w6[13]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[46] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[46]_i_1_n_0 ),
        .Q(w6[14]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[47] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[47]_i_1_n_0 ),
        .Q(w6[15]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[48] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[48]_i_1_n_0 ),
        .Q(w6[16]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[49] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[49]_i_1_n_0 ),
        .Q(w6[17]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[4] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[4]_i_1_n_0 ),
        .Q(Q[4]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[50] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[50]_i_1_n_0 ),
        .Q(w6[18]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[51] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[51]_i_1_n_0 ),
        .Q(w6[19]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[52] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[52]_i_1_n_0 ),
        .Q(w6[20]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[53] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[53]_i_1_n_0 ),
        .Q(w6[21]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[54] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[54]_i_1_n_0 ),
        .Q(w6[22]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[55] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[55]_i_1_n_0 ),
        .Q(w6[23]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[56] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[56]_i_1_n_0 ),
        .Q(w6[24]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[57] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[57]_i_1_n_0 ),
        .Q(w6[25]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[58] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[58]_i_1_n_0 ),
        .Q(w6[26]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[59] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[59]_i_1_n_0 ),
        .Q(w6[27]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[5] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[5]_i_1_n_0 ),
        .Q(Q[5]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[60] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[60]_i_1_n_0 ),
        .Q(w6[28]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[61] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[61]_i_1_n_0 ),
        .Q(w6[29]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[62] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[62]_i_1_n_0 ),
        .Q(w6[30]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[63] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[63]_i_1_n_0 ),
        .Q(w6[31]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[64] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[64]_i_1_n_0 ),
        .Q(w5[0]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[65] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[65]_i_1_n_0 ),
        .Q(w5[1]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[66] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[66]_i_1_n_0 ),
        .Q(w5[2]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[67] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[67]_i_1_n_0 ),
        .Q(w5[3]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[68] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[68]_i_1_n_0 ),
        .Q(w5[4]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[69] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[69]_i_1_n_0 ),
        .Q(w5[5]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[6] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[6]_i_1_n_0 ),
        .Q(Q[6]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[70] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[70]_i_1_n_0 ),
        .Q(w5[6]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[71] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[71]_i_1_n_0 ),
        .Q(w5[7]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[72] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[72]_i_1_n_0 ),
        .Q(w5[8]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[73] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[73]_i_1_n_0 ),
        .Q(w5[9]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[74] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[74]_i_1_n_0 ),
        .Q(w5[10]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[75] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[75]_i_1_n_0 ),
        .Q(w5[11]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[76] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[76]_i_1_n_0 ),
        .Q(w5[12]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[77] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[77]_i_1_n_0 ),
        .Q(w5[13]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[78] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[78]_i_1_n_0 ),
        .Q(w5[14]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[79] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[79]_i_1_n_0 ),
        .Q(w5[15]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[7] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[7]_i_1_n_0 ),
        .Q(Q[7]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[80] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[80]_i_1_n_0 ),
        .Q(w5[16]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[81] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[81]_i_1_n_0 ),
        .Q(w5[17]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[82] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[82]_i_1_n_0 ),
        .Q(w5[18]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[83] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[83]_i_1_n_0 ),
        .Q(w5[19]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[84] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[84]_i_1_n_0 ),
        .Q(w5[20]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[85] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[85]_i_1_n_0 ),
        .Q(w5[21]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[86] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[86]_i_1_n_0 ),
        .Q(w5[22]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[87] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[87]_i_1_n_0 ),
        .Q(w5[23]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[88] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[88]_i_1_n_0 ),
        .Q(w5[24]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[89] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[89]_i_1_n_0 ),
        .Q(w5[25]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[8] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[8]_i_1_n_0 ),
        .Q(Q[8]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[90] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[90]_i_1_n_0 ),
        .Q(w5[26]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[91] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[91]_i_1_n_0 ),
        .Q(w5[27]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[92] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[92]_i_1_n_0 ),
        .Q(w5[28]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[93] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[93]_i_1_n_0 ),
        .Q(w5[29]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[94] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[94]_i_1_n_0 ),
        .Q(w5[30]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[95] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[95]_i_1_n_0 ),
        .Q(w5[31]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[96] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[96]_i_1_n_0 ),
        .Q(w4[0]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[97] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[97]_i_1_n_0 ),
        .Q(w4[1]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[98] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[98]_i_1_n_0 ),
        .Q(w4[2]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[99] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[99]_i_1_n_0 ),
        .Q(w4[3]));
  FDCE #(
    .INIT(1'b0)) 
    \prev_key1_reg_reg[9] 
       (.C(clk_i),
        .CE(prev_key1_we1_out),
        .CLR(rst_i),
        .D(\prev_key1_reg[9]_i_1_n_0 ),
        .Q(Q[9]));
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT4 #(
    .INIT(16'hB3BB)) 
    \rcon_reg[0]_i_1 
       (.I0(\rcon_reg_reg[7]_0 [7]),
        .I1(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I2(\round_ctr_reg_reg[0]_rep_n_0 ),
        .I3(p_1_in[2]),
        .O(rcon_new[0]));
  LUT5 #(
    .INIT(32'h00D0D000)) 
    \rcon_reg[1]_i_1 
       (.I0(p_1_in[2]),
        .I1(\round_ctr_reg_reg[0]_rep_n_0 ),
        .I2(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I3(\rcon_reg_reg[7]_0 [0]),
        .I4(\rcon_reg_reg[7]_0 [7]),
        .O(rcon_new[1]));
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT4 #(
    .INIT(16'hB3BB)) 
    \rcon_reg[2]_i_1 
       (.I0(\rcon_reg_reg[7]_0 [1]),
        .I1(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I2(\round_ctr_reg_reg[0]_rep_n_0 ),
        .I3(p_1_in[2]),
        .O(rcon_new[2]));
  LUT5 #(
    .INIT(32'h6F0F6F6F)) 
    \rcon_reg[3]_i_1 
       (.I0(\rcon_reg_reg[7]_0 [7]),
        .I1(\rcon_reg_reg[7]_0 [2]),
        .I2(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I3(\round_ctr_reg_reg[0]_rep_n_0 ),
        .I4(p_1_in[2]),
        .O(rcon_new[3]));
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT5 #(
    .INIT(32'h00D0D000)) 
    \rcon_reg[4]_i_1 
       (.I0(p_1_in[2]),
        .I1(\round_ctr_reg_reg[0]_rep_n_0 ),
        .I2(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I3(\rcon_reg_reg[7]_0 [3]),
        .I4(\rcon_reg_reg[7]_0 [7]),
        .O(rcon_new[4]));
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT4 #(
    .INIT(16'hD000)) 
    \rcon_reg[5]_i_1 
       (.I0(p_1_in[2]),
        .I1(\round_ctr_reg_reg[0]_rep_n_0 ),
        .I2(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I3(\rcon_reg_reg[7]_0 [4]),
        .O(rcon_new[5]));
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT4 #(
    .INIT(16'hD000)) 
    \rcon_reg[6]_i_1 
       (.I0(p_1_in[2]),
        .I1(\round_ctr_reg_reg[0]_rep_n_0 ),
        .I2(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I3(\rcon_reg_reg[7]_0 [5]),
        .O(rcon_new[6]));
  LUT3 #(
    .INIT(8'hDF)) 
    \rcon_reg[7]_i_1 
       (.I0(p_1_in[2]),
        .I1(\round_ctr_reg_reg[0]_rep_n_0 ),
        .I2(\round_ctr_reg[3]_i_3__1_n_0 ),
        .O(\rcon_reg[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT4 #(
    .INIT(16'hB3BB)) 
    \rcon_reg[7]_i_2 
       (.I0(\rcon_reg_reg[7]_0 [6]),
        .I1(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I2(\round_ctr_reg_reg[0]_rep_n_0 ),
        .I3(p_1_in[2]),
        .O(rcon_new[7]));
  FDCE #(
    .INIT(1'b0)) 
    \rcon_reg_reg[0] 
       (.C(clk_i),
        .CE(\rcon_reg[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(rcon_new[0]),
        .Q(\rcon_reg_reg[7]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \rcon_reg_reg[1] 
       (.C(clk_i),
        .CE(\rcon_reg[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(rcon_new[1]),
        .Q(\rcon_reg_reg[7]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \rcon_reg_reg[2] 
       (.C(clk_i),
        .CE(\rcon_reg[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(rcon_new[2]),
        .Q(\rcon_reg_reg[7]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \rcon_reg_reg[3] 
       (.C(clk_i),
        .CE(\rcon_reg[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(rcon_new[3]),
        .Q(\rcon_reg_reg[7]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \rcon_reg_reg[4] 
       (.C(clk_i),
        .CE(\rcon_reg[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(rcon_new[4]),
        .Q(\rcon_reg_reg[7]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \rcon_reg_reg[5] 
       (.C(clk_i),
        .CE(\rcon_reg[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(rcon_new[5]),
        .Q(\rcon_reg_reg[7]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \rcon_reg_reg[6] 
       (.C(clk_i),
        .CE(\rcon_reg[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(rcon_new[6]),
        .Q(\rcon_reg_reg[7]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \rcon_reg_reg[7] 
       (.C(clk_i),
        .CE(\rcon_reg[7]_i_1_n_0 ),
        .CLR(rst_i),
        .D(rcon_new[7]),
        .Q(\rcon_reg_reg[7]_0 [7]));
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT4 #(
    .INIT(16'hFBA0)) 
    ready_reg_i_1__1
       (.I0(key_mem_ctrl_reg[0]),
        .I1(p_1_in[0]),
        .I2(key_mem_ctrl_reg[1]),
        .I3(key_ready),
        .O(ready_reg_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h3033300088888888)) 
    ready_reg_i_1__2
       (.I0(key_ready),
        .I1(ready_reg_reg_0[0]),
        .I2(enc_ready),
        .I3(p_1_in[1]),
        .I4(dec_ready),
        .I5(ready_reg_reg_0[1]),
        .O(ready_new));
  FDCE #(
    .INIT(1'b0)) 
    ready_reg_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(ready_reg_i_1__1_n_0),
        .Q(key_ready));
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT4 #(
    .INIT(16'h4044)) 
    \round_ctr_reg[0]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[0] ),
        .I1(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I2(key_mem_ctrl_reg[1]),
        .I3(key_mem_ctrl_reg[0]),
        .O(round_ctr_new[0]));
  LUT4 #(
    .INIT(16'h4044)) 
    \round_ctr_reg[0]_rep_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[0] ),
        .I1(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I2(key_mem_ctrl_reg[1]),
        .I3(key_mem_ctrl_reg[0]),
        .O(\round_ctr_reg[0]_rep_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h4044)) 
    \round_ctr_reg[0]_rep_i_1__0 
       (.I0(\round_ctr_reg_reg_n_0_[0] ),
        .I1(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I2(key_mem_ctrl_reg[1]),
        .I3(key_mem_ctrl_reg[0]),
        .O(\round_ctr_reg[0]_rep_i_1__0_n_0 ));
  LUT4 #(
    .INIT(16'h4044)) 
    \round_ctr_reg[0]_rep_i_1__1 
       (.I0(\round_ctr_reg_reg_n_0_[0] ),
        .I1(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I2(key_mem_ctrl_reg[1]),
        .I3(key_mem_ctrl_reg[0]),
        .O(\round_ctr_reg[0]_rep_i_1__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT5 #(
    .INIT(32'h60006060)) 
    \round_ctr_reg[1]_i_1 
       (.I0(\round_ctr_reg_reg_n_0_[0] ),
        .I1(p_0_in0),
        .I2(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I3(key_mem_ctrl_reg[1]),
        .I4(key_mem_ctrl_reg[0]),
        .O(round_ctr_new[1]));
  LUT6 #(
    .INIT(64'h7800000078007800)) 
    \round_ctr_reg[2]_i_1 
       (.I0(p_0_in0),
        .I1(\round_ctr_reg_reg_n_0_[0] ),
        .I2(\round_ctr_reg_reg_n_0_[2] ),
        .I3(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I4(key_mem_ctrl_reg[1]),
        .I5(key_mem_ctrl_reg[0]),
        .O(round_ctr_new[2]));
  LUT3 #(
    .INIT(8'hF4)) 
    \round_ctr_reg[3]_i_1 
       (.I0(key_mem_ctrl_reg[1]),
        .I1(key_mem_ctrl_reg[0]),
        .I2(\round_ctr_reg[3]_i_3__1_n_0 ),
        .O(round_ctr_we));
  LUT6 #(
    .INIT(64'h000000007F800000)) 
    \round_ctr_reg[3]_i_2 
       (.I0(\round_ctr_reg_reg_n_0_[0] ),
        .I1(p_0_in0),
        .I2(\round_ctr_reg_reg_n_0_[2] ),
        .I3(\round_ctr_reg_reg_n_0_[3] ),
        .I4(\round_ctr_reg[3]_i_3__1_n_0 ),
        .I5(\round_ctr_reg[3]_i_4__0_n_0 ),
        .O(round_ctr_new[3]));
  LUT2 #(
    .INIT(4'h2)) 
    \round_ctr_reg[3]_i_3__1 
       (.I0(key_mem_ctrl_reg[1]),
        .I1(key_mem_ctrl_reg[0]),
        .O(\round_ctr_reg[3]_i_3__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \round_ctr_reg[3]_i_4__0 
       (.I0(key_mem_ctrl_reg[0]),
        .I1(key_mem_ctrl_reg[1]),
        .O(\round_ctr_reg[3]_i_4__0_n_0 ));
  (* ORIG_CELL_NAME = "round_ctr_reg_reg[0]" *) 
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[0] 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(round_ctr_new[0]),
        .Q(\round_ctr_reg_reg_n_0_[0] ));
  (* ORIG_CELL_NAME = "round_ctr_reg_reg[0]" *) 
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[0]_rep 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(\round_ctr_reg[0]_rep_i_1_n_0 ),
        .Q(\round_ctr_reg_reg[0]_rep_n_0 ));
  (* ORIG_CELL_NAME = "round_ctr_reg_reg[0]" *) 
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[0]_rep__0 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(\round_ctr_reg[0]_rep_i_1__0_n_0 ),
        .Q(\round_ctr_reg_reg[0]_rep__0_n_0 ));
  (* ORIG_CELL_NAME = "round_ctr_reg_reg[0]" *) 
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[0]_rep__1 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(\round_ctr_reg[0]_rep_i_1__1_n_0 ),
        .Q(\round_ctr_reg_reg[0]_rep__1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[1] 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(round_ctr_new[1]),
        .Q(p_0_in0));
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[2] 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(round_ctr_new[2]),
        .Q(\round_ctr_reg_reg_n_0_[2] ));
  FDCE #(
    .INIT(1'b0)) 
    \round_ctr_reg_reg[3] 
       (.C(clk_i),
        .CE(round_ctr_we),
        .CLR(rst_i),
        .D(round_ctr_new[3]),
        .Q(\round_ctr_reg_reg_n_0_[3] ));
endmodule

(* ORIG_REF_NAME = "aes_sbox" *) 
module switch_elements_aes_sbox
   (new_sboxw,
    \block_w3_reg[31]_i_3 ,
    \block_w2_reg_reg[0]_i_5_0 ,
    \block_w2_reg_reg[0]_i_5_1 ,
    \block_w2_reg_reg[0]_i_5_2 ,
    \block_w2_reg_reg[0]_i_5_3 ,
    \block_w2_reg_reg[1]_i_5_0 ,
    \block_w2_reg_reg[1]_i_5_1 ,
    \block_w2_reg_reg[1]_i_5_2 ,
    \block_w2_reg_reg[1]_i_5_3 ,
    \block_w2_reg_reg[2]_i_5_0 ,
    \block_w2_reg_reg[2]_i_5_1 ,
    \block_w2_reg_reg[2]_i_5_2 ,
    \block_w2_reg_reg[2]_i_5_3 ,
    \block_w2_reg_reg[3]_i_5_0 ,
    \block_w2_reg_reg[3]_i_5_1 ,
    \block_w2_reg_reg[3]_i_5_2 ,
    \block_w2_reg_reg[3]_i_5_3 ,
    \block_w2_reg_reg[4]_i_6_0 ,
    \block_w2_reg_reg[4]_i_6_1 ,
    \block_w2_reg_reg[4]_i_6_2 ,
    \block_w2_reg_reg[4]_i_6_3 ,
    \block_w2_reg_reg[5]_i_5_0 ,
    \block_w2_reg_reg[5]_i_5_1 ,
    \block_w2_reg_reg[5]_i_5_2 ,
    \block_w2_reg_reg[5]_i_5_3 ,
    \block_w2_reg_reg[6]_i_5_0 ,
    \block_w2_reg_reg[6]_i_5_1 ,
    \block_w2_reg_reg[6]_i_5_2 ,
    \block_w2_reg_reg[6]_i_5_3 ,
    \block_w2_reg_reg[7]_i_5_0 ,
    \block_w2_reg_reg[7]_i_5_1 ,
    \block_w2_reg_reg[7]_i_5_2 ,
    \block_w2_reg_reg[7]_i_5_3 ,
    \sbox_inferred__0/block_w2_reg_reg[8]_i_5_0 ,
    \sbox_inferred__0/block_w2_reg_reg[8]_i_5_1 ,
    \sbox_inferred__0/block_w2_reg_reg[8]_i_5_2 ,
    \sbox_inferred__0/block_w2_reg_reg[8]_i_5_3 ,
    \sbox_inferred__0/block_w2_reg_reg[9]_i_6_0 ,
    \sbox_inferred__0/block_w2_reg_reg[9]_i_6_1 ,
    \sbox_inferred__0/block_w2_reg_reg[9]_i_6_2 ,
    \sbox_inferred__0/block_w2_reg_reg[9]_i_6_3 ,
    \sbox_inferred__0/block_w2_reg_reg[10]_i_5_0 ,
    \sbox_inferred__0/block_w2_reg_reg[10]_i_5_1 ,
    \sbox_inferred__0/block_w2_reg_reg[10]_i_5_2 ,
    \sbox_inferred__0/block_w2_reg_reg[10]_i_5_3 ,
    \sbox_inferred__0/block_w2_reg_reg[11]_i_5_0 ,
    \sbox_inferred__0/block_w2_reg_reg[11]_i_5_1 ,
    \sbox_inferred__0/block_w2_reg_reg[11]_i_5_2 ,
    \sbox_inferred__0/block_w2_reg_reg[11]_i_5_3 ,
    \sbox_inferred__0/block_w2_reg_reg[12]_i_5_0 ,
    \sbox_inferred__0/block_w2_reg_reg[12]_i_5_1 ,
    \sbox_inferred__0/block_w2_reg_reg[12]_i_5_2 ,
    \sbox_inferred__0/block_w2_reg_reg[12]_i_5_3 ,
    \sbox_inferred__0/block_w2_reg_reg[13]_i_5_0 ,
    \sbox_inferred__0/block_w2_reg_reg[13]_i_5_1 ,
    \sbox_inferred__0/block_w2_reg_reg[13]_i_5_2 ,
    \sbox_inferred__0/block_w2_reg_reg[13]_i_5_3 ,
    \sbox_inferred__0/block_w2_reg_reg[14]_i_5_0 ,
    \sbox_inferred__0/block_w2_reg_reg[14]_i_5_1 ,
    \sbox_inferred__0/block_w2_reg_reg[14]_i_5_2 ,
    \sbox_inferred__0/block_w2_reg_reg[14]_i_5_3 ,
    \sbox_inferred__0/block_w2_reg_reg[15]_i_5_0 ,
    \sbox_inferred__0/block_w2_reg_reg[15]_i_5_1 ,
    \sbox_inferred__0/block_w2_reg_reg[15]_i_5_2 ,
    \sbox_inferred__0/block_w2_reg_reg[15]_i_5_3 ,
    \sbox_inferred__1/block_w2_reg_reg[16]_i_5_0 ,
    \sbox_inferred__1/block_w2_reg_reg[16]_i_5_1 ,
    \sbox_inferred__1/block_w2_reg_reg[16]_i_5_2 ,
    \sbox_inferred__1/block_w2_reg_reg[16]_i_5_3 ,
    \sbox_inferred__1/block_w2_reg_reg[17]_i_5_0 ,
    \sbox_inferred__1/block_w2_reg_reg[17]_i_5_1 ,
    \sbox_inferred__1/block_w2_reg_reg[17]_i_5_2 ,
    \sbox_inferred__1/block_w2_reg_reg[17]_i_5_3 ,
    \sbox_inferred__1/block_w2_reg_reg[18]_i_5_0 ,
    \sbox_inferred__1/block_w2_reg_reg[18]_i_5_1 ,
    \sbox_inferred__1/block_w2_reg_reg[18]_i_5_2 ,
    \sbox_inferred__1/block_w2_reg_reg[18]_i_5_3 ,
    \sbox_inferred__1/block_w2_reg_reg[19]_i_5_0 ,
    \sbox_inferred__1/block_w2_reg_reg[19]_i_5_1 ,
    \sbox_inferred__1/block_w2_reg_reg[19]_i_5_2 ,
    \sbox_inferred__1/block_w2_reg_reg[19]_i_5_3 ,
    \sbox_inferred__1/block_w2_reg_reg[20]_i_6_0 ,
    \sbox_inferred__1/block_w2_reg_reg[20]_i_6_1 ,
    \sbox_inferred__1/block_w2_reg_reg[20]_i_6_2 ,
    \sbox_inferred__1/block_w2_reg_reg[20]_i_6_3 ,
    \sbox_inferred__1/block_w2_reg_reg[21]_i_5_0 ,
    \sbox_inferred__1/block_w2_reg_reg[21]_i_5_1 ,
    \sbox_inferred__1/block_w2_reg_reg[21]_i_5_2 ,
    \sbox_inferred__1/block_w2_reg_reg[21]_i_5_3 ,
    \sbox_inferred__1/block_w2_reg_reg[22]_i_5_0 ,
    \sbox_inferred__1/block_w2_reg_reg[22]_i_5_1 ,
    \sbox_inferred__1/block_w2_reg_reg[22]_i_5_2 ,
    \sbox_inferred__1/block_w2_reg_reg[22]_i_5_3 ,
    \sbox_inferred__1/block_w2_reg_reg[23]_i_5_0 ,
    \sbox_inferred__1/block_w2_reg_reg[23]_i_5_1 ,
    \sbox_inferred__1/block_w2_reg_reg[23]_i_5_2 ,
    \sbox_inferred__1/block_w2_reg_reg[23]_i_5_3 ,
    \sbox_inferred__2/block_w2_reg_reg[24]_i_5_0 ,
    \sbox_inferred__2/block_w2_reg_reg[24]_i_5_1 ,
    \sbox_inferred__2/block_w2_reg_reg[24]_i_5_2 ,
    \sbox_inferred__2/block_w2_reg_reg[24]_i_5_3 ,
    \sbox_inferred__2/block_w2_reg_reg[25]_i_6_0 ,
    \sbox_inferred__2/block_w2_reg_reg[25]_i_6_1 ,
    \sbox_inferred__2/block_w2_reg_reg[25]_i_6_2 ,
    \sbox_inferred__2/block_w2_reg_reg[25]_i_6_3 ,
    \sbox_inferred__2/block_w2_reg_reg[26]_i_5_0 ,
    \sbox_inferred__2/block_w2_reg_reg[26]_i_5_1 ,
    \sbox_inferred__2/block_w2_reg_reg[26]_i_5_2 ,
    \sbox_inferred__2/block_w2_reg_reg[26]_i_5_3 ,
    \sbox_inferred__2/block_w2_reg_reg[27]_i_5_0 ,
    \sbox_inferred__2/block_w2_reg_reg[27]_i_5_1 ,
    \sbox_inferred__2/block_w2_reg_reg[27]_i_5_2 ,
    \sbox_inferred__2/block_w2_reg_reg[27]_i_5_3 ,
    \sbox_inferred__2/block_w2_reg_reg[28]_i_5_0 ,
    \sbox_inferred__2/block_w2_reg_reg[28]_i_5_1 ,
    \sbox_inferred__2/block_w2_reg_reg[28]_i_5_2 ,
    \sbox_inferred__2/block_w2_reg_reg[28]_i_5_3 ,
    \sbox_inferred__2/block_w2_reg_reg[29]_i_5_0 ,
    \sbox_inferred__2/block_w2_reg_reg[29]_i_5_1 ,
    \sbox_inferred__2/block_w2_reg_reg[29]_i_5_2 ,
    \sbox_inferred__2/block_w2_reg_reg[29]_i_5_3 ,
    \sbox_inferred__2/block_w2_reg_reg[30]_i_5_0 ,
    \sbox_inferred__2/block_w2_reg_reg[30]_i_5_1 ,
    \sbox_inferred__2/block_w2_reg_reg[30]_i_5_2 ,
    \sbox_inferred__2/block_w2_reg_reg[30]_i_5_3 ,
    \sbox_inferred__2/block_w2_reg_reg[31]_i_10_0 ,
    \sbox_inferred__2/block_w2_reg_reg[31]_i_10_1 ,
    \sbox_inferred__2/block_w2_reg_reg[31]_i_10_2 ,
    \sbox_inferred__2/block_w2_reg_reg[31]_i_10_3 );
  output [31:0]new_sboxw;
  input [7:0]\block_w3_reg[31]_i_3 ;
  input \block_w2_reg_reg[0]_i_5_0 ;
  input \block_w2_reg_reg[0]_i_5_1 ;
  input \block_w2_reg_reg[0]_i_5_2 ;
  input \block_w2_reg_reg[0]_i_5_3 ;
  input \block_w2_reg_reg[1]_i_5_0 ;
  input \block_w2_reg_reg[1]_i_5_1 ;
  input \block_w2_reg_reg[1]_i_5_2 ;
  input \block_w2_reg_reg[1]_i_5_3 ;
  input \block_w2_reg_reg[2]_i_5_0 ;
  input \block_w2_reg_reg[2]_i_5_1 ;
  input \block_w2_reg_reg[2]_i_5_2 ;
  input \block_w2_reg_reg[2]_i_5_3 ;
  input \block_w2_reg_reg[3]_i_5_0 ;
  input \block_w2_reg_reg[3]_i_5_1 ;
  input \block_w2_reg_reg[3]_i_5_2 ;
  input \block_w2_reg_reg[3]_i_5_3 ;
  input \block_w2_reg_reg[4]_i_6_0 ;
  input \block_w2_reg_reg[4]_i_6_1 ;
  input \block_w2_reg_reg[4]_i_6_2 ;
  input \block_w2_reg_reg[4]_i_6_3 ;
  input \block_w2_reg_reg[5]_i_5_0 ;
  input \block_w2_reg_reg[5]_i_5_1 ;
  input \block_w2_reg_reg[5]_i_5_2 ;
  input \block_w2_reg_reg[5]_i_5_3 ;
  input \block_w2_reg_reg[6]_i_5_0 ;
  input \block_w2_reg_reg[6]_i_5_1 ;
  input \block_w2_reg_reg[6]_i_5_2 ;
  input \block_w2_reg_reg[6]_i_5_3 ;
  input \block_w2_reg_reg[7]_i_5_0 ;
  input \block_w2_reg_reg[7]_i_5_1 ;
  input \block_w2_reg_reg[7]_i_5_2 ;
  input \block_w2_reg_reg[7]_i_5_3 ;
  input \sbox_inferred__0/block_w2_reg_reg[8]_i_5_0 ;
  input \sbox_inferred__0/block_w2_reg_reg[8]_i_5_1 ;
  input \sbox_inferred__0/block_w2_reg_reg[8]_i_5_2 ;
  input \sbox_inferred__0/block_w2_reg_reg[8]_i_5_3 ;
  input \sbox_inferred__0/block_w2_reg_reg[9]_i_6_0 ;
  input \sbox_inferred__0/block_w2_reg_reg[9]_i_6_1 ;
  input \sbox_inferred__0/block_w2_reg_reg[9]_i_6_2 ;
  input \sbox_inferred__0/block_w2_reg_reg[9]_i_6_3 ;
  input \sbox_inferred__0/block_w2_reg_reg[10]_i_5_0 ;
  input \sbox_inferred__0/block_w2_reg_reg[10]_i_5_1 ;
  input \sbox_inferred__0/block_w2_reg_reg[10]_i_5_2 ;
  input \sbox_inferred__0/block_w2_reg_reg[10]_i_5_3 ;
  input \sbox_inferred__0/block_w2_reg_reg[11]_i_5_0 ;
  input \sbox_inferred__0/block_w2_reg_reg[11]_i_5_1 ;
  input \sbox_inferred__0/block_w2_reg_reg[11]_i_5_2 ;
  input \sbox_inferred__0/block_w2_reg_reg[11]_i_5_3 ;
  input \sbox_inferred__0/block_w2_reg_reg[12]_i_5_0 ;
  input \sbox_inferred__0/block_w2_reg_reg[12]_i_5_1 ;
  input \sbox_inferred__0/block_w2_reg_reg[12]_i_5_2 ;
  input \sbox_inferred__0/block_w2_reg_reg[12]_i_5_3 ;
  input \sbox_inferred__0/block_w2_reg_reg[13]_i_5_0 ;
  input \sbox_inferred__0/block_w2_reg_reg[13]_i_5_1 ;
  input \sbox_inferred__0/block_w2_reg_reg[13]_i_5_2 ;
  input \sbox_inferred__0/block_w2_reg_reg[13]_i_5_3 ;
  input \sbox_inferred__0/block_w2_reg_reg[14]_i_5_0 ;
  input \sbox_inferred__0/block_w2_reg_reg[14]_i_5_1 ;
  input \sbox_inferred__0/block_w2_reg_reg[14]_i_5_2 ;
  input \sbox_inferred__0/block_w2_reg_reg[14]_i_5_3 ;
  input \sbox_inferred__0/block_w2_reg_reg[15]_i_5_0 ;
  input \sbox_inferred__0/block_w2_reg_reg[15]_i_5_1 ;
  input \sbox_inferred__0/block_w2_reg_reg[15]_i_5_2 ;
  input \sbox_inferred__0/block_w2_reg_reg[15]_i_5_3 ;
  input \sbox_inferred__1/block_w2_reg_reg[16]_i_5_0 ;
  input \sbox_inferred__1/block_w2_reg_reg[16]_i_5_1 ;
  input \sbox_inferred__1/block_w2_reg_reg[16]_i_5_2 ;
  input \sbox_inferred__1/block_w2_reg_reg[16]_i_5_3 ;
  input \sbox_inferred__1/block_w2_reg_reg[17]_i_5_0 ;
  input \sbox_inferred__1/block_w2_reg_reg[17]_i_5_1 ;
  input \sbox_inferred__1/block_w2_reg_reg[17]_i_5_2 ;
  input \sbox_inferred__1/block_w2_reg_reg[17]_i_5_3 ;
  input \sbox_inferred__1/block_w2_reg_reg[18]_i_5_0 ;
  input \sbox_inferred__1/block_w2_reg_reg[18]_i_5_1 ;
  input \sbox_inferred__1/block_w2_reg_reg[18]_i_5_2 ;
  input \sbox_inferred__1/block_w2_reg_reg[18]_i_5_3 ;
  input \sbox_inferred__1/block_w2_reg_reg[19]_i_5_0 ;
  input \sbox_inferred__1/block_w2_reg_reg[19]_i_5_1 ;
  input \sbox_inferred__1/block_w2_reg_reg[19]_i_5_2 ;
  input \sbox_inferred__1/block_w2_reg_reg[19]_i_5_3 ;
  input \sbox_inferred__1/block_w2_reg_reg[20]_i_6_0 ;
  input \sbox_inferred__1/block_w2_reg_reg[20]_i_6_1 ;
  input \sbox_inferred__1/block_w2_reg_reg[20]_i_6_2 ;
  input \sbox_inferred__1/block_w2_reg_reg[20]_i_6_3 ;
  input \sbox_inferred__1/block_w2_reg_reg[21]_i_5_0 ;
  input \sbox_inferred__1/block_w2_reg_reg[21]_i_5_1 ;
  input \sbox_inferred__1/block_w2_reg_reg[21]_i_5_2 ;
  input \sbox_inferred__1/block_w2_reg_reg[21]_i_5_3 ;
  input \sbox_inferred__1/block_w2_reg_reg[22]_i_5_0 ;
  input \sbox_inferred__1/block_w2_reg_reg[22]_i_5_1 ;
  input \sbox_inferred__1/block_w2_reg_reg[22]_i_5_2 ;
  input \sbox_inferred__1/block_w2_reg_reg[22]_i_5_3 ;
  input \sbox_inferred__1/block_w2_reg_reg[23]_i_5_0 ;
  input \sbox_inferred__1/block_w2_reg_reg[23]_i_5_1 ;
  input \sbox_inferred__1/block_w2_reg_reg[23]_i_5_2 ;
  input \sbox_inferred__1/block_w2_reg_reg[23]_i_5_3 ;
  input \sbox_inferred__2/block_w2_reg_reg[24]_i_5_0 ;
  input \sbox_inferred__2/block_w2_reg_reg[24]_i_5_1 ;
  input \sbox_inferred__2/block_w2_reg_reg[24]_i_5_2 ;
  input \sbox_inferred__2/block_w2_reg_reg[24]_i_5_3 ;
  input \sbox_inferred__2/block_w2_reg_reg[25]_i_6_0 ;
  input \sbox_inferred__2/block_w2_reg_reg[25]_i_6_1 ;
  input \sbox_inferred__2/block_w2_reg_reg[25]_i_6_2 ;
  input \sbox_inferred__2/block_w2_reg_reg[25]_i_6_3 ;
  input \sbox_inferred__2/block_w2_reg_reg[26]_i_5_0 ;
  input \sbox_inferred__2/block_w2_reg_reg[26]_i_5_1 ;
  input \sbox_inferred__2/block_w2_reg_reg[26]_i_5_2 ;
  input \sbox_inferred__2/block_w2_reg_reg[26]_i_5_3 ;
  input \sbox_inferred__2/block_w2_reg_reg[27]_i_5_0 ;
  input \sbox_inferred__2/block_w2_reg_reg[27]_i_5_1 ;
  input \sbox_inferred__2/block_w2_reg_reg[27]_i_5_2 ;
  input \sbox_inferred__2/block_w2_reg_reg[27]_i_5_3 ;
  input \sbox_inferred__2/block_w2_reg_reg[28]_i_5_0 ;
  input \sbox_inferred__2/block_w2_reg_reg[28]_i_5_1 ;
  input \sbox_inferred__2/block_w2_reg_reg[28]_i_5_2 ;
  input \sbox_inferred__2/block_w2_reg_reg[28]_i_5_3 ;
  input \sbox_inferred__2/block_w2_reg_reg[29]_i_5_0 ;
  input \sbox_inferred__2/block_w2_reg_reg[29]_i_5_1 ;
  input \sbox_inferred__2/block_w2_reg_reg[29]_i_5_2 ;
  input \sbox_inferred__2/block_w2_reg_reg[29]_i_5_3 ;
  input \sbox_inferred__2/block_w2_reg_reg[30]_i_5_0 ;
  input \sbox_inferred__2/block_w2_reg_reg[30]_i_5_1 ;
  input \sbox_inferred__2/block_w2_reg_reg[30]_i_5_2 ;
  input \sbox_inferred__2/block_w2_reg_reg[30]_i_5_3 ;
  input \sbox_inferred__2/block_w2_reg_reg[31]_i_10_0 ;
  input \sbox_inferred__2/block_w2_reg_reg[31]_i_10_1 ;
  input \sbox_inferred__2/block_w2_reg_reg[31]_i_10_2 ;
  input \sbox_inferred__2/block_w2_reg_reg[31]_i_10_3 ;

  wire \block_w2_reg_reg[0]_i_10_n_0 ;
  wire \block_w2_reg_reg[0]_i_5_0 ;
  wire \block_w2_reg_reg[0]_i_5_1 ;
  wire \block_w2_reg_reg[0]_i_5_2 ;
  wire \block_w2_reg_reg[0]_i_5_3 ;
  wire \block_w2_reg_reg[0]_i_9_n_0 ;
  wire \block_w2_reg_reg[1]_i_10_n_0 ;
  wire \block_w2_reg_reg[1]_i_11_n_0 ;
  wire \block_w2_reg_reg[1]_i_5_0 ;
  wire \block_w2_reg_reg[1]_i_5_1 ;
  wire \block_w2_reg_reg[1]_i_5_2 ;
  wire \block_w2_reg_reg[1]_i_5_3 ;
  wire \block_w2_reg_reg[2]_i_10_n_0 ;
  wire \block_w2_reg_reg[2]_i_5_0 ;
  wire \block_w2_reg_reg[2]_i_5_1 ;
  wire \block_w2_reg_reg[2]_i_5_2 ;
  wire \block_w2_reg_reg[2]_i_5_3 ;
  wire \block_w2_reg_reg[2]_i_9_n_0 ;
  wire \block_w2_reg_reg[3]_i_10_n_0 ;
  wire \block_w2_reg_reg[3]_i_11_n_0 ;
  wire \block_w2_reg_reg[3]_i_5_0 ;
  wire \block_w2_reg_reg[3]_i_5_1 ;
  wire \block_w2_reg_reg[3]_i_5_2 ;
  wire \block_w2_reg_reg[3]_i_5_3 ;
  wire \block_w2_reg_reg[4]_i_11_n_0 ;
  wire \block_w2_reg_reg[4]_i_12_n_0 ;
  wire \block_w2_reg_reg[4]_i_6_0 ;
  wire \block_w2_reg_reg[4]_i_6_1 ;
  wire \block_w2_reg_reg[4]_i_6_2 ;
  wire \block_w2_reg_reg[4]_i_6_3 ;
  wire \block_w2_reg_reg[5]_i_10_n_0 ;
  wire \block_w2_reg_reg[5]_i_5_0 ;
  wire \block_w2_reg_reg[5]_i_5_1 ;
  wire \block_w2_reg_reg[5]_i_5_2 ;
  wire \block_w2_reg_reg[5]_i_5_3 ;
  wire \block_w2_reg_reg[5]_i_9_n_0 ;
  wire \block_w2_reg_reg[6]_i_10_n_0 ;
  wire \block_w2_reg_reg[6]_i_5_0 ;
  wire \block_w2_reg_reg[6]_i_5_1 ;
  wire \block_w2_reg_reg[6]_i_5_2 ;
  wire \block_w2_reg_reg[6]_i_5_3 ;
  wire \block_w2_reg_reg[6]_i_9_n_0 ;
  wire \block_w2_reg_reg[7]_i_10_n_0 ;
  wire \block_w2_reg_reg[7]_i_11_n_0 ;
  wire \block_w2_reg_reg[7]_i_5_0 ;
  wire \block_w2_reg_reg[7]_i_5_1 ;
  wire \block_w2_reg_reg[7]_i_5_2 ;
  wire \block_w2_reg_reg[7]_i_5_3 ;
  wire [7:0]\block_w3_reg[31]_i_3 ;
  wire [31:0]new_sboxw;
  wire \sbox_inferred__0/block_w2_reg_reg[10]_i_10_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[10]_i_5_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[10]_i_5_1 ;
  wire \sbox_inferred__0/block_w2_reg_reg[10]_i_5_2 ;
  wire \sbox_inferred__0/block_w2_reg_reg[10]_i_5_3 ;
  wire \sbox_inferred__0/block_w2_reg_reg[10]_i_9_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[11]_i_10_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[11]_i_11_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[11]_i_5_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[11]_i_5_1 ;
  wire \sbox_inferred__0/block_w2_reg_reg[11]_i_5_2 ;
  wire \sbox_inferred__0/block_w2_reg_reg[11]_i_5_3 ;
  wire \sbox_inferred__0/block_w2_reg_reg[12]_i_10_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[12]_i_11_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[12]_i_5_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[12]_i_5_1 ;
  wire \sbox_inferred__0/block_w2_reg_reg[12]_i_5_2 ;
  wire \sbox_inferred__0/block_w2_reg_reg[12]_i_5_3 ;
  wire \sbox_inferred__0/block_w2_reg_reg[13]_i_10_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[13]_i_5_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[13]_i_5_1 ;
  wire \sbox_inferred__0/block_w2_reg_reg[13]_i_5_2 ;
  wire \sbox_inferred__0/block_w2_reg_reg[13]_i_5_3 ;
  wire \sbox_inferred__0/block_w2_reg_reg[13]_i_9_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[14]_i_10_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[14]_i_5_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[14]_i_5_1 ;
  wire \sbox_inferred__0/block_w2_reg_reg[14]_i_5_2 ;
  wire \sbox_inferred__0/block_w2_reg_reg[14]_i_5_3 ;
  wire \sbox_inferred__0/block_w2_reg_reg[14]_i_9_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[15]_i_10_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[15]_i_11_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[15]_i_5_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[15]_i_5_1 ;
  wire \sbox_inferred__0/block_w2_reg_reg[15]_i_5_2 ;
  wire \sbox_inferred__0/block_w2_reg_reg[15]_i_5_3 ;
  wire \sbox_inferred__0/block_w2_reg_reg[8]_i_10_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[8]_i_5_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[8]_i_5_1 ;
  wire \sbox_inferred__0/block_w2_reg_reg[8]_i_5_2 ;
  wire \sbox_inferred__0/block_w2_reg_reg[8]_i_5_3 ;
  wire \sbox_inferred__0/block_w2_reg_reg[8]_i_9_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[9]_i_11_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[9]_i_12_n_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[9]_i_6_0 ;
  wire \sbox_inferred__0/block_w2_reg_reg[9]_i_6_1 ;
  wire \sbox_inferred__0/block_w2_reg_reg[9]_i_6_2 ;
  wire \sbox_inferred__0/block_w2_reg_reg[9]_i_6_3 ;
  wire \sbox_inferred__1/block_w2_reg_reg[16]_i_10_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[16]_i_5_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[16]_i_5_1 ;
  wire \sbox_inferred__1/block_w2_reg_reg[16]_i_5_2 ;
  wire \sbox_inferred__1/block_w2_reg_reg[16]_i_5_3 ;
  wire \sbox_inferred__1/block_w2_reg_reg[16]_i_9_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[17]_i_10_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[17]_i_11_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[17]_i_5_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[17]_i_5_1 ;
  wire \sbox_inferred__1/block_w2_reg_reg[17]_i_5_2 ;
  wire \sbox_inferred__1/block_w2_reg_reg[17]_i_5_3 ;
  wire \sbox_inferred__1/block_w2_reg_reg[18]_i_10_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[18]_i_5_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[18]_i_5_1 ;
  wire \sbox_inferred__1/block_w2_reg_reg[18]_i_5_2 ;
  wire \sbox_inferred__1/block_w2_reg_reg[18]_i_5_3 ;
  wire \sbox_inferred__1/block_w2_reg_reg[18]_i_9_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[19]_i_10_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[19]_i_11_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[19]_i_5_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[19]_i_5_1 ;
  wire \sbox_inferred__1/block_w2_reg_reg[19]_i_5_2 ;
  wire \sbox_inferred__1/block_w2_reg_reg[19]_i_5_3 ;
  wire \sbox_inferred__1/block_w2_reg_reg[20]_i_11_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[20]_i_12_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[20]_i_6_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[20]_i_6_1 ;
  wire \sbox_inferred__1/block_w2_reg_reg[20]_i_6_2 ;
  wire \sbox_inferred__1/block_w2_reg_reg[20]_i_6_3 ;
  wire \sbox_inferred__1/block_w2_reg_reg[21]_i_10_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[21]_i_5_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[21]_i_5_1 ;
  wire \sbox_inferred__1/block_w2_reg_reg[21]_i_5_2 ;
  wire \sbox_inferred__1/block_w2_reg_reg[21]_i_5_3 ;
  wire \sbox_inferred__1/block_w2_reg_reg[21]_i_9_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[22]_i_10_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[22]_i_5_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[22]_i_5_1 ;
  wire \sbox_inferred__1/block_w2_reg_reg[22]_i_5_2 ;
  wire \sbox_inferred__1/block_w2_reg_reg[22]_i_5_3 ;
  wire \sbox_inferred__1/block_w2_reg_reg[22]_i_9_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[23]_i_10_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[23]_i_11_n_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[23]_i_5_0 ;
  wire \sbox_inferred__1/block_w2_reg_reg[23]_i_5_1 ;
  wire \sbox_inferred__1/block_w2_reg_reg[23]_i_5_2 ;
  wire \sbox_inferred__1/block_w2_reg_reg[23]_i_5_3 ;
  wire \sbox_inferred__2/block_w2_reg_reg[24]_i_10_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[24]_i_5_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[24]_i_5_1 ;
  wire \sbox_inferred__2/block_w2_reg_reg[24]_i_5_2 ;
  wire \sbox_inferred__2/block_w2_reg_reg[24]_i_5_3 ;
  wire \sbox_inferred__2/block_w2_reg_reg[24]_i_9_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[25]_i_11_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[25]_i_12_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[25]_i_6_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[25]_i_6_1 ;
  wire \sbox_inferred__2/block_w2_reg_reg[25]_i_6_2 ;
  wire \sbox_inferred__2/block_w2_reg_reg[25]_i_6_3 ;
  wire \sbox_inferred__2/block_w2_reg_reg[26]_i_10_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[26]_i_5_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[26]_i_5_1 ;
  wire \sbox_inferred__2/block_w2_reg_reg[26]_i_5_2 ;
  wire \sbox_inferred__2/block_w2_reg_reg[26]_i_5_3 ;
  wire \sbox_inferred__2/block_w2_reg_reg[26]_i_9_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[27]_i_12_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[27]_i_13_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[27]_i_5_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[27]_i_5_1 ;
  wire \sbox_inferred__2/block_w2_reg_reg[27]_i_5_2 ;
  wire \sbox_inferred__2/block_w2_reg_reg[27]_i_5_3 ;
  wire \sbox_inferred__2/block_w2_reg_reg[28]_i_11_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[28]_i_12_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[28]_i_5_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[28]_i_5_1 ;
  wire \sbox_inferred__2/block_w2_reg_reg[28]_i_5_2 ;
  wire \sbox_inferred__2/block_w2_reg_reg[28]_i_5_3 ;
  wire \sbox_inferred__2/block_w2_reg_reg[29]_i_10_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[29]_i_5_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[29]_i_5_1 ;
  wire \sbox_inferred__2/block_w2_reg_reg[29]_i_5_2 ;
  wire \sbox_inferred__2/block_w2_reg_reg[29]_i_5_3 ;
  wire \sbox_inferred__2/block_w2_reg_reg[29]_i_9_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[30]_i_10_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[30]_i_5_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[30]_i_5_1 ;
  wire \sbox_inferred__2/block_w2_reg_reg[30]_i_5_2 ;
  wire \sbox_inferred__2/block_w2_reg_reg[30]_i_5_3 ;
  wire \sbox_inferred__2/block_w2_reg_reg[30]_i_9_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[31]_i_10_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[31]_i_10_1 ;
  wire \sbox_inferred__2/block_w2_reg_reg[31]_i_10_2 ;
  wire \sbox_inferred__2/block_w2_reg_reg[31]_i_10_3 ;
  wire \sbox_inferred__2/block_w2_reg_reg[31]_i_17_n_0 ;
  wire \sbox_inferred__2/block_w2_reg_reg[31]_i_18_n_0 ;

  MUXF7 \block_w2_reg_reg[0]_i_10 
       (.I0(\block_w2_reg_reg[0]_i_5_2 ),
        .I1(\block_w2_reg_reg[0]_i_5_3 ),
        .O(\block_w2_reg_reg[0]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF8 \block_w2_reg_reg[0]_i_5 
       (.I0(\block_w2_reg_reg[0]_i_9_n_0 ),
        .I1(\block_w2_reg_reg[0]_i_10_n_0 ),
        .O(new_sboxw[0]),
        .S(\block_w3_reg[31]_i_3 [1]));
  MUXF7 \block_w2_reg_reg[0]_i_9 
       (.I0(\block_w2_reg_reg[0]_i_5_0 ),
        .I1(\block_w2_reg_reg[0]_i_5_1 ),
        .O(\block_w2_reg_reg[0]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF7 \block_w2_reg_reg[1]_i_10 
       (.I0(\block_w2_reg_reg[1]_i_5_0 ),
        .I1(\block_w2_reg_reg[1]_i_5_1 ),
        .O(\block_w2_reg_reg[1]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF7 \block_w2_reg_reg[1]_i_11 
       (.I0(\block_w2_reg_reg[1]_i_5_2 ),
        .I1(\block_w2_reg_reg[1]_i_5_3 ),
        .O(\block_w2_reg_reg[1]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF8 \block_w2_reg_reg[1]_i_5 
       (.I0(\block_w2_reg_reg[1]_i_10_n_0 ),
        .I1(\block_w2_reg_reg[1]_i_11_n_0 ),
        .O(new_sboxw[1]),
        .S(\block_w3_reg[31]_i_3 [1]));
  MUXF7 \block_w2_reg_reg[2]_i_10 
       (.I0(\block_w2_reg_reg[2]_i_5_2 ),
        .I1(\block_w2_reg_reg[2]_i_5_3 ),
        .O(\block_w2_reg_reg[2]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF8 \block_w2_reg_reg[2]_i_5 
       (.I0(\block_w2_reg_reg[2]_i_9_n_0 ),
        .I1(\block_w2_reg_reg[2]_i_10_n_0 ),
        .O(new_sboxw[2]),
        .S(\block_w3_reg[31]_i_3 [1]));
  MUXF7 \block_w2_reg_reg[2]_i_9 
       (.I0(\block_w2_reg_reg[2]_i_5_0 ),
        .I1(\block_w2_reg_reg[2]_i_5_1 ),
        .O(\block_w2_reg_reg[2]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF7 \block_w2_reg_reg[3]_i_10 
       (.I0(\block_w2_reg_reg[3]_i_5_0 ),
        .I1(\block_w2_reg_reg[3]_i_5_1 ),
        .O(\block_w2_reg_reg[3]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF7 \block_w2_reg_reg[3]_i_11 
       (.I0(\block_w2_reg_reg[3]_i_5_2 ),
        .I1(\block_w2_reg_reg[3]_i_5_3 ),
        .O(\block_w2_reg_reg[3]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF8 \block_w2_reg_reg[3]_i_5 
       (.I0(\block_w2_reg_reg[3]_i_10_n_0 ),
        .I1(\block_w2_reg_reg[3]_i_11_n_0 ),
        .O(new_sboxw[3]),
        .S(\block_w3_reg[31]_i_3 [1]));
  MUXF7 \block_w2_reg_reg[4]_i_11 
       (.I0(\block_w2_reg_reg[4]_i_6_0 ),
        .I1(\block_w2_reg_reg[4]_i_6_1 ),
        .O(\block_w2_reg_reg[4]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF7 \block_w2_reg_reg[4]_i_12 
       (.I0(\block_w2_reg_reg[4]_i_6_2 ),
        .I1(\block_w2_reg_reg[4]_i_6_3 ),
        .O(\block_w2_reg_reg[4]_i_12_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF8 \block_w2_reg_reg[4]_i_6 
       (.I0(\block_w2_reg_reg[4]_i_11_n_0 ),
        .I1(\block_w2_reg_reg[4]_i_12_n_0 ),
        .O(new_sboxw[4]),
        .S(\block_w3_reg[31]_i_3 [1]));
  MUXF7 \block_w2_reg_reg[5]_i_10 
       (.I0(\block_w2_reg_reg[5]_i_5_2 ),
        .I1(\block_w2_reg_reg[5]_i_5_3 ),
        .O(\block_w2_reg_reg[5]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF8 \block_w2_reg_reg[5]_i_5 
       (.I0(\block_w2_reg_reg[5]_i_9_n_0 ),
        .I1(\block_w2_reg_reg[5]_i_10_n_0 ),
        .O(new_sboxw[5]),
        .S(\block_w3_reg[31]_i_3 [1]));
  MUXF7 \block_w2_reg_reg[5]_i_9 
       (.I0(\block_w2_reg_reg[5]_i_5_0 ),
        .I1(\block_w2_reg_reg[5]_i_5_1 ),
        .O(\block_w2_reg_reg[5]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF7 \block_w2_reg_reg[6]_i_10 
       (.I0(\block_w2_reg_reg[6]_i_5_2 ),
        .I1(\block_w2_reg_reg[6]_i_5_3 ),
        .O(\block_w2_reg_reg[6]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF8 \block_w2_reg_reg[6]_i_5 
       (.I0(\block_w2_reg_reg[6]_i_9_n_0 ),
        .I1(\block_w2_reg_reg[6]_i_10_n_0 ),
        .O(new_sboxw[6]),
        .S(\block_w3_reg[31]_i_3 [1]));
  MUXF7 \block_w2_reg_reg[6]_i_9 
       (.I0(\block_w2_reg_reg[6]_i_5_0 ),
        .I1(\block_w2_reg_reg[6]_i_5_1 ),
        .O(\block_w2_reg_reg[6]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF7 \block_w2_reg_reg[7]_i_10 
       (.I0(\block_w2_reg_reg[7]_i_5_0 ),
        .I1(\block_w2_reg_reg[7]_i_5_1 ),
        .O(\block_w2_reg_reg[7]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF7 \block_w2_reg_reg[7]_i_11 
       (.I0(\block_w2_reg_reg[7]_i_5_2 ),
        .I1(\block_w2_reg_reg[7]_i_5_3 ),
        .O(\block_w2_reg_reg[7]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [0]));
  MUXF8 \block_w2_reg_reg[7]_i_5 
       (.I0(\block_w2_reg_reg[7]_i_10_n_0 ),
        .I1(\block_w2_reg_reg[7]_i_11_n_0 ),
        .O(new_sboxw[7]),
        .S(\block_w3_reg[31]_i_3 [1]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[10]_i_10 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[10]_i_5_2 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[10]_i_5_3 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[10]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF8 \sbox_inferred__0/block_w2_reg_reg[10]_i_5 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[10]_i_9_n_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[10]_i_10_n_0 ),
        .O(new_sboxw[10]),
        .S(\block_w3_reg[31]_i_3 [3]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[10]_i_9 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[10]_i_5_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[10]_i_5_1 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[10]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[11]_i_10 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[11]_i_5_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[11]_i_5_1 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[11]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[11]_i_11 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[11]_i_5_2 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[11]_i_5_3 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[11]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF8 \sbox_inferred__0/block_w2_reg_reg[11]_i_5 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[11]_i_10_n_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[11]_i_11_n_0 ),
        .O(new_sboxw[11]),
        .S(\block_w3_reg[31]_i_3 [3]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[12]_i_10 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[12]_i_5_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[12]_i_5_1 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[12]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[12]_i_11 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[12]_i_5_2 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[12]_i_5_3 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[12]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF8 \sbox_inferred__0/block_w2_reg_reg[12]_i_5 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[12]_i_10_n_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[12]_i_11_n_0 ),
        .O(new_sboxw[12]),
        .S(\block_w3_reg[31]_i_3 [3]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[13]_i_10 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[13]_i_5_2 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[13]_i_5_3 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[13]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF8 \sbox_inferred__0/block_w2_reg_reg[13]_i_5 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[13]_i_9_n_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[13]_i_10_n_0 ),
        .O(new_sboxw[13]),
        .S(\block_w3_reg[31]_i_3 [3]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[13]_i_9 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[13]_i_5_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[13]_i_5_1 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[13]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[14]_i_10 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[14]_i_5_2 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[14]_i_5_3 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[14]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF8 \sbox_inferred__0/block_w2_reg_reg[14]_i_5 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[14]_i_9_n_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[14]_i_10_n_0 ),
        .O(new_sboxw[14]),
        .S(\block_w3_reg[31]_i_3 [3]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[14]_i_9 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[14]_i_5_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[14]_i_5_1 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[14]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[15]_i_10 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[15]_i_5_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[15]_i_5_1 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[15]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[15]_i_11 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[15]_i_5_2 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[15]_i_5_3 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[15]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF8 \sbox_inferred__0/block_w2_reg_reg[15]_i_5 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[15]_i_10_n_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[15]_i_11_n_0 ),
        .O(new_sboxw[15]),
        .S(\block_w3_reg[31]_i_3 [3]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[8]_i_10 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[8]_i_5_2 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[8]_i_5_3 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[8]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF8 \sbox_inferred__0/block_w2_reg_reg[8]_i_5 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[8]_i_9_n_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[8]_i_10_n_0 ),
        .O(new_sboxw[8]),
        .S(\block_w3_reg[31]_i_3 [3]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[8]_i_9 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[8]_i_5_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[8]_i_5_1 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[8]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[9]_i_11 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[9]_i_6_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[9]_i_6_1 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[9]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF7 \sbox_inferred__0/block_w2_reg_reg[9]_i_12 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[9]_i_6_2 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[9]_i_6_3 ),
        .O(\sbox_inferred__0/block_w2_reg_reg[9]_i_12_n_0 ),
        .S(\block_w3_reg[31]_i_3 [2]));
  MUXF8 \sbox_inferred__0/block_w2_reg_reg[9]_i_6 
       (.I0(\sbox_inferred__0/block_w2_reg_reg[9]_i_11_n_0 ),
        .I1(\sbox_inferred__0/block_w2_reg_reg[9]_i_12_n_0 ),
        .O(new_sboxw[9]),
        .S(\block_w3_reg[31]_i_3 [3]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[16]_i_10 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[16]_i_5_2 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[16]_i_5_3 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[16]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF8 \sbox_inferred__1/block_w2_reg_reg[16]_i_5 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[16]_i_9_n_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[16]_i_10_n_0 ),
        .O(new_sboxw[16]),
        .S(\block_w3_reg[31]_i_3 [5]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[16]_i_9 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[16]_i_5_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[16]_i_5_1 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[16]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[17]_i_10 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[17]_i_5_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[17]_i_5_1 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[17]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[17]_i_11 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[17]_i_5_2 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[17]_i_5_3 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[17]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF8 \sbox_inferred__1/block_w2_reg_reg[17]_i_5 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[17]_i_10_n_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[17]_i_11_n_0 ),
        .O(new_sboxw[17]),
        .S(\block_w3_reg[31]_i_3 [5]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[18]_i_10 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[18]_i_5_2 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[18]_i_5_3 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[18]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF8 \sbox_inferred__1/block_w2_reg_reg[18]_i_5 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[18]_i_9_n_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[18]_i_10_n_0 ),
        .O(new_sboxw[18]),
        .S(\block_w3_reg[31]_i_3 [5]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[18]_i_9 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[18]_i_5_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[18]_i_5_1 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[18]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[19]_i_10 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[19]_i_5_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[19]_i_5_1 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[19]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[19]_i_11 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[19]_i_5_2 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[19]_i_5_3 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[19]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF8 \sbox_inferred__1/block_w2_reg_reg[19]_i_5 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[19]_i_10_n_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[19]_i_11_n_0 ),
        .O(new_sboxw[19]),
        .S(\block_w3_reg[31]_i_3 [5]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[20]_i_11 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[20]_i_6_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[20]_i_6_1 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[20]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[20]_i_12 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[20]_i_6_2 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[20]_i_6_3 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[20]_i_12_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF8 \sbox_inferred__1/block_w2_reg_reg[20]_i_6 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[20]_i_11_n_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[20]_i_12_n_0 ),
        .O(new_sboxw[20]),
        .S(\block_w3_reg[31]_i_3 [5]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[21]_i_10 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[21]_i_5_2 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[21]_i_5_3 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[21]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF8 \sbox_inferred__1/block_w2_reg_reg[21]_i_5 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[21]_i_9_n_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[21]_i_10_n_0 ),
        .O(new_sboxw[21]),
        .S(\block_w3_reg[31]_i_3 [5]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[21]_i_9 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[21]_i_5_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[21]_i_5_1 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[21]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[22]_i_10 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[22]_i_5_2 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[22]_i_5_3 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[22]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF8 \sbox_inferred__1/block_w2_reg_reg[22]_i_5 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[22]_i_9_n_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[22]_i_10_n_0 ),
        .O(new_sboxw[22]),
        .S(\block_w3_reg[31]_i_3 [5]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[22]_i_9 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[22]_i_5_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[22]_i_5_1 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[22]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[23]_i_10 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[23]_i_5_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[23]_i_5_1 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[23]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF7 \sbox_inferred__1/block_w2_reg_reg[23]_i_11 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[23]_i_5_2 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[23]_i_5_3 ),
        .O(\sbox_inferred__1/block_w2_reg_reg[23]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [4]));
  MUXF8 \sbox_inferred__1/block_w2_reg_reg[23]_i_5 
       (.I0(\sbox_inferred__1/block_w2_reg_reg[23]_i_10_n_0 ),
        .I1(\sbox_inferred__1/block_w2_reg_reg[23]_i_11_n_0 ),
        .O(new_sboxw[23]),
        .S(\block_w3_reg[31]_i_3 [5]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[24]_i_10 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[24]_i_5_2 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[24]_i_5_3 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[24]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF8 \sbox_inferred__2/block_w2_reg_reg[24]_i_5 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[24]_i_9_n_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[24]_i_10_n_0 ),
        .O(new_sboxw[24]),
        .S(\block_w3_reg[31]_i_3 [7]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[24]_i_9 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[24]_i_5_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[24]_i_5_1 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[24]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[25]_i_11 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[25]_i_6_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[25]_i_6_1 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[25]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[25]_i_12 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[25]_i_6_2 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[25]_i_6_3 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[25]_i_12_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF8 \sbox_inferred__2/block_w2_reg_reg[25]_i_6 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[25]_i_11_n_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[25]_i_12_n_0 ),
        .O(new_sboxw[25]),
        .S(\block_w3_reg[31]_i_3 [7]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[26]_i_10 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[26]_i_5_2 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[26]_i_5_3 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[26]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF8 \sbox_inferred__2/block_w2_reg_reg[26]_i_5 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[26]_i_9_n_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[26]_i_10_n_0 ),
        .O(new_sboxw[26]),
        .S(\block_w3_reg[31]_i_3 [7]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[26]_i_9 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[26]_i_5_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[26]_i_5_1 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[26]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[27]_i_12 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[27]_i_5_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[27]_i_5_1 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[27]_i_12_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[27]_i_13 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[27]_i_5_2 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[27]_i_5_3 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[27]_i_13_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF8 \sbox_inferred__2/block_w2_reg_reg[27]_i_5 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[27]_i_12_n_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[27]_i_13_n_0 ),
        .O(new_sboxw[27]),
        .S(\block_w3_reg[31]_i_3 [7]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[28]_i_11 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[28]_i_5_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[28]_i_5_1 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[28]_i_11_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[28]_i_12 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[28]_i_5_2 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[28]_i_5_3 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[28]_i_12_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF8 \sbox_inferred__2/block_w2_reg_reg[28]_i_5 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[28]_i_11_n_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[28]_i_12_n_0 ),
        .O(new_sboxw[28]),
        .S(\block_w3_reg[31]_i_3 [7]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[29]_i_10 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[29]_i_5_2 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[29]_i_5_3 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[29]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF8 \sbox_inferred__2/block_w2_reg_reg[29]_i_5 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[29]_i_9_n_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[29]_i_10_n_0 ),
        .O(new_sboxw[29]),
        .S(\block_w3_reg[31]_i_3 [7]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[29]_i_9 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[29]_i_5_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[29]_i_5_1 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[29]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[30]_i_10 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[30]_i_5_2 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[30]_i_5_3 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[30]_i_10_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF8 \sbox_inferred__2/block_w2_reg_reg[30]_i_5 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[30]_i_9_n_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[30]_i_10_n_0 ),
        .O(new_sboxw[30]),
        .S(\block_w3_reg[31]_i_3 [7]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[30]_i_9 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[30]_i_5_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[30]_i_5_1 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[30]_i_9_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF8 \sbox_inferred__2/block_w2_reg_reg[31]_i_10 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[31]_i_17_n_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[31]_i_18_n_0 ),
        .O(new_sboxw[31]),
        .S(\block_w3_reg[31]_i_3 [7]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[31]_i_17 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[31]_i_10_0 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[31]_i_10_1 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[31]_i_17_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
  MUXF7 \sbox_inferred__2/block_w2_reg_reg[31]_i_18 
       (.I0(\sbox_inferred__2/block_w2_reg_reg[31]_i_10_2 ),
        .I1(\sbox_inferred__2/block_w2_reg_reg[31]_i_10_3 ),
        .O(\sbox_inferred__2/block_w2_reg_reg[31]_i_18_n_0 ),
        .S(\block_w3_reg[31]_i_3 [6]));
endmodule
`ifndef GLBL
`define GLBL
`timescale  1 ps / 1 ps

module glbl ();

    parameter ROC_WIDTH = 100000;
    parameter TOC_WIDTH = 0;

//--------   STARTUP Globals --------------
    wire GSR;
    wire GTS;
    wire GWE;
    wire PRLD;
    tri1 p_up_tmp;
    tri (weak1, strong0) PLL_LOCKG = p_up_tmp;

    wire PROGB_GLBL;
    wire CCLKO_GLBL;
    wire FCSBO_GLBL;
    wire [3:0] DO_GLBL;
    wire [3:0] DI_GLBL;
   
    reg GSR_int;
    reg GTS_int;
    reg PRLD_int;

//--------   JTAG Globals --------------
    wire JTAG_TDO_GLBL;
    wire JTAG_TCK_GLBL;
    wire JTAG_TDI_GLBL;
    wire JTAG_TMS_GLBL;
    wire JTAG_TRST_GLBL;

    reg JTAG_CAPTURE_GLBL;
    reg JTAG_RESET_GLBL;
    reg JTAG_SHIFT_GLBL;
    reg JTAG_UPDATE_GLBL;
    reg JTAG_RUNTEST_GLBL;

    reg JTAG_SEL1_GLBL = 0;
    reg JTAG_SEL2_GLBL = 0 ;
    reg JTAG_SEL3_GLBL = 0;
    reg JTAG_SEL4_GLBL = 0;

    reg JTAG_USER_TDO1_GLBL = 1'bz;
    reg JTAG_USER_TDO2_GLBL = 1'bz;
    reg JTAG_USER_TDO3_GLBL = 1'bz;
    reg JTAG_USER_TDO4_GLBL = 1'bz;

    assign (strong1, weak0) GSR = GSR_int;
    assign (strong1, weak0) GTS = GTS_int;
    assign (weak1, weak0) PRLD = PRLD_int;

    initial begin
	GSR_int = 1'b1;
	PRLD_int = 1'b1;
	#(ROC_WIDTH)
	GSR_int = 1'b0;
	PRLD_int = 1'b0;
    end

    initial begin
	GTS_int = 1'b1;
	#(TOC_WIDTH)
	GTS_int = 1'b0;
    end

endmodule
`endif
