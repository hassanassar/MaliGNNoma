`timescale 1 ps / 1 ps
`define XIL_TIMING

module RAM64M8_UNIQ_BASE_
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39684
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39685
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39686
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39687
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39688
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39689
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39690
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39691
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39692
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39693
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39694
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39695
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39696
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39697
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39698
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39699
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39700
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39701
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39702
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39703
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39704
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39705
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39706
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39707
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39708
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39709
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39710
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39711
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39712
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39713
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39714
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39715
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39716
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39717
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39718
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39719
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39720
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39721
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39722
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39723
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39724
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39725
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39726
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39727
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39728
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39729
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39730
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39731
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39732
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39733
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39734
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39735
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39736
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39737
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39738
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39739
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39740
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39741
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39742
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39743
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39744
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39745
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39746
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39747
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39748
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39749
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39750
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39751
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39752
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39753
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39754
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39755
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39756
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39757
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39758
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39759
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39760
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39761
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39762
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39763
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39764
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39765
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39766
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39767
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39768
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39769
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39770
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39771
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39772
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39773
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39774
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39775
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39776
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39777
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39778
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39779
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39780
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39781
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39782
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39783
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39784
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39785
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39786
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39787
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39788
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39789
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39790
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39791
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39792
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39793
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39794
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39795
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39796
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39797
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39798
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39799
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39800
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39801
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39802
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39803
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39804
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39805
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39806
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39807
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39808
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39809
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39810
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39811
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39812
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39813
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39814
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39815
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39816
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39817
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39818
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39819
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39820
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39821
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39822
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39823
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39824
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39825
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39826
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39827
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39828
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39829
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39830
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39831
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39832
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39833
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39834
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39835
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39836
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39837
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39838
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39839
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39840
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39841
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39842
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39843
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39844
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39845
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39846
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39847
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39848
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39849
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39850
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39851
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39852
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39853
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39854
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39855
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39856
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39857
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39858
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39859
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39860
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39861
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39862
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39863
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39864
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39865
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39866
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39867
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39868
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39869
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39870
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39871
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39872
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39873
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39874
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39875
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39876
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39877
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39878
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39879
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39880
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39881
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39882
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39883
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39884
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39885
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39886
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39887
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39888
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39889
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39890
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39891
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39892
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39893
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39894
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39895
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39896
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39897
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39898
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39899
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39900
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39901
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39902
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39903
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39904
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39905
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39906
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39907
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39908
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39909
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39910
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39911
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39912
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39913
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39914
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39915
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39916
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39917
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39918
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39919
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39920
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39921
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39922
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39923
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39924
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39925
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39926
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39927
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39928
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39929
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39930
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39931
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

module RAM64M8_HD39932
   (DOA,
    DOB,
    DOC,
    DOD,
    DOE,
    DOF,
    DOG,
    DOH,
    ADDRA,
    ADDRB,
    ADDRC,
    ADDRD,
    ADDRE,
    ADDRF,
    ADDRG,
    ADDRH,
    DIA,
    DIB,
    DIC,
    DID,
    DIE,
    DIF,
    DIG,
    DIH,
    WCLK,
    WE);
  output DOA;
  output DOB;
  output DOC;
  output DOD;
  output DOE;
  output DOF;
  output DOG;
  output DOH;
  input [5:0]ADDRA;
  input [5:0]ADDRB;
  input [5:0]ADDRC;
  input [5:0]ADDRD;
  input [5:0]ADDRE;
  input [5:0]ADDRF;
  input [5:0]ADDRG;
  input [5:0]ADDRH;
  input DIA;
  input DIB;
  input DIC;
  input DID;
  input DIE;
  input DIF;
  input DIG;
  input DIH;
  input WCLK;
  input WE;

  wire ADDRA0;
  wire ADDRA1;
  wire ADDRA2;
  wire ADDRA3;
  wire ADDRA4;
  wire ADDRA5;
  wire ADDRB0;
  wire ADDRB1;
  wire ADDRB2;
  wire ADDRB3;
  wire ADDRB4;
  wire ADDRB5;
  wire ADDRC0;
  wire ADDRC1;
  wire ADDRC2;
  wire ADDRC3;
  wire ADDRC4;
  wire ADDRC5;
  wire ADDRD0;
  wire ADDRD1;
  wire ADDRD2;
  wire ADDRD3;
  wire ADDRD4;
  wire ADDRD5;
  wire ADDRE0;
  wire ADDRE1;
  wire ADDRE2;
  wire ADDRE3;
  wire ADDRE4;
  wire ADDRE5;
  wire ADDRF0;
  wire ADDRF1;
  wire ADDRF2;
  wire ADDRF3;
  wire ADDRF4;
  wire ADDRF5;
  wire ADDRG0;
  wire ADDRG1;
  wire ADDRG2;
  wire ADDRG3;
  wire ADDRG4;
  wire ADDRG5;
  wire ADDRH0;
  wire ADDRH1;
  wire ADDRH2;
  wire ADDRH3;
  wire ADDRH4;
  wire ADDRH5;
  wire DIA;
  wire DIB;
  wire DIC;
  wire DID;
  wire DIE;
  wire DIF;
  wire DIG;
  wire DIH;
  wire DOA;
  wire DOB;
  wire DOC;
  wire DOD;
  wire DOE;
  wire DOF;
  wire DOG;
  wire DOH;
  wire WCLK;
  wire WE;
  wire NLW_RAMA_WADR6_UNCONNECTED;
  wire NLW_RAMA_WADR7_UNCONNECTED;
  wire NLW_RAMB_WADR6_UNCONNECTED;
  wire NLW_RAMB_WADR7_UNCONNECTED;
  wire NLW_RAMC_WADR6_UNCONNECTED;
  wire NLW_RAMC_WADR7_UNCONNECTED;
  wire NLW_RAMD_WADR6_UNCONNECTED;
  wire NLW_RAMD_WADR7_UNCONNECTED;
  wire NLW_RAME_WADR6_UNCONNECTED;
  wire NLW_RAME_WADR7_UNCONNECTED;
  wire NLW_RAMF_WADR6_UNCONNECTED;
  wire NLW_RAMF_WADR7_UNCONNECTED;
  wire NLW_RAMG_WADR6_UNCONNECTED;
  wire NLW_RAMG_WADR7_UNCONNECTED;
  wire NLW_RAMH_WADR6_UNCONNECTED;
  wire NLW_RAMH_WADR7_UNCONNECTED;

  assign ADDRA0 = ADDRA[0];
  assign ADDRA1 = ADDRA[1];
  assign ADDRA2 = ADDRA[2];
  assign ADDRA3 = ADDRA[3];
  assign ADDRA4 = ADDRA[4];
  assign ADDRA5 = ADDRA[5];
  assign ADDRB0 = ADDRB[0];
  assign ADDRB1 = ADDRB[1];
  assign ADDRB2 = ADDRB[2];
  assign ADDRB3 = ADDRB[3];
  assign ADDRB4 = ADDRB[4];
  assign ADDRB5 = ADDRB[5];
  assign ADDRC0 = ADDRC[0];
  assign ADDRC1 = ADDRC[1];
  assign ADDRC2 = ADDRC[2];
  assign ADDRC3 = ADDRC[3];
  assign ADDRC4 = ADDRC[4];
  assign ADDRC5 = ADDRC[5];
  assign ADDRD0 = ADDRD[0];
  assign ADDRD1 = ADDRD[1];
  assign ADDRD2 = ADDRD[2];
  assign ADDRD3 = ADDRD[3];
  assign ADDRD4 = ADDRD[4];
  assign ADDRD5 = ADDRD[5];
  assign ADDRE0 = ADDRE[0];
  assign ADDRE1 = ADDRE[1];
  assign ADDRE2 = ADDRE[2];
  assign ADDRE3 = ADDRE[3];
  assign ADDRE4 = ADDRE[4];
  assign ADDRE5 = ADDRE[5];
  assign ADDRF0 = ADDRF[0];
  assign ADDRF1 = ADDRF[1];
  assign ADDRF2 = ADDRF[2];
  assign ADDRF3 = ADDRF[3];
  assign ADDRF4 = ADDRF[4];
  assign ADDRF5 = ADDRF[5];
  assign ADDRG0 = ADDRG[0];
  assign ADDRG1 = ADDRG[1];
  assign ADDRG2 = ADDRG[2];
  assign ADDRG3 = ADDRG[3];
  assign ADDRG4 = ADDRG[4];
  assign ADDRG5 = ADDRG[5];
  assign ADDRH0 = ADDRH[0];
  assign ADDRH1 = ADDRH[1];
  assign ADDRH2 = ADDRH[2];
  assign ADDRH3 = ADDRH[3];
  assign ADDRH4 = ADDRH[4];
  assign ADDRH5 = ADDRH[5];
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMA
       (.CLK(WCLK),
        .I(DIA),
        .O(DOA),
        .RADR0(ADDRA0),
        .RADR1(ADDRA1),
        .RADR2(ADDRA2),
        .RADR3(ADDRA3),
        .RADR4(ADDRA4),
        .RADR5(ADDRA5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMA_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMA_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMB
       (.CLK(WCLK),
        .I(DIB),
        .O(DOB),
        .RADR0(ADDRB0),
        .RADR1(ADDRB1),
        .RADR2(ADDRB2),
        .RADR3(ADDRB3),
        .RADR4(ADDRB4),
        .RADR5(ADDRB5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMB_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMB_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMC
       (.CLK(WCLK),
        .I(DIC),
        .O(DOC),
        .RADR0(ADDRC0),
        .RADR1(ADDRC1),
        .RADR2(ADDRC2),
        .RADR3(ADDRC3),
        .RADR4(ADDRC4),
        .RADR5(ADDRC5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMC_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMC_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMD
       (.CLK(WCLK),
        .I(DID),
        .O(DOD),
        .RADR0(ADDRD0),
        .RADR1(ADDRD1),
        .RADR2(ADDRD2),
        .RADR3(ADDRD3),
        .RADR4(ADDRD4),
        .RADR5(ADDRD5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMD_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMD_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAME
       (.CLK(WCLK),
        .I(DIE),
        .O(DOE),
        .RADR0(ADDRE0),
        .RADR1(ADDRE1),
        .RADR2(ADDRE2),
        .RADR3(ADDRE3),
        .RADR4(ADDRE4),
        .RADR5(ADDRE5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAME_WADR6_UNCONNECTED),
        .WADR7(NLW_RAME_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMF
       (.CLK(WCLK),
        .I(DIF),
        .O(DOF),
        .RADR0(ADDRF0),
        .RADR1(ADDRF1),
        .RADR2(ADDRF2),
        .RADR3(ADDRF3),
        .RADR4(ADDRF4),
        .RADR5(ADDRF5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMF_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMF_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMG
       (.CLK(WCLK),
        .I(DIG),
        .O(DOG),
        .RADR0(ADDRG0),
        .RADR1(ADDRG1),
        .RADR2(ADDRG2),
        .RADR3(ADDRG3),
        .RADR4(ADDRG4),
        .RADR5(ADDRG5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMG_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMG_WADR7_UNCONNECTED),
        .WE(WE));
  RAMD64E #(
    .INIT(64'h0000000000000000),
    .IS_CLK_INVERTED(1'b0),
    .RAM_ADDRESS_MASK(2'b11),
    .RAM_ADDRESS_SPACE(2'b11)) 
    RAMH
       (.CLK(WCLK),
        .I(DIH),
        .O(DOH),
        .RADR0(ADDRH0),
        .RADR1(ADDRH1),
        .RADR2(ADDRH2),
        .RADR3(ADDRH3),
        .RADR4(ADDRH4),
        .RADR5(ADDRH5),
        .WADR0(ADDRH0),
        .WADR1(ADDRH1),
        .WADR2(ADDRH2),
        .WADR3(ADDRH3),
        .WADR4(ADDRH4),
        .WADR5(ADDRH5),
        .WADR6(NLW_RAMH_WADR6_UNCONNECTED),
        .WADR7(NLW_RAMH_WADR7_UNCONNECTED),
        .WE(WE));
endmodule

(* dont_touch = "true" *) 
(* NotValidForBitStream *)
module switch_elements
   (enable_i,
    clk_i,
    rst_i,
    info_o);
  input [31:0]enable_i;
  input clk_i;
  input rst_i;
  output [31:0]info_o;

  wire clk_i;
  wire [31:0]enable_i;
  (* DONT_TOUCH *) wire [31:0]info_s;
  wire \info_s[0]_i_1_n_0 ;
  wire \info_s[10]_i_1_n_0 ;
  wire \info_s[11]_i_1_n_0 ;
  wire \info_s[12]_i_1_n_0 ;
  wire \info_s[13]_i_1_n_0 ;
  wire \info_s[14]_i_1_n_0 ;
  wire \info_s[15]_i_1_n_0 ;
  wire \info_s[16]_i_1_n_0 ;
  wire \info_s[17]_i_1_n_0 ;
  wire \info_s[18]_i_1_n_0 ;
  wire \info_s[19]_i_1_n_0 ;
  wire \info_s[1]_i_1_n_0 ;
  wire \info_s[20]_i_1_n_0 ;
  wire \info_s[21]_i_1_n_0 ;
  wire \info_s[22]_i_1_n_0 ;
  wire \info_s[23]_i_1_n_0 ;
  wire \info_s[24]_i_1_n_0 ;
  wire \info_s[25]_i_1_n_0 ;
  wire \info_s[26]_i_1_n_0 ;
  wire \info_s[27]_i_1_n_0 ;
  wire \info_s[28]_i_1_n_0 ;
  wire \info_s[29]_i_1_n_0 ;
  wire \info_s[2]_i_1_n_0 ;
  wire \info_s[30]_i_1_n_0 ;
  wire \info_s[31]_i_1_n_0 ;
  wire \info_s[3]_i_1_n_0 ;
  wire \info_s[4]_i_1_n_0 ;
  wire \info_s[5]_i_1_n_0 ;
  wire \info_s[6]_i_1_n_0 ;
  wire \info_s[7]_i_1_n_0 ;
  wire \info_s[8]_i_1_n_0 ;
  wire \info_s[9]_i_1_n_0 ;
  (* DONT_TOUCH *) wire [31:0]\info_v[0] ;
  wire rst_i;

  assign info_o[31:0] = info_s;
  (* DONT_TOUCH *) 
  switch_elements_switch_elements3 \activity_blocks[0].switch 
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .info_o(\info_v[0] ),
        .rst_i(rst_i));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[0]_i_1 
       (.I0(\info_v[0] [0]),
        .I1(info_s[0]),
        .O(\info_s[0]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[10]_i_1 
       (.I0(\info_v[0] [10]),
        .I1(info_s[10]),
        .O(\info_s[10]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[11]_i_1 
       (.I0(\info_v[0] [11]),
        .I1(info_s[11]),
        .O(\info_s[11]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[12]_i_1 
       (.I0(\info_v[0] [12]),
        .I1(info_s[12]),
        .O(\info_s[12]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[13]_i_1 
       (.I0(\info_v[0] [13]),
        .I1(info_s[13]),
        .O(\info_s[13]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[14]_i_1 
       (.I0(\info_v[0] [14]),
        .I1(info_s[14]),
        .O(\info_s[14]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[15]_i_1 
       (.I0(\info_v[0] [15]),
        .I1(info_s[15]),
        .O(\info_s[15]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[16]_i_1 
       (.I0(\info_v[0] [16]),
        .I1(info_s[16]),
        .O(\info_s[16]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[17]_i_1 
       (.I0(\info_v[0] [17]),
        .I1(info_s[17]),
        .O(\info_s[17]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[18]_i_1 
       (.I0(\info_v[0] [18]),
        .I1(info_s[18]),
        .O(\info_s[18]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[19]_i_1 
       (.I0(\info_v[0] [19]),
        .I1(info_s[19]),
        .O(\info_s[19]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[1]_i_1 
       (.I0(\info_v[0] [1]),
        .I1(info_s[1]),
        .O(\info_s[1]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[20]_i_1 
       (.I0(\info_v[0] [20]),
        .I1(info_s[20]),
        .O(\info_s[20]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[21]_i_1 
       (.I0(\info_v[0] [21]),
        .I1(info_s[21]),
        .O(\info_s[21]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[22]_i_1 
       (.I0(\info_v[0] [22]),
        .I1(info_s[22]),
        .O(\info_s[22]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[23]_i_1 
       (.I0(\info_v[0] [23]),
        .I1(info_s[23]),
        .O(\info_s[23]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[24]_i_1 
       (.I0(\info_v[0] [24]),
        .I1(info_s[24]),
        .O(\info_s[24]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[25]_i_1 
       (.I0(\info_v[0] [25]),
        .I1(info_s[25]),
        .O(\info_s[25]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[26]_i_1 
       (.I0(\info_v[0] [26]),
        .I1(info_s[26]),
        .O(\info_s[26]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[27]_i_1 
       (.I0(\info_v[0] [27]),
        .I1(info_s[27]),
        .O(\info_s[27]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[28]_i_1 
       (.I0(\info_v[0] [28]),
        .I1(info_s[28]),
        .O(\info_s[28]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[29]_i_1 
       (.I0(\info_v[0] [29]),
        .I1(info_s[29]),
        .O(\info_s[29]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[2]_i_1 
       (.I0(\info_v[0] [2]),
        .I1(info_s[2]),
        .O(\info_s[2]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[30]_i_1 
       (.I0(\info_v[0] [30]),
        .I1(info_s[30]),
        .O(\info_s[30]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[31]_i_1 
       (.I0(\info_v[0] [31]),
        .I1(info_s[31]),
        .O(\info_s[31]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[3]_i_1 
       (.I0(\info_v[0] [3]),
        .I1(info_s[3]),
        .O(\info_s[3]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[4]_i_1 
       (.I0(\info_v[0] [4]),
        .I1(info_s[4]),
        .O(\info_s[4]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[5]_i_1 
       (.I0(\info_v[0] [5]),
        .I1(info_s[5]),
        .O(\info_s[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[6]_i_1 
       (.I0(\info_v[0] [6]),
        .I1(info_s[6]),
        .O(\info_s[6]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[7]_i_1 
       (.I0(\info_v[0] [7]),
        .I1(info_s[7]),
        .O(\info_s[7]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[8]_i_1 
       (.I0(\info_v[0] [8]),
        .I1(info_s[8]),
        .O(\info_s[8]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \info_s[9]_i_1 
       (.I0(\info_v[0] [9]),
        .I1(info_s[9]),
        .O(\info_s[9]_i_1_n_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[0]_i_1_n_0 ),
        .Q(info_s[0]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[10]_i_1_n_0 ),
        .Q(info_s[10]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[11]_i_1_n_0 ),
        .Q(info_s[11]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[12]_i_1_n_0 ),
        .Q(info_s[12]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[13]_i_1_n_0 ),
        .Q(info_s[13]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[14]_i_1_n_0 ),
        .Q(info_s[14]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[15]_i_1_n_0 ),
        .Q(info_s[15]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[16]_i_1_n_0 ),
        .Q(info_s[16]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[17]_i_1_n_0 ),
        .Q(info_s[17]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[18]_i_1_n_0 ),
        .Q(info_s[18]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[19]_i_1_n_0 ),
        .Q(info_s[19]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[1]_i_1_n_0 ),
        .Q(info_s[1]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[20]_i_1_n_0 ),
        .Q(info_s[20]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[21]_i_1_n_0 ),
        .Q(info_s[21]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[22]_i_1_n_0 ),
        .Q(info_s[22]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[23]_i_1_n_0 ),
        .Q(info_s[23]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[24]_i_1_n_0 ),
        .Q(info_s[24]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[25]_i_1_n_0 ),
        .Q(info_s[25]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[26]_i_1_n_0 ),
        .Q(info_s[26]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[27]_i_1_n_0 ),
        .Q(info_s[27]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[28]_i_1_n_0 ),
        .Q(info_s[28]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[29]_i_1_n_0 ),
        .Q(info_s[29]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[2]_i_1_n_0 ),
        .Q(info_s[2]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[30]_i_1_n_0 ),
        .Q(info_s[30]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[31]_i_1_n_0 ),
        .Q(info_s[31]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[3]_i_1_n_0 ),
        .Q(info_s[3]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[4]_i_1_n_0 ),
        .Q(info_s[4]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[5]_i_1_n_0 ),
        .Q(info_s[5]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[6]_i_1_n_0 ),
        .Q(info_s[6]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[7]_i_1_n_0 ),
        .Q(info_s[7]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[8]_i_1_n_0 ),
        .Q(info_s[8]),
        .R(1'b0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \info_s_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\info_s[9]_i_1_n_0 ),
        .Q(info_s[9]),
        .R(1'b0));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8" *) 
module switch_elements_cf_fft_512_8
   (p_6_out,
    rst_i,
    enable_i,
    clk_i,
    enable_s,
    DOUTADOUT,
    n14__56_carry);
  output [31:0]p_6_out;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [31:0]enable_s;
  input [15:0]DOUTADOUT;
  input [15:0]n14__56_carry;

  wire [15:0]DOUTADOUT;
  wire clk_i;
  wire [0:0]enable_i;
  wire [31:0]enable_s;
  wire [15:0]n14__56_carry;
  wire [31:0]p_6_out;
  wire rst_i;

  switch_elements_cf_fft_512_8_1 s1
       (.DOUTADOUT(DOUTADOUT),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .enable_s(enable_s),
        .n14__56_carry(n14__56_carry),
        .p_6_out(p_6_out),
        .rst_i(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_1" *) 
module switch_elements_cf_fft_512_8_1
   (p_6_out,
    rst_i,
    enable_i,
    clk_i,
    enable_s,
    DOUTADOUT,
    n14__56_carry);
  output [31:0]p_6_out;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [31:0]enable_s;
  input [15:0]DOUTADOUT;
  input [15:0]n14__56_carry;

  wire [7:0]A;
  wire [15:0]DOUTADOUT;
  wire clk_i;
  wire [0:0]enable_i;
  wire [31:0]enable_s;
  wire [31:0]inf4_s;
  wire [15:0]n110_out;
  wire [15:0]n14__56_carry;
  wire [31:0]p_6_out;
  wire rst_i;
  wire [15:0]s1_2;
  wire [15:0]s1_3;
  wire s1_n_0;
  wire s3_n_16;
  wire s3_n_17;
  wire s3_n_18;
  wire s3_n_19;
  wire s3_n_20;
  wire s3_n_21;
  wire s3_n_22;
  wire s3_n_23;

  switch_elements_cf_fft_512_8_21 s1
       (.D(s1_2),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .\n1_reg[15] (n110_out),
        .n22(A),
        .\n4_reg[7] ({s3_n_16,s3_n_17,s3_n_18,s3_n_19,s3_n_20,s3_n_21,s3_n_22,s3_n_23}),
        .\n9_reg[0] (s1_n_0),
        .rst_i(rst_i),
        .s1_3(s1_3));
  switch_elements_cf_fft_512_8_5 s2
       (.DOUTADOUT(DOUTADOUT),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .enable_s(enable_s),
        .i2(s1_2),
        .i3(s1_3),
        .inf4_s(inf4_s),
        .n14__56_carry(n14__56_carry),
        .p_6_out(p_6_out),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_2 s3
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i2({inf4_s[15:0],inf4_s[31:16]}),
        .n22(s1_n_0),
        .\n5_reg[0] (n110_out),
        .\n5_reg[0]_0 ({s3_n_16,s3_n_17,s3_n_18,s3_n_19,s3_n_20,s3_n_21,s3_n_22,s3_n_23}),
        .\n5_reg[0]_1 (A),
        .rst_i(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_10" *) 
module switch_elements_cf_fft_512_8_10
   (i1,
    rst_i,
    enable_i,
    clk_i,
    s7_3,
    D);
  output [29:0]i1;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]s7_3;
  input [15:0]D;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [7:0]n10;
  wire [7:0]n15;
  wire \n16[3]_i_10_n_0 ;
  wire \n16[3]_i_11_n_0 ;
  wire \n16[3]_i_12_n_0 ;
  wire \n16[3]_i_13_n_0 ;
  wire \n16[3]_i_14__0_n_0 ;
  wire \n16[3]_i_15__0_n_0 ;
  wire \n16[3]_i_16_n_0 ;
  wire \n16[3]_i_18_n_0 ;
  wire \n16[3]_i_19_n_0 ;
  wire \n16[3]_i_20_n_0 ;
  wire \n16[3]_i_21_n_0 ;
  wire \n16[3]_i_22_n_0 ;
  wire \n16[3]_i_23__0_n_0 ;
  wire \n16[3]_i_24__0_n_0 ;
  wire \n16[3]_i_25__0_n_0 ;
  wire \n16[3]_i_26__0_n_0 ;
  wire \n16[3]_i_27_n_0 ;
  wire \n16[3]_i_28__0_n_0 ;
  wire \n16[3]_i_2_n_0 ;
  wire \n16[3]_i_3_n_0 ;
  wire \n16[3]_i_4_n_0 ;
  wire \n16[3]_i_5_n_0 ;
  wire \n16[3]_i_6__0_n_0 ;
  wire \n16[3]_i_7_n_0 ;
  wire \n16[3]_i_8_n_0 ;
  wire \n16[3]_i_9_n_0 ;
  wire \n16[7]_i_13__0_n_0 ;
  wire \n16[7]_i_14_n_0 ;
  wire \n16[7]_i_15__0_n_0 ;
  wire \n16[7]_i_16__0_n_0 ;
  wire \n16[7]_i_17_n_0 ;
  wire \n16[7]_i_18_n_0 ;
  wire \n16[7]_i_19__0_n_0 ;
  wire \n16[7]_i_20__0_n_0 ;
  wire \n16[7]_i_21__0_n_0 ;
  wire \n16[7]_i_22_n_0 ;
  wire \n16[7]_i_23__0_n_0 ;
  wire \n16[7]_i_24_n_0 ;
  wire \n16[7]_i_25_n_0 ;
  wire \n16[7]_i_26_n_0 ;
  wire \n16[7]_i_27_n_0 ;
  wire \n16[7]_i_28_n_0 ;
  wire \n16[7]_i_29__0_n_0 ;
  wire \n16[7]_i_2_n_0 ;
  wire \n16[7]_i_30__0_n_0 ;
  wire \n16[7]_i_31__0_n_0 ;
  wire \n16[7]_i_32__0_n_0 ;
  wire \n16[7]_i_33_n_0 ;
  wire \n16[7]_i_34__0_n_0 ;
  wire \n16[7]_i_35__0_n_0 ;
  wire \n16[7]_i_36_n_0 ;
  wire \n16[7]_i_37__0_n_0 ;
  wire \n16[7]_i_38__0_n_0 ;
  wire \n16[7]_i_3_n_0 ;
  wire \n16[7]_i_4_n_0 ;
  wire \n16[7]_i_5__0_n_0 ;
  wire \n16[7]_i_6__0_n_0 ;
  wire \n16[7]_i_7__0_n_0 ;
  wire \n16[7]_i_8_n_0 ;
  wire \n16_reg[3]_i_17_n_0 ;
  wire \n16_reg[3]_i_17_n_1 ;
  wire \n16_reg[3]_i_17_n_10 ;
  wire \n16_reg[3]_i_17_n_11 ;
  wire \n16_reg[3]_i_17_n_12 ;
  wire \n16_reg[3]_i_17_n_15 ;
  wire \n16_reg[3]_i_17_n_2 ;
  wire \n16_reg[3]_i_17_n_3 ;
  wire \n16_reg[3]_i_17_n_4 ;
  wire \n16_reg[3]_i_17_n_5 ;
  wire \n16_reg[3]_i_17_n_6 ;
  wire \n16_reg[3]_i_17_n_7 ;
  wire \n16_reg[3]_i_17_n_8 ;
  wire \n16_reg[3]_i_17_n_9 ;
  wire \n16_reg[3]_i_1_n_0 ;
  wire \n16_reg[3]_i_1_n_1 ;
  wire \n16_reg[3]_i_1_n_2 ;
  wire \n16_reg[3]_i_1_n_3 ;
  wire \n16_reg[3]_i_1_n_4 ;
  wire \n16_reg[3]_i_1_n_5 ;
  wire \n16_reg[3]_i_1_n_6 ;
  wire \n16_reg[3]_i_1_n_7 ;
  wire \n16_reg[7]_i_10_n_1 ;
  wire \n16_reg[7]_i_10_n_10 ;
  wire \n16_reg[7]_i_10_n_11 ;
  wire \n16_reg[7]_i_10_n_12 ;
  wire \n16_reg[7]_i_10_n_13 ;
  wire \n16_reg[7]_i_10_n_14 ;
  wire \n16_reg[7]_i_10_n_15 ;
  wire \n16_reg[7]_i_10_n_2 ;
  wire \n16_reg[7]_i_10_n_3 ;
  wire \n16_reg[7]_i_10_n_4 ;
  wire \n16_reg[7]_i_10_n_5 ;
  wire \n16_reg[7]_i_10_n_6 ;
  wire \n16_reg[7]_i_10_n_7 ;
  wire \n16_reg[7]_i_10_n_8 ;
  wire \n16_reg[7]_i_10_n_9 ;
  wire \n16_reg[7]_i_11_n_0 ;
  wire \n16_reg[7]_i_11_n_1 ;
  wire \n16_reg[7]_i_11_n_10 ;
  wire \n16_reg[7]_i_11_n_11 ;
  wire \n16_reg[7]_i_11_n_12 ;
  wire \n16_reg[7]_i_11_n_13 ;
  wire \n16_reg[7]_i_11_n_14 ;
  wire \n16_reg[7]_i_11_n_2 ;
  wire \n16_reg[7]_i_11_n_3 ;
  wire \n16_reg[7]_i_11_n_4 ;
  wire \n16_reg[7]_i_11_n_5 ;
  wire \n16_reg[7]_i_11_n_6 ;
  wire \n16_reg[7]_i_11_n_7 ;
  wire \n16_reg[7]_i_11_n_8 ;
  wire \n16_reg[7]_i_11_n_9 ;
  wire \n16_reg[7]_i_12_n_14 ;
  wire \n16_reg[7]_i_12_n_15 ;
  wire \n16_reg[7]_i_12_n_5 ;
  wire \n16_reg[7]_i_12_n_7 ;
  wire \n16_reg[7]_i_1_n_5 ;
  wire \n16_reg[7]_i_1_n_6 ;
  wire \n16_reg[7]_i_1_n_7 ;
  wire \n16_reg[7]_i_9_n_14 ;
  wire \n16_reg[7]_i_9_n_15 ;
  wire \n16_reg[7]_i_9_n_5 ;
  wire \n16_reg[7]_i_9_n_7 ;
  wire \n16_reg_n_0_[0] ;
  wire \n16_reg_n_0_[1] ;
  wire \n16_reg_n_0_[2] ;
  wire \n16_reg_n_0_[3] ;
  wire \n16_reg_n_0_[4] ;
  wire \n16_reg_n_0_[5] ;
  wire \n16_reg_n_0_[6] ;
  wire \n16_reg_n_0_[7] ;
  wire \n1_reg_n_0_[0] ;
  wire \n1_reg_n_0_[1] ;
  wire \n1_reg_n_0_[2] ;
  wire \n1_reg_n_0_[3] ;
  wire \n1_reg_n_0_[4] ;
  wire \n1_reg_n_0_[5] ;
  wire \n1_reg_n_0_[6] ;
  wire \n1_reg_n_0_[7] ;
  wire [7:0]n2;
  wire [7:0]n202_out;
  wire [7:0]n21;
  wire \n21[7]_i_2__0_n_0 ;
  wire \n21[7]_i_3__0_n_0 ;
  wire \n21[7]_i_4__0_n_0 ;
  wire \n21[7]_i_5__0_n_0 ;
  wire \n21[7]_i_6__0_n_0 ;
  wire \n21[7]_i_7__0_n_0 ;
  wire \n21[7]_i_8__0_n_0 ;
  wire \n21[7]_i_9__0_n_0 ;
  wire \n21_reg[7]_i_1__0_n_1 ;
  wire \n21_reg[7]_i_1__0_n_2 ;
  wire \n21_reg[7]_i_1__0_n_3 ;
  wire \n21_reg[7]_i_1__0_n_4 ;
  wire \n21_reg[7]_i_1__0_n_5 ;
  wire \n21_reg[7]_i_1__0_n_6 ;
  wire \n21_reg[7]_i_1__0_n_7 ;
  wire n22__0_n_0;
  wire n22__1_n_0;
  wire n22__2_n_0;
  wire n22__3_n_0;
  wire n22__4_n_0;
  wire n22__5_n_0;
  wire n22__6_n_0;
  wire n22_n_0;
  wire [7:0]n26;
  wire [7:0]n27;
  wire \n27[3]_i_10_n_0 ;
  wire \n27[3]_i_11_n_0 ;
  wire \n27[3]_i_12_n_0 ;
  wire \n27[3]_i_13_n_0 ;
  wire \n27[3]_i_14__0_n_0 ;
  wire \n27[3]_i_15__0_n_0 ;
  wire \n27[3]_i_16_n_0 ;
  wire \n27[3]_i_18_n_0 ;
  wire \n27[3]_i_19_n_0 ;
  wire \n27[3]_i_20_n_0 ;
  wire \n27[3]_i_21_n_0 ;
  wire \n27[3]_i_22_n_0 ;
  wire \n27[3]_i_23__0_n_0 ;
  wire \n27[3]_i_24__0_n_0 ;
  wire \n27[3]_i_25__0_n_0 ;
  wire \n27[3]_i_26__0_n_0 ;
  wire \n27[3]_i_27_n_0 ;
  wire \n27[3]_i_28__0_n_0 ;
  wire \n27[3]_i_2_n_0 ;
  wire \n27[3]_i_3_n_0 ;
  wire \n27[3]_i_4_n_0 ;
  wire \n27[3]_i_5_n_0 ;
  wire \n27[3]_i_6__0_n_0 ;
  wire \n27[3]_i_7_n_0 ;
  wire \n27[3]_i_8_n_0 ;
  wire \n27[3]_i_9_n_0 ;
  wire \n27[7]_i_13__0_n_0 ;
  wire \n27[7]_i_14_n_0 ;
  wire \n27[7]_i_15__0_n_0 ;
  wire \n27[7]_i_16__0_n_0 ;
  wire \n27[7]_i_17_n_0 ;
  wire \n27[7]_i_18_n_0 ;
  wire \n27[7]_i_19__0_n_0 ;
  wire \n27[7]_i_20__0_n_0 ;
  wire \n27[7]_i_21__0_n_0 ;
  wire \n27[7]_i_22_n_0 ;
  wire \n27[7]_i_23__0_n_0 ;
  wire \n27[7]_i_24_n_0 ;
  wire \n27[7]_i_25_n_0 ;
  wire \n27[7]_i_26_n_0 ;
  wire \n27[7]_i_27_n_0 ;
  wire \n27[7]_i_28_n_0 ;
  wire \n27[7]_i_29__0_n_0 ;
  wire \n27[7]_i_2_n_0 ;
  wire \n27[7]_i_30__0_n_0 ;
  wire \n27[7]_i_31__0_n_0 ;
  wire \n27[7]_i_32__0_n_0 ;
  wire \n27[7]_i_33_n_0 ;
  wire \n27[7]_i_34__0_n_0 ;
  wire \n27[7]_i_35__0_n_0 ;
  wire \n27[7]_i_36_n_0 ;
  wire \n27[7]_i_37__0_n_0 ;
  wire \n27[7]_i_38__0_n_0 ;
  wire \n27[7]_i_3_n_0 ;
  wire \n27[7]_i_4_n_0 ;
  wire \n27[7]_i_5__0_n_0 ;
  wire \n27[7]_i_6__0_n_0 ;
  wire \n27[7]_i_7__0_n_0 ;
  wire \n27[7]_i_8_n_0 ;
  wire \n27_reg[3]_i_17_n_0 ;
  wire \n27_reg[3]_i_17_n_1 ;
  wire \n27_reg[3]_i_17_n_10 ;
  wire \n27_reg[3]_i_17_n_11 ;
  wire \n27_reg[3]_i_17_n_12 ;
  wire \n27_reg[3]_i_17_n_15 ;
  wire \n27_reg[3]_i_17_n_2 ;
  wire \n27_reg[3]_i_17_n_3 ;
  wire \n27_reg[3]_i_17_n_4 ;
  wire \n27_reg[3]_i_17_n_5 ;
  wire \n27_reg[3]_i_17_n_6 ;
  wire \n27_reg[3]_i_17_n_7 ;
  wire \n27_reg[3]_i_17_n_8 ;
  wire \n27_reg[3]_i_17_n_9 ;
  wire \n27_reg[3]_i_1_n_0 ;
  wire \n27_reg[3]_i_1_n_1 ;
  wire \n27_reg[3]_i_1_n_2 ;
  wire \n27_reg[3]_i_1_n_3 ;
  wire \n27_reg[3]_i_1_n_4 ;
  wire \n27_reg[3]_i_1_n_5 ;
  wire \n27_reg[3]_i_1_n_6 ;
  wire \n27_reg[3]_i_1_n_7 ;
  wire \n27_reg[7]_i_10_n_1 ;
  wire \n27_reg[7]_i_10_n_10 ;
  wire \n27_reg[7]_i_10_n_11 ;
  wire \n27_reg[7]_i_10_n_12 ;
  wire \n27_reg[7]_i_10_n_13 ;
  wire \n27_reg[7]_i_10_n_14 ;
  wire \n27_reg[7]_i_10_n_15 ;
  wire \n27_reg[7]_i_10_n_2 ;
  wire \n27_reg[7]_i_10_n_3 ;
  wire \n27_reg[7]_i_10_n_4 ;
  wire \n27_reg[7]_i_10_n_5 ;
  wire \n27_reg[7]_i_10_n_6 ;
  wire \n27_reg[7]_i_10_n_7 ;
  wire \n27_reg[7]_i_10_n_8 ;
  wire \n27_reg[7]_i_10_n_9 ;
  wire \n27_reg[7]_i_11_n_0 ;
  wire \n27_reg[7]_i_11_n_1 ;
  wire \n27_reg[7]_i_11_n_10 ;
  wire \n27_reg[7]_i_11_n_11 ;
  wire \n27_reg[7]_i_11_n_12 ;
  wire \n27_reg[7]_i_11_n_13 ;
  wire \n27_reg[7]_i_11_n_14 ;
  wire \n27_reg[7]_i_11_n_2 ;
  wire \n27_reg[7]_i_11_n_3 ;
  wire \n27_reg[7]_i_11_n_4 ;
  wire \n27_reg[7]_i_11_n_5 ;
  wire \n27_reg[7]_i_11_n_6 ;
  wire \n27_reg[7]_i_11_n_7 ;
  wire \n27_reg[7]_i_11_n_8 ;
  wire \n27_reg[7]_i_11_n_9 ;
  wire \n27_reg[7]_i_12_n_14 ;
  wire \n27_reg[7]_i_12_n_15 ;
  wire \n27_reg[7]_i_12_n_5 ;
  wire \n27_reg[7]_i_12_n_7 ;
  wire \n27_reg[7]_i_1_n_5 ;
  wire \n27_reg[7]_i_1_n_6 ;
  wire \n27_reg[7]_i_1_n_7 ;
  wire \n27_reg[7]_i_9_n_14 ;
  wire \n27_reg[7]_i_9_n_15 ;
  wire \n27_reg[7]_i_9_n_5 ;
  wire \n27_reg[7]_i_9_n_7 ;
  wire [7:0]n29;
  wire [7:7]n30;
  wire [7:0]n31;
  wire \n33[10]_i_1__4_n_0 ;
  wire \n33[11]_i_1__4_n_0 ;
  wire \n33[12]_i_1__4_n_0 ;
  wire \n33[12]_i_2__4_n_0 ;
  wire \n33[13]_i_1__4_n_0 ;
  wire \n33[14]_i_1__4_n_0 ;
  wire \n33[14]_i_2__4_n_0 ;
  wire \n33[15]_i_2__4_n_0 ;
  wire \n33[2]_i_1__4_n_0 ;
  wire \n33[3]_i_1__4_n_0 ;
  wire \n33[4]_i_1__4_n_0 ;
  wire \n33[4]_i_2__4_n_0 ;
  wire \n33[5]_i_1__4_n_0 ;
  wire \n33[6]_i_1__4_n_0 ;
  wire \n33[6]_i_2__4_n_0 ;
  wire \n33[7]_i_2__4_n_0 ;
  wire \n33[9]_i_1__4_n_0 ;
  wire [7:0]n341_out;
  wire [7:1]n350_out;
  wire \n37[12]_i_2__4_n_0 ;
  wire \n37[14]_i_2__4_n_0 ;
  wire \n37[15]_i_2__4_n_0 ;
  wire \n37[4]_i_2__4_n_0 ;
  wire \n37[6]_i_2__4_n_0 ;
  wire \n37[7]_i_2__4_n_0 ;
  wire \n4_reg_n_0_[0] ;
  wire \n4_reg_n_0_[1] ;
  wire \n4_reg_n_0_[2] ;
  wire \n4_reg_n_0_[3] ;
  wire \n4_reg_n_0_[4] ;
  wire \n4_reg_n_0_[5] ;
  wire \n4_reg_n_0_[6] ;
  wire \n4_reg_n_0_[7] ;
  wire \n7_reg_n_0_[0] ;
  wire \n7_reg_n_0_[1] ;
  wire \n7_reg_n_0_[2] ;
  wire \n7_reg_n_0_[3] ;
  wire \n7_reg_n_0_[4] ;
  wire \n7_reg_n_0_[5] ;
  wire \n7_reg_n_0_[6] ;
  wire \n7_reg_n_0_[7] ;
  wire \n8_reg_n_0_[0] ;
  wire \n8_reg_n_0_[1] ;
  wire \n8_reg_n_0_[2] ;
  wire \n8_reg_n_0_[3] ;
  wire \n8_reg_n_0_[4] ;
  wire \n8_reg_n_0_[5] ;
  wire \n8_reg_n_0_[6] ;
  wire \n8_reg_n_0_[7] ;
  wire \n9_reg_n_0_[0] ;
  wire \n9_reg_n_0_[1] ;
  wire \n9_reg_n_0_[2] ;
  wire \n9_reg_n_0_[3] ;
  wire \n9_reg_n_0_[4] ;
  wire \n9_reg_n_0_[5] ;
  wire \n9_reg_n_0_[6] ;
  wire \n9_reg_n_0_[7] ;
  wire rst_i;
  wire [15:0]s7_3;
  wire [3:0]\NLW_n16_reg[3]_i_1_O_UNCONNECTED ;
  wire [2:1]\NLW_n16_reg[3]_i_17_O_UNCONNECTED ;
  wire [7:3]\NLW_n16_reg[7]_i_1_CO_UNCONNECTED ;
  wire [7:4]\NLW_n16_reg[7]_i_1_O_UNCONNECTED ;
  wire [7:7]\NLW_n16_reg[7]_i_10_CO_UNCONNECTED ;
  wire [0:0]\NLW_n16_reg[7]_i_11_O_UNCONNECTED ;
  wire [7:1]\NLW_n16_reg[7]_i_12_CO_UNCONNECTED ;
  wire [7:2]\NLW_n16_reg[7]_i_12_O_UNCONNECTED ;
  wire [7:1]\NLW_n16_reg[7]_i_9_CO_UNCONNECTED ;
  wire [7:2]\NLW_n16_reg[7]_i_9_O_UNCONNECTED ;
  wire [7:7]\NLW_n21_reg[7]_i_1__0_CO_UNCONNECTED ;
  wire [3:0]\NLW_n27_reg[3]_i_1_O_UNCONNECTED ;
  wire [2:1]\NLW_n27_reg[3]_i_17_O_UNCONNECTED ;
  wire [7:3]\NLW_n27_reg[7]_i_1_CO_UNCONNECTED ;
  wire [7:4]\NLW_n27_reg[7]_i_1_O_UNCONNECTED ;
  wire [7:7]\NLW_n27_reg[7]_i_10_CO_UNCONNECTED ;
  wire [0:0]\NLW_n27_reg[7]_i_11_O_UNCONNECTED ;
  wire [7:1]\NLW_n27_reg[7]_i_12_CO_UNCONNECTED ;
  wire [7:2]\NLW_n27_reg[7]_i_12_O_UNCONNECTED ;
  wire [7:1]\NLW_n27_reg[7]_i_9_CO_UNCONNECTED ;
  wire [7:2]\NLW_n27_reg[7]_i_9_O_UNCONNECTED ;

  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[0] ),
        .Q(n10[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[1] ),
        .Q(n10[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[2] ),
        .Q(n10[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[3] ),
        .Q(n10[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[4] ),
        .Q(n10[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[5] ),
        .Q(n10[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[6] ),
        .Q(n10[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[7] ),
        .Q(n10[7]),
        .R(rst_i));
  (* HLUTNM = "lutpair55" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_10 
       (.I0(\n16_reg[7]_i_10_n_13 ),
        .I1(\n16_reg[7]_i_11_n_9 ),
        .I2(\n16_reg[7]_i_12_n_14 ),
        .I3(\n16[3]_i_3_n_0 ),
        .O(\n16[3]_i_10_n_0 ));
  (* HLUTNM = "lutpair54" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_11 
       (.I0(\n16_reg[7]_i_10_n_14 ),
        .I1(\n16_reg[7]_i_11_n_10 ),
        .I2(\n16_reg[7]_i_12_n_15 ),
        .I3(\n16[3]_i_4_n_0 ),
        .O(\n16[3]_i_11_n_0 ));
  (* HLUTNM = "lutpair53" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_12 
       (.I0(\n16_reg[7]_i_10_n_15 ),
        .I1(\n16_reg[7]_i_11_n_11 ),
        .I2(\n16_reg[3]_i_17_n_8 ),
        .I3(\n16[3]_i_5_n_0 ),
        .O(\n16[3]_i_12_n_0 ));
  (* HLUTNM = "lutpair52" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_13 
       (.I0(n22__6_n_0),
        .I1(\n16_reg[7]_i_11_n_12 ),
        .I2(\n16_reg[3]_i_17_n_9 ),
        .I3(\n16[3]_i_6__0_n_0 ),
        .O(\n16[3]_i_13_n_0 ));
  (* HLUTNM = "lutpair99" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n16[3]_i_14__0 
       (.I0(\n16_reg[7]_i_11_n_13 ),
        .I1(\n16_reg[3]_i_17_n_10 ),
        .I2(\n16_reg[3]_i_17_n_11 ),
        .I3(\n16_reg[7]_i_11_n_14 ),
        .O(\n16[3]_i_14__0_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n16[3]_i_15__0 
       (.I0(\n16_reg[3]_i_17_n_12 ),
        .I1(\n16_reg[3]_i_17_n_15 ),
        .I2(\n16_reg[7]_i_11_n_14 ),
        .I3(\n16_reg[3]_i_17_n_11 ),
        .O(\n16[3]_i_15__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n16[3]_i_16 
       (.I0(\n16_reg[3]_i_17_n_12 ),
        .I1(\n16_reg[3]_i_17_n_15 ),
        .O(\n16[3]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_18 
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(n22__1_n_0),
        .O(\n16[3]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_19 
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__2_n_0),
        .O(\n16[3]_i_19_n_0 ));
  (* HLUTNM = "lutpair55" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_2 
       (.I0(\n16_reg[7]_i_10_n_13 ),
        .I1(\n16_reg[7]_i_11_n_9 ),
        .I2(\n16_reg[7]_i_12_n_14 ),
        .O(\n16[3]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_20 
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(n22__3_n_0),
        .O(\n16[3]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n16[3]_i_21 
       (.I0(n22__4_n_0),
        .I1(n22__5_n_0),
        .I2(n22__3_n_0),
        .O(\n16[3]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h9669)) 
    \n16[3]_i_22 
       (.I0(\n16[7]_i_23__0_n_0 ),
        .I1(n22__0_n_0),
        .I2(n22__1_n_0),
        .I3(n22_n_0),
        .O(\n16[3]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[3]_i_23__0 
       (.I0(n22__3_n_0),
        .I1(n22__1_n_0),
        .I2(n22__2_n_0),
        .I3(n22__0_n_0),
        .O(\n16[3]_i_23__0_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[3]_i_24__0 
       (.I0(n22__4_n_0),
        .I1(n22__2_n_0),
        .I2(n22__3_n_0),
        .I3(n22__1_n_0),
        .O(\n16[3]_i_24__0_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[3]_i_25__0 
       (.I0(n22__5_n_0),
        .I1(n22__3_n_0),
        .I2(n22__4_n_0),
        .I3(n22__2_n_0),
        .O(\n16[3]_i_25__0_n_0 ));
  LUT4 #(
    .INIT(16'h6696)) 
    \n16[3]_i_26__0 
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__5_n_0),
        .I3(n22__6_n_0),
        .O(\n16[3]_i_26__0_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n16[3]_i_27 
       (.I0(n22__6_n_0),
        .I1(n22__5_n_0),
        .I2(n22__4_n_0),
        .O(\n16[3]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n16[3]_i_28__0 
       (.I0(n22__5_n_0),
        .I1(n22__6_n_0),
        .O(\n16[3]_i_28__0_n_0 ));
  (* HLUTNM = "lutpair54" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_3 
       (.I0(\n16_reg[7]_i_10_n_14 ),
        .I1(\n16_reg[7]_i_11_n_10 ),
        .I2(\n16_reg[7]_i_12_n_15 ),
        .O(\n16[3]_i_3_n_0 ));
  (* HLUTNM = "lutpair53" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_4 
       (.I0(\n16_reg[7]_i_10_n_15 ),
        .I1(\n16_reg[7]_i_11_n_11 ),
        .I2(\n16_reg[3]_i_17_n_8 ),
        .O(\n16[3]_i_4_n_0 ));
  (* HLUTNM = "lutpair52" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_5 
       (.I0(n22__6_n_0),
        .I1(\n16_reg[7]_i_11_n_12 ),
        .I2(\n16_reg[3]_i_17_n_9 ),
        .O(\n16[3]_i_5_n_0 ));
  (* HLUTNM = "lutpair99" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \n16[3]_i_6__0 
       (.I0(\n16_reg[7]_i_11_n_13 ),
        .I1(\n16_reg[3]_i_17_n_10 ),
        .O(\n16[3]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n16[3]_i_7 
       (.I0(\n16_reg[3]_i_17_n_11 ),
        .I1(\n16_reg[7]_i_11_n_14 ),
        .O(\n16[3]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n16[3]_i_8 
       (.I0(\n16_reg[3]_i_17_n_12 ),
        .I1(\n16_reg[3]_i_17_n_15 ),
        .O(\n16[3]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_9 
       (.I0(\n16[3]_i_2_n_0 ),
        .I1(\n16_reg[7]_i_11_n_8 ),
        .I2(\n16_reg[7]_i_10_n_12 ),
        .I3(\n16_reg[7]_i_12_n_5 ),
        .O(\n16[3]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \n16[7]_i_13__0 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_13__0_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \n16[7]_i_14 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(\n16[7]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \n16[7]_i_15__0 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_15__0_n_0 ));
  LUT3 #(
    .INIT(8'h4D)) 
    \n16[7]_i_16__0 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(\n16[7]_i_16__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n16[7]_i_17 
       (.I0(n22_n_0),
        .O(\n16[7]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n16[7]_i_18 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n16[7]_i_19__0 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .O(\n16[7]_i_19__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n16[7]_i_2 
       (.I0(\n16_reg[7]_i_9_n_14 ),
        .I1(\n16_reg[7]_i_10_n_10 ),
        .O(\n16[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n16[7]_i_20__0 
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .O(\n16[7]_i_20__0_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n16[7]_i_21__0 
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .O(\n16[7]_i_21__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n16[7]_i_22 
       (.I0(n22__5_n_0),
        .O(\n16[7]_i_22_n_0 ));
  (* HLUTNM = "lutpair98" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_23__0 
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .O(\n16[7]_i_23__0_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_24 
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(n22__1_n_0),
        .O(\n16[7]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_25 
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__2_n_0),
        .O(\n16[7]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_26 
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(n22__3_n_0),
        .O(\n16[7]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n16[7]_i_27 
       (.I0(n22__4_n_0),
        .I1(n22__5_n_0),
        .I2(n22__3_n_0),
        .O(\n16[7]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h9669)) 
    \n16[7]_i_28 
       (.I0(\n16[7]_i_23__0_n_0 ),
        .I1(n22__0_n_0),
        .I2(n22__1_n_0),
        .I3(n22_n_0),
        .O(\n16[7]_i_28_n_0 ));
  (* HLUTNM = "lutpair98" *) 
  LUT4 #(
    .INIT(16'h781E)) 
    \n16[7]_i_29__0 
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(n22__3_n_0),
        .O(\n16[7]_i_29__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n16[7]_i_3 
       (.I0(\n16_reg[7]_i_9_n_15 ),
        .I1(\n16_reg[7]_i_10_n_11 ),
        .O(\n16[7]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[7]_i_30__0 
       (.I0(n22__4_n_0),
        .I1(n22__2_n_0),
        .I2(n22__3_n_0),
        .I3(n22__1_n_0),
        .O(\n16[7]_i_30__0_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[7]_i_31__0 
       (.I0(n22__5_n_0),
        .I1(n22__3_n_0),
        .I2(n22__4_n_0),
        .I3(n22__2_n_0),
        .O(\n16[7]_i_31__0_n_0 ));
  LUT4 #(
    .INIT(16'h6696)) 
    \n16[7]_i_32__0 
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__5_n_0),
        .I3(n22__6_n_0),
        .O(\n16[7]_i_32__0_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n16[7]_i_33 
       (.I0(n22__6_n_0),
        .I1(n22__5_n_0),
        .I2(n22__4_n_0),
        .O(\n16[7]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n16[7]_i_34__0 
       (.I0(n22__5_n_0),
        .I1(n22__6_n_0),
        .O(\n16[7]_i_34__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \n16[7]_i_35__0 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_35__0_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \n16[7]_i_36 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(\n16[7]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \n16[7]_i_37__0 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_37__0_n_0 ));
  LUT3 #(
    .INIT(8'h4D)) 
    \n16[7]_i_38__0 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(\n16[7]_i_38__0_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_4 
       (.I0(\n16_reg[7]_i_10_n_12 ),
        .I1(\n16_reg[7]_i_11_n_8 ),
        .I2(\n16_reg[7]_i_12_n_5 ),
        .O(\n16[7]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \n16[7]_i_5__0 
       (.I0(\n16_reg[7]_i_9_n_5 ),
        .I1(\n16_reg[7]_i_10_n_9 ),
        .I2(\n16_reg[7]_i_10_n_8 ),
        .O(\n16[7]_i_5__0_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n16[7]_i_6__0 
       (.I0(\n16_reg[7]_i_9_n_14 ),
        .I1(\n16_reg[7]_i_10_n_10 ),
        .I2(\n16_reg[7]_i_10_n_9 ),
        .I3(\n16_reg[7]_i_9_n_5 ),
        .O(\n16[7]_i_6__0_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n16[7]_i_7__0 
       (.I0(\n16_reg[7]_i_9_n_15 ),
        .I1(\n16_reg[7]_i_10_n_11 ),
        .I2(\n16_reg[7]_i_10_n_10 ),
        .I3(\n16_reg[7]_i_9_n_14 ),
        .O(\n16[7]_i_7__0_n_0 ));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    \n16[7]_i_8 
       (.I0(\n16_reg[7]_i_12_n_5 ),
        .I1(\n16_reg[7]_i_11_n_8 ),
        .I2(\n16_reg[7]_i_10_n_12 ),
        .I3(\n16_reg[7]_i_10_n_11 ),
        .I4(\n16_reg[7]_i_9_n_15 ),
        .O(\n16[7]_i_8_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[0]),
        .Q(\n16_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[1]),
        .Q(\n16_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[2]),
        .Q(\n16_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[3]),
        .Q(\n16_reg_n_0_[3] ),
        .R(rst_i));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[3]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n16_reg[3]_i_1_n_0 ,\n16_reg[3]_i_1_n_1 ,\n16_reg[3]_i_1_n_2 ,\n16_reg[3]_i_1_n_3 ,\n16_reg[3]_i_1_n_4 ,\n16_reg[3]_i_1_n_5 ,\n16_reg[3]_i_1_n_6 ,\n16_reg[3]_i_1_n_7 }),
        .DI({\n16[3]_i_2_n_0 ,\n16[3]_i_3_n_0 ,\n16[3]_i_4_n_0 ,\n16[3]_i_5_n_0 ,\n16[3]_i_6__0_n_0 ,\n16[3]_i_7_n_0 ,\n16[3]_i_8_n_0 ,1'b0}),
        .O({n15[3:0],\NLW_n16_reg[3]_i_1_O_UNCONNECTED [3:0]}),
        .S({\n16[3]_i_9_n_0 ,\n16[3]_i_10_n_0 ,\n16[3]_i_11_n_0 ,\n16[3]_i_12_n_0 ,\n16[3]_i_13_n_0 ,\n16[3]_i_14__0_n_0 ,\n16[3]_i_15__0_n_0 ,\n16[3]_i_16_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[3]_i_17 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n16_reg[3]_i_17_n_0 ,\n16_reg[3]_i_17_n_1 ,\n16_reg[3]_i_17_n_2 ,\n16_reg[3]_i_17_n_3 ,\n16_reg[3]_i_17_n_4 ,\n16_reg[3]_i_17_n_5 ,\n16_reg[3]_i_17_n_6 ,\n16_reg[3]_i_17_n_7 }),
        .DI({\n16[7]_i_23__0_n_0 ,\n16[3]_i_18_n_0 ,\n16[3]_i_19_n_0 ,\n16[3]_i_20_n_0 ,\n16[3]_i_21_n_0 ,n22__4_n_0,n22__5_n_0,1'b0}),
        .O({\n16_reg[3]_i_17_n_8 ,\n16_reg[3]_i_17_n_9 ,\n16_reg[3]_i_17_n_10 ,\n16_reg[3]_i_17_n_11 ,\n16_reg[3]_i_17_n_12 ,\NLW_n16_reg[3]_i_17_O_UNCONNECTED [2:1],\n16_reg[3]_i_17_n_15 }),
        .S({\n16[3]_i_22_n_0 ,\n16[3]_i_23__0_n_0 ,\n16[3]_i_24__0_n_0 ,\n16[3]_i_25__0_n_0 ,\n16[3]_i_26__0_n_0 ,\n16[3]_i_27_n_0 ,\n16[3]_i_28__0_n_0 ,n22__6_n_0}));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[4]),
        .Q(\n16_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[5]),
        .Q(\n16_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[6]),
        .Q(\n16_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[7]),
        .Q(\n16_reg_n_0_[7] ),
        .R(rst_i));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_1 
       (.CI(\n16_reg[3]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n16_reg[7]_i_1_CO_UNCONNECTED [7:3],\n16_reg[7]_i_1_n_5 ,\n16_reg[7]_i_1_n_6 ,\n16_reg[7]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,\n16[7]_i_2_n_0 ,\n16[7]_i_3_n_0 ,\n16[7]_i_4_n_0 }),
        .O({\NLW_n16_reg[7]_i_1_O_UNCONNECTED [7:4],n15[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,\n16[7]_i_5__0_n_0 ,\n16[7]_i_6__0_n_0 ,\n16[7]_i_7__0_n_0 ,\n16[7]_i_8_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_10 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\NLW_n16_reg[7]_i_10_CO_UNCONNECTED [7],\n16_reg[7]_i_10_n_1 ,\n16_reg[7]_i_10_n_2 ,\n16_reg[7]_i_10_n_3 ,\n16_reg[7]_i_10_n_4 ,\n16_reg[7]_i_10_n_5 ,\n16_reg[7]_i_10_n_6 ,\n16_reg[7]_i_10_n_7 }),
        .DI({1'b0,n22__0_n_0,n22__1_n_0,n22__2_n_0,n22__3_n_0,1'b1,1'b0,1'b1}),
        .O({\n16_reg[7]_i_10_n_8 ,\n16_reg[7]_i_10_n_9 ,\n16_reg[7]_i_10_n_10 ,\n16_reg[7]_i_10_n_11 ,\n16_reg[7]_i_10_n_12 ,\n16_reg[7]_i_10_n_13 ,\n16_reg[7]_i_10_n_14 ,\n16_reg[7]_i_10_n_15 }),
        .S({\n16[7]_i_17_n_0 ,\n16[7]_i_18_n_0 ,\n16[7]_i_19__0_n_0 ,\n16[7]_i_20__0_n_0 ,\n16[7]_i_21__0_n_0 ,n22__3_n_0,n22__4_n_0,\n16[7]_i_22_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_11 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n16_reg[7]_i_11_n_0 ,\n16_reg[7]_i_11_n_1 ,\n16_reg[7]_i_11_n_2 ,\n16_reg[7]_i_11_n_3 ,\n16_reg[7]_i_11_n_4 ,\n16_reg[7]_i_11_n_5 ,\n16_reg[7]_i_11_n_6 ,\n16_reg[7]_i_11_n_7 }),
        .DI({\n16[7]_i_23__0_n_0 ,\n16[7]_i_24_n_0 ,\n16[7]_i_25_n_0 ,\n16[7]_i_26_n_0 ,\n16[7]_i_27_n_0 ,n22__4_n_0,n22__5_n_0,1'b0}),
        .O({\n16_reg[7]_i_11_n_8 ,\n16_reg[7]_i_11_n_9 ,\n16_reg[7]_i_11_n_10 ,\n16_reg[7]_i_11_n_11 ,\n16_reg[7]_i_11_n_12 ,\n16_reg[7]_i_11_n_13 ,\n16_reg[7]_i_11_n_14 ,\NLW_n16_reg[7]_i_11_O_UNCONNECTED [0]}),
        .S({\n16[7]_i_28_n_0 ,\n16[7]_i_29__0_n_0 ,\n16[7]_i_30__0_n_0 ,\n16[7]_i_31__0_n_0 ,\n16[7]_i_32__0_n_0 ,\n16[7]_i_33_n_0 ,\n16[7]_i_34__0_n_0 ,n22__6_n_0}));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_12 
       (.CI(\n16_reg[3]_i_17_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n16_reg[7]_i_12_CO_UNCONNECTED [7:3],\n16_reg[7]_i_12_n_5 ,\NLW_n16_reg[7]_i_12_CO_UNCONNECTED [1],\n16_reg[7]_i_12_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\n16[7]_i_35__0_n_0 ,\n16[7]_i_36_n_0 }),
        .O({\NLW_n16_reg[7]_i_12_O_UNCONNECTED [7:2],\n16_reg[7]_i_12_n_14 ,\n16_reg[7]_i_12_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,\n16[7]_i_37__0_n_0 ,\n16[7]_i_38__0_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_9 
       (.CI(\n16_reg[7]_i_11_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n16_reg[7]_i_9_CO_UNCONNECTED [7:3],\n16_reg[7]_i_9_n_5 ,\NLW_n16_reg[7]_i_9_CO_UNCONNECTED [1],\n16_reg[7]_i_9_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\n16[7]_i_13__0_n_0 ,\n16[7]_i_14_n_0 }),
        .O({\NLW_n16_reg[7]_i_9_O_UNCONNECTED [7:2],\n16_reg[7]_i_9_n_14 ,\n16_reg[7]_i_9_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,\n16[7]_i_15__0_n_0 ,\n16[7]_i_16__0_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[0]),
        .Q(\n1_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[10]),
        .Q(n2[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[11]),
        .Q(n2[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[12]),
        .Q(n2[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[13]),
        .Q(n2[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[14]),
        .Q(n2[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[15]),
        .Q(n2[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[1]),
        .Q(\n1_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[2]),
        .Q(\n1_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[3]),
        .Q(\n1_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[4]),
        .Q(\n1_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[5]),
        .Q(\n1_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[6]),
        .Q(\n1_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[7]),
        .Q(\n1_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[8]),
        .Q(n2[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[9]),
        .Q(n2[1]),
        .R(rst_i));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_2__0 
       (.I0(\n16_reg_n_0_[7] ),
        .O(\n21[7]_i_2__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_3__0 
       (.I0(\n16_reg_n_0_[6] ),
        .O(\n21[7]_i_3__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_4__0 
       (.I0(\n16_reg_n_0_[5] ),
        .O(\n21[7]_i_4__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_5__0 
       (.I0(\n16_reg_n_0_[4] ),
        .O(\n21[7]_i_5__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_6__0 
       (.I0(\n16_reg_n_0_[3] ),
        .O(\n21[7]_i_6__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_7__0 
       (.I0(\n16_reg_n_0_[2] ),
        .O(\n21[7]_i_7__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_8__0 
       (.I0(\n16_reg_n_0_[1] ),
        .O(\n21[7]_i_8__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_9__0 
       (.I0(\n16_reg_n_0_[0] ),
        .O(\n21[7]_i_9__0_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[0]),
        .Q(n21[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[1]),
        .Q(n21[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[2]),
        .Q(n21[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[3]),
        .Q(n21[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[4]),
        .Q(n21[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[5]),
        .Q(n21[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[6]),
        .Q(n21[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[7]),
        .Q(n21[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n21_reg[7]_i_1__0 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\NLW_n21_reg[7]_i_1__0_CO_UNCONNECTED [7],\n21_reg[7]_i_1__0_n_1 ,\n21_reg[7]_i_1__0_n_2 ,\n21_reg[7]_i_1__0_n_3 ,\n21_reg[7]_i_1__0_n_4 ,\n21_reg[7]_i_1__0_n_5 ,\n21_reg[7]_i_1__0_n_6 ,\n21_reg[7]_i_1__0_n_7 }),
        .DI({1'b0,\n16_reg_n_0_[6] ,\n16_reg_n_0_[5] ,\n16_reg_n_0_[4] ,\n16_reg_n_0_[3] ,\n16_reg_n_0_[2] ,\n16_reg_n_0_[1] ,\n16_reg_n_0_[0] }),
        .O(n202_out),
        .S({\n21[7]_i_2__0_n_0 ,\n21[7]_i_3__0_n_0 ,\n21[7]_i_4__0_n_0 ,\n21[7]_i_5__0_n_0 ,\n21[7]_i_6__0_n_0 ,\n21[7]_i_7__0_n_0 ,\n21[7]_i_8__0_n_0 ,\n21[7]_i_9__0_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    n22
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[15]),
        .Q(n22_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__0
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[14]),
        .Q(n22__0_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__1
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[13]),
        .Q(n22__1_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__2
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[12]),
        .Q(n22__2_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__3
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[11]),
        .Q(n22__3_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__4
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[10]),
        .Q(n22__4_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__5
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[9]),
        .Q(n22__5_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__6
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[8]),
        .Q(n22__6_n_0),
        .R(rst_i));
  (* HLUTNM = "lutpair51" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_10 
       (.I0(\n27_reg[7]_i_10_n_13 ),
        .I1(\n27_reg[7]_i_11_n_9 ),
        .I2(\n27_reg[7]_i_12_n_14 ),
        .I3(\n27[3]_i_3_n_0 ),
        .O(\n27[3]_i_10_n_0 ));
  (* HLUTNM = "lutpair50" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_11 
       (.I0(\n27_reg[7]_i_10_n_14 ),
        .I1(\n27_reg[7]_i_11_n_10 ),
        .I2(\n27_reg[7]_i_12_n_15 ),
        .I3(\n27[3]_i_4_n_0 ),
        .O(\n27[3]_i_11_n_0 ));
  (* HLUTNM = "lutpair49" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_12 
       (.I0(\n27_reg[7]_i_10_n_15 ),
        .I1(\n27_reg[7]_i_11_n_11 ),
        .I2(\n27_reg[3]_i_17_n_8 ),
        .I3(\n27[3]_i_5_n_0 ),
        .O(\n27[3]_i_12_n_0 ));
  (* HLUTNM = "lutpair48" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_13 
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n27_reg[7]_i_11_n_12 ),
        .I2(\n27_reg[3]_i_17_n_9 ),
        .I3(\n27[3]_i_6__0_n_0 ),
        .O(\n27[3]_i_13_n_0 ));
  (* HLUTNM = "lutpair97" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n27[3]_i_14__0 
       (.I0(\n27_reg[7]_i_11_n_13 ),
        .I1(\n27_reg[3]_i_17_n_10 ),
        .I2(\n27_reg[3]_i_17_n_11 ),
        .I3(\n27_reg[7]_i_11_n_14 ),
        .O(\n27[3]_i_14__0_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n27[3]_i_15__0 
       (.I0(\n27_reg[3]_i_17_n_12 ),
        .I1(\n27_reg[3]_i_17_n_15 ),
        .I2(\n27_reg[7]_i_11_n_14 ),
        .I3(\n27_reg[3]_i_17_n_11 ),
        .O(\n27[3]_i_15__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n27[3]_i_16 
       (.I0(\n27_reg[3]_i_17_n_12 ),
        .I1(\n27_reg[3]_i_17_n_15 ),
        .O(\n27[3]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_18 
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[5] ),
        .O(\n27[3]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_19 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[4] ),
        .O(\n27[3]_i_19_n_0 ));
  (* HLUTNM = "lutpair51" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_2 
       (.I0(\n27_reg[7]_i_10_n_13 ),
        .I1(\n27_reg[7]_i_11_n_9 ),
        .I2(\n27_reg[7]_i_12_n_14 ),
        .O(\n27[3]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_20 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[2] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(\n27[3]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n27[3]_i_21 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(\n27[3]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h9669)) 
    \n27[3]_i_22 
       (.I0(\n27[7]_i_23__0_n_0 ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[5] ),
        .I3(\n4_reg_n_0_[7] ),
        .O(\n27[3]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[3]_i_23__0 
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[5] ),
        .I2(\n4_reg_n_0_[4] ),
        .I3(\n4_reg_n_0_[6] ),
        .O(\n27[3]_i_23__0_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[3]_i_24__0 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[3] ),
        .I3(\n4_reg_n_0_[5] ),
        .O(\n27[3]_i_24__0_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[3]_i_25__0 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[2] ),
        .I3(\n4_reg_n_0_[4] ),
        .O(\n27[3]_i_25__0_n_0 ));
  LUT4 #(
    .INIT(16'h6696)) 
    \n27[3]_i_26__0 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[1] ),
        .I3(\n4_reg_n_0_[0] ),
        .O(\n27[3]_i_26__0_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n27[3]_i_27 
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[2] ),
        .O(\n27[3]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n27[3]_i_28__0 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[0] ),
        .O(\n27[3]_i_28__0_n_0 ));
  (* HLUTNM = "lutpair50" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_3 
       (.I0(\n27_reg[7]_i_10_n_14 ),
        .I1(\n27_reg[7]_i_11_n_10 ),
        .I2(\n27_reg[7]_i_12_n_15 ),
        .O(\n27[3]_i_3_n_0 ));
  (* HLUTNM = "lutpair49" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_4 
       (.I0(\n27_reg[7]_i_10_n_15 ),
        .I1(\n27_reg[7]_i_11_n_11 ),
        .I2(\n27_reg[3]_i_17_n_8 ),
        .O(\n27[3]_i_4_n_0 ));
  (* HLUTNM = "lutpair48" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_5 
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n27_reg[7]_i_11_n_12 ),
        .I2(\n27_reg[3]_i_17_n_9 ),
        .O(\n27[3]_i_5_n_0 ));
  (* HLUTNM = "lutpair97" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \n27[3]_i_6__0 
       (.I0(\n27_reg[7]_i_11_n_13 ),
        .I1(\n27_reg[3]_i_17_n_10 ),
        .O(\n27[3]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n27[3]_i_7 
       (.I0(\n27_reg[3]_i_17_n_11 ),
        .I1(\n27_reg[7]_i_11_n_14 ),
        .O(\n27[3]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n27[3]_i_8 
       (.I0(\n27_reg[3]_i_17_n_12 ),
        .I1(\n27_reg[3]_i_17_n_15 ),
        .O(\n27[3]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_9 
       (.I0(\n27[3]_i_2_n_0 ),
        .I1(\n27_reg[7]_i_11_n_8 ),
        .I2(\n27_reg[7]_i_10_n_12 ),
        .I3(\n27_reg[7]_i_12_n_5 ),
        .O(\n27[3]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \n27[7]_i_13__0 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_13__0_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \n27[7]_i_14 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \n27[7]_i_15__0 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_15__0_n_0 ));
  LUT3 #(
    .INIT(8'h4D)) 
    \n27[7]_i_16__0 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_16__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n27[7]_i_17 
       (.I0(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n27[7]_i_18 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n27[7]_i_19__0 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .O(\n27[7]_i_19__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n27[7]_i_2 
       (.I0(\n27_reg[7]_i_9_n_14 ),
        .I1(\n27_reg[7]_i_10_n_10 ),
        .O(\n27[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n27[7]_i_20__0 
       (.I0(\n4_reg_n_0_[4] ),
        .I1(\n4_reg_n_0_[5] ),
        .O(\n27[7]_i_20__0_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n27[7]_i_21__0 
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[4] ),
        .O(\n27[7]_i_21__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n27[7]_i_22 
       (.I0(\n4_reg_n_0_[1] ),
        .O(\n27[7]_i_22_n_0 ));
  (* HLUTNM = "lutpair96" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_23__0 
       (.I0(\n4_reg_n_0_[4] ),
        .I1(\n4_reg_n_0_[5] ),
        .I2(\n4_reg_n_0_[6] ),
        .O(\n27[7]_i_23__0_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_24 
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[5] ),
        .O(\n27[7]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_25 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[4] ),
        .O(\n27[7]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_26 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[2] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(\n27[7]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n27[7]_i_27 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(\n27[7]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h9669)) 
    \n27[7]_i_28 
       (.I0(\n27[7]_i_23__0_n_0 ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[5] ),
        .I3(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_28_n_0 ));
  (* HLUTNM = "lutpair96" *) 
  LUT4 #(
    .INIT(16'h781E)) 
    \n27[7]_i_29__0 
       (.I0(\n4_reg_n_0_[4] ),
        .I1(\n4_reg_n_0_[5] ),
        .I2(\n4_reg_n_0_[6] ),
        .I3(\n4_reg_n_0_[3] ),
        .O(\n27[7]_i_29__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n27[7]_i_3 
       (.I0(\n27_reg[7]_i_9_n_15 ),
        .I1(\n27_reg[7]_i_10_n_11 ),
        .O(\n27[7]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[7]_i_30__0 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[3] ),
        .I3(\n4_reg_n_0_[5] ),
        .O(\n27[7]_i_30__0_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[7]_i_31__0 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[2] ),
        .I3(\n4_reg_n_0_[4] ),
        .O(\n27[7]_i_31__0_n_0 ));
  LUT4 #(
    .INIT(16'h6696)) 
    \n27[7]_i_32__0 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[1] ),
        .I3(\n4_reg_n_0_[0] ),
        .O(\n27[7]_i_32__0_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n27[7]_i_33 
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[2] ),
        .O(\n27[7]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n27[7]_i_34__0 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[0] ),
        .O(\n27[7]_i_34__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \n27[7]_i_35__0 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_35__0_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \n27[7]_i_36 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \n27[7]_i_37__0 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_37__0_n_0 ));
  LUT3 #(
    .INIT(8'h4D)) 
    \n27[7]_i_38__0 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_38__0_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_4 
       (.I0(\n27_reg[7]_i_10_n_12 ),
        .I1(\n27_reg[7]_i_11_n_8 ),
        .I2(\n27_reg[7]_i_12_n_5 ),
        .O(\n27[7]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \n27[7]_i_5__0 
       (.I0(\n27_reg[7]_i_9_n_5 ),
        .I1(\n27_reg[7]_i_10_n_9 ),
        .I2(\n27_reg[7]_i_10_n_8 ),
        .O(\n27[7]_i_5__0_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n27[7]_i_6__0 
       (.I0(\n27_reg[7]_i_9_n_14 ),
        .I1(\n27_reg[7]_i_10_n_10 ),
        .I2(\n27_reg[7]_i_10_n_9 ),
        .I3(\n27_reg[7]_i_9_n_5 ),
        .O(\n27[7]_i_6__0_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n27[7]_i_7__0 
       (.I0(\n27_reg[7]_i_9_n_15 ),
        .I1(\n27_reg[7]_i_10_n_11 ),
        .I2(\n27_reg[7]_i_10_n_10 ),
        .I3(\n27_reg[7]_i_9_n_14 ),
        .O(\n27[7]_i_7__0_n_0 ));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    \n27[7]_i_8 
       (.I0(\n27_reg[7]_i_12_n_5 ),
        .I1(\n27_reg[7]_i_11_n_8 ),
        .I2(\n27_reg[7]_i_10_n_12 ),
        .I3(\n27_reg[7]_i_10_n_11 ),
        .I4(\n27_reg[7]_i_9_n_15 ),
        .O(\n27[7]_i_8_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[0]),
        .Q(n27[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[1]),
        .Q(n27[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[2]),
        .Q(n27[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[3]),
        .Q(n27[3]),
        .R(rst_i));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[3]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n27_reg[3]_i_1_n_0 ,\n27_reg[3]_i_1_n_1 ,\n27_reg[3]_i_1_n_2 ,\n27_reg[3]_i_1_n_3 ,\n27_reg[3]_i_1_n_4 ,\n27_reg[3]_i_1_n_5 ,\n27_reg[3]_i_1_n_6 ,\n27_reg[3]_i_1_n_7 }),
        .DI({\n27[3]_i_2_n_0 ,\n27[3]_i_3_n_0 ,\n27[3]_i_4_n_0 ,\n27[3]_i_5_n_0 ,\n27[3]_i_6__0_n_0 ,\n27[3]_i_7_n_0 ,\n27[3]_i_8_n_0 ,1'b0}),
        .O({n26[3:0],\NLW_n27_reg[3]_i_1_O_UNCONNECTED [3:0]}),
        .S({\n27[3]_i_9_n_0 ,\n27[3]_i_10_n_0 ,\n27[3]_i_11_n_0 ,\n27[3]_i_12_n_0 ,\n27[3]_i_13_n_0 ,\n27[3]_i_14__0_n_0 ,\n27[3]_i_15__0_n_0 ,\n27[3]_i_16_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[3]_i_17 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n27_reg[3]_i_17_n_0 ,\n27_reg[3]_i_17_n_1 ,\n27_reg[3]_i_17_n_2 ,\n27_reg[3]_i_17_n_3 ,\n27_reg[3]_i_17_n_4 ,\n27_reg[3]_i_17_n_5 ,\n27_reg[3]_i_17_n_6 ,\n27_reg[3]_i_17_n_7 }),
        .DI({\n27[7]_i_23__0_n_0 ,\n27[3]_i_18_n_0 ,\n27[3]_i_19_n_0 ,\n27[3]_i_20_n_0 ,\n27[3]_i_21_n_0 ,\n4_reg_n_0_[2] ,\n4_reg_n_0_[1] ,1'b0}),
        .O({\n27_reg[3]_i_17_n_8 ,\n27_reg[3]_i_17_n_9 ,\n27_reg[3]_i_17_n_10 ,\n27_reg[3]_i_17_n_11 ,\n27_reg[3]_i_17_n_12 ,\NLW_n27_reg[3]_i_17_O_UNCONNECTED [2:1],\n27_reg[3]_i_17_n_15 }),
        .S({\n27[3]_i_22_n_0 ,\n27[3]_i_23__0_n_0 ,\n27[3]_i_24__0_n_0 ,\n27[3]_i_25__0_n_0 ,\n27[3]_i_26__0_n_0 ,\n27[3]_i_27_n_0 ,\n27[3]_i_28__0_n_0 ,\n4_reg_n_0_[0] }));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[4]),
        .Q(n27[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[5]),
        .Q(n27[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[6]),
        .Q(n27[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[7]),
        .Q(n27[7]),
        .R(rst_i));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_1 
       (.CI(\n27_reg[3]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n27_reg[7]_i_1_CO_UNCONNECTED [7:3],\n27_reg[7]_i_1_n_5 ,\n27_reg[7]_i_1_n_6 ,\n27_reg[7]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,\n27[7]_i_2_n_0 ,\n27[7]_i_3_n_0 ,\n27[7]_i_4_n_0 }),
        .O({\NLW_n27_reg[7]_i_1_O_UNCONNECTED [7:4],n26[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,\n27[7]_i_5__0_n_0 ,\n27[7]_i_6__0_n_0 ,\n27[7]_i_7__0_n_0 ,\n27[7]_i_8_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_10 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\NLW_n27_reg[7]_i_10_CO_UNCONNECTED [7],\n27_reg[7]_i_10_n_1 ,\n27_reg[7]_i_10_n_2 ,\n27_reg[7]_i_10_n_3 ,\n27_reg[7]_i_10_n_4 ,\n27_reg[7]_i_10_n_5 ,\n27_reg[7]_i_10_n_6 ,\n27_reg[7]_i_10_n_7 }),
        .DI({1'b0,\n4_reg_n_0_[6] ,\n4_reg_n_0_[5] ,\n4_reg_n_0_[4] ,\n4_reg_n_0_[3] ,1'b1,1'b0,1'b1}),
        .O({\n27_reg[7]_i_10_n_8 ,\n27_reg[7]_i_10_n_9 ,\n27_reg[7]_i_10_n_10 ,\n27_reg[7]_i_10_n_11 ,\n27_reg[7]_i_10_n_12 ,\n27_reg[7]_i_10_n_13 ,\n27_reg[7]_i_10_n_14 ,\n27_reg[7]_i_10_n_15 }),
        .S({\n27[7]_i_17_n_0 ,\n27[7]_i_18_n_0 ,\n27[7]_i_19__0_n_0 ,\n27[7]_i_20__0_n_0 ,\n27[7]_i_21__0_n_0 ,\n4_reg_n_0_[3] ,\n4_reg_n_0_[2] ,\n27[7]_i_22_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_11 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n27_reg[7]_i_11_n_0 ,\n27_reg[7]_i_11_n_1 ,\n27_reg[7]_i_11_n_2 ,\n27_reg[7]_i_11_n_3 ,\n27_reg[7]_i_11_n_4 ,\n27_reg[7]_i_11_n_5 ,\n27_reg[7]_i_11_n_6 ,\n27_reg[7]_i_11_n_7 }),
        .DI({\n27[7]_i_23__0_n_0 ,\n27[7]_i_24_n_0 ,\n27[7]_i_25_n_0 ,\n27[7]_i_26_n_0 ,\n27[7]_i_27_n_0 ,\n4_reg_n_0_[2] ,\n4_reg_n_0_[1] ,1'b0}),
        .O({\n27_reg[7]_i_11_n_8 ,\n27_reg[7]_i_11_n_9 ,\n27_reg[7]_i_11_n_10 ,\n27_reg[7]_i_11_n_11 ,\n27_reg[7]_i_11_n_12 ,\n27_reg[7]_i_11_n_13 ,\n27_reg[7]_i_11_n_14 ,\NLW_n27_reg[7]_i_11_O_UNCONNECTED [0]}),
        .S({\n27[7]_i_28_n_0 ,\n27[7]_i_29__0_n_0 ,\n27[7]_i_30__0_n_0 ,\n27[7]_i_31__0_n_0 ,\n27[7]_i_32__0_n_0 ,\n27[7]_i_33_n_0 ,\n27[7]_i_34__0_n_0 ,\n4_reg_n_0_[0] }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_12 
       (.CI(\n27_reg[3]_i_17_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n27_reg[7]_i_12_CO_UNCONNECTED [7:3],\n27_reg[7]_i_12_n_5 ,\NLW_n27_reg[7]_i_12_CO_UNCONNECTED [1],\n27_reg[7]_i_12_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\n27[7]_i_35__0_n_0 ,\n27[7]_i_36_n_0 }),
        .O({\NLW_n27_reg[7]_i_12_O_UNCONNECTED [7:2],\n27_reg[7]_i_12_n_14 ,\n27_reg[7]_i_12_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,\n27[7]_i_37__0_n_0 ,\n27[7]_i_38__0_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_9 
       (.CI(\n27_reg[7]_i_11_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n27_reg[7]_i_9_CO_UNCONNECTED [7:3],\n27_reg[7]_i_9_n_5 ,\NLW_n27_reg[7]_i_9_CO_UNCONNECTED [1],\n27_reg[7]_i_9_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\n27[7]_i_13__0_n_0 ,\n27[7]_i_14_n_0 }),
        .O({\NLW_n27_reg[7]_i_9_O_UNCONNECTED [7:2],\n27_reg[7]_i_9_n_14 ,\n27_reg[7]_i_9_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,\n27[7]_i_15__0_n_0 ,\n27[7]_i_16__0_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[0]),
        .Q(n29[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[1]),
        .Q(n29[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[2]),
        .Q(n29[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[3]),
        .Q(n29[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[4]),
        .Q(n29[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[5]),
        .Q(n29[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[6]),
        .Q(n29[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[7]),
        .Q(n29[7]),
        .R(rst_i));
  LUT2 #(
    .INIT(4'h6)) 
    \n33[0]_i_1__4 
       (.I0(n29[0]),
        .I1(n10[0]),
        .O(n31[0]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[10]_i_1__4 
       (.I0(n21[2]),
        .I1(\n8_reg_n_0_[2] ),
        .I2(\n8_reg_n_0_[1] ),
        .I3(n21[1]),
        .I4(\n8_reg_n_0_[0] ),
        .I5(n21[0]),
        .O(\n33[10]_i_1__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[11]_i_1__4 
       (.I0(n21[3]),
        .I1(\n8_reg_n_0_[3] ),
        .I2(\n33[12]_i_2__4_n_0 ),
        .O(\n33[11]_i_1__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[12]_i_1__4 
       (.I0(n21[4]),
        .I1(\n8_reg_n_0_[4] ),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[3]),
        .I4(\n33[12]_i_2__4_n_0 ),
        .O(\n33[12]_i_1__4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[12]_i_2__4 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n33[12]_i_2__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[13]_i_1__4 
       (.I0(n21[5]),
        .I1(\n8_reg_n_0_[5] ),
        .I2(\n33[14]_i_2__4_n_0 ),
        .O(\n33[13]_i_1__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[14]_i_1__4 
       (.I0(n21[6]),
        .I1(\n8_reg_n_0_[6] ),
        .I2(\n8_reg_n_0_[5] ),
        .I3(n21[5]),
        .I4(\n33[14]_i_2__4_n_0 ),
        .O(\n33[14]_i_1__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[14]_i_2__4 
       (.I0(\n33[12]_i_2__4_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n33[14]_i_2__4_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[15]_i_1__4 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n33[15]_i_2__4_n_0 ),
        .O(n30));
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[15]_i_2__4 
       (.I0(\n33[14]_i_2__4_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n33[15]_i_2__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[1]_i_1__4 
       (.I0(n29[1]),
        .I1(n10[1]),
        .I2(n10[0]),
        .I3(n29[0]),
        .O(n31[1]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[2]_i_1__4 
       (.I0(n29[2]),
        .I1(n10[2]),
        .I2(n10[1]),
        .I3(n29[1]),
        .I4(n10[0]),
        .I5(n29[0]),
        .O(\n33[2]_i_1__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[3]_i_1__4 
       (.I0(n29[3]),
        .I1(n10[3]),
        .I2(\n33[4]_i_2__4_n_0 ),
        .O(\n33[3]_i_1__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[4]_i_1__4 
       (.I0(n29[4]),
        .I1(n10[4]),
        .I2(n10[3]),
        .I3(n29[3]),
        .I4(\n33[4]_i_2__4_n_0 ),
        .O(\n33[4]_i_1__4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[4]_i_2__4 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n33[4]_i_2__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[5]_i_1__4 
       (.I0(n29[5]),
        .I1(n10[5]),
        .I2(\n33[6]_i_2__4_n_0 ),
        .O(\n33[5]_i_1__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[6]_i_1__4 
       (.I0(n29[6]),
        .I1(n10[6]),
        .I2(n10[5]),
        .I3(n29[5]),
        .I4(\n33[6]_i_2__4_n_0 ),
        .O(\n33[6]_i_1__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[6]_i_2__4 
       (.I0(\n33[4]_i_2__4_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n33[6]_i_2__4_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[7]_i_1__4 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n33[7]_i_2__4_n_0 ),
        .O(n31[7]));
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[7]_i_2__4 
       (.I0(\n33[6]_i_2__4_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n33[7]_i_2__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[9]_i_1__4 
       (.I0(n21[1]),
        .I1(\n8_reg_n_0_[1] ),
        .I2(\n8_reg_n_0_[0] ),
        .I3(n21[0]),
        .O(\n33[9]_i_1__4_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[0]),
        .Q(i1[15]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[10]_i_1__4_n_0 ),
        .Q(i1[24]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[11]_i_1__4_n_0 ),
        .Q(i1[25]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[12]_i_1__4_n_0 ),
        .Q(i1[26]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[13]_i_1__4_n_0 ),
        .Q(i1[27]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[14]_i_1__4_n_0 ),
        .Q(i1[28]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n30),
        .Q(i1[29]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[1]),
        .Q(i1[16]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[2]_i_1__4_n_0 ),
        .Q(i1[17]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[3]_i_1__4_n_0 ),
        .Q(i1[18]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[4]_i_1__4_n_0 ),
        .Q(i1[19]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[5]_i_1__4_n_0 ),
        .Q(i1[20]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[6]_i_1__4_n_0 ),
        .Q(i1[21]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[7]),
        .Q(i1[22]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[9]_i_1__4_n_0 ),
        .Q(i1[23]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[10]_i_1__4 
       (.I0(\n8_reg_n_0_[1] ),
        .I1(n21[1]),
        .I2(n21[0]),
        .I3(\n8_reg_n_0_[0] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(n341_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[11]_i_1__4 
       (.I0(\n37[12]_i_2__4_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .O(n341_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[12]_i_1__4 
       (.I0(\n8_reg_n_0_[3] ),
        .I1(n21[3]),
        .I2(\n37[12]_i_2__4_n_0 ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(n341_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[12]_i_2__4 
       (.I0(\n8_reg_n_0_[0] ),
        .I1(n21[0]),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n37[12]_i_2__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[13]_i_1__4 
       (.I0(\n37[14]_i_2__4_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(n341_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[14]_i_1__4 
       (.I0(\n8_reg_n_0_[5] ),
        .I1(n21[5]),
        .I2(\n37[14]_i_2__4_n_0 ),
        .I3(n21[6]),
        .I4(\n8_reg_n_0_[6] ),
        .O(n341_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[14]_i_2__4 
       (.I0(\n37[12]_i_2__4_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n37[14]_i_2__4_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[15]_i_1__4 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n37[15]_i_2__4_n_0 ),
        .O(n341_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[15]_i_2__4 
       (.I0(\n37[14]_i_2__4_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n37[15]_i_2__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[1]_i_1__4 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .O(n350_out[1]));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[2]_i_1__4 
       (.I0(n10[1]),
        .I1(n29[1]),
        .I2(n29[0]),
        .I3(n10[0]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(n350_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[3]_i_1__4 
       (.I0(\n37[4]_i_2__4_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .O(n350_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[4]_i_1__4 
       (.I0(n10[3]),
        .I1(n29[3]),
        .I2(\n37[4]_i_2__4_n_0 ),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(n350_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[4]_i_2__4 
       (.I0(n10[0]),
        .I1(n29[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n37[4]_i_2__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[5]_i_1__4 
       (.I0(\n37[6]_i_2__4_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(n350_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[6]_i_1__4 
       (.I0(n10[5]),
        .I1(n29[5]),
        .I2(\n37[6]_i_2__4_n_0 ),
        .I3(n29[6]),
        .I4(n10[6]),
        .O(n350_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[6]_i_2__4 
       (.I0(\n37[4]_i_2__4_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n37[6]_i_2__4_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[7]_i_1__4 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n37[7]_i_2__4_n_0 ),
        .O(n350_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[7]_i_2__4 
       (.I0(\n37[6]_i_2__4_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n37[7]_i_2__4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n37[8]_i_1__1 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .O(n341_out[0]));
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[9]_i_1__4 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .O(n341_out[1]));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[2]),
        .Q(i1[9]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[3]),
        .Q(i1[10]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[4]),
        .Q(i1[11]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[5]),
        .Q(i1[12]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[6]),
        .Q(i1[13]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[7]),
        .Q(i1[14]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[1]),
        .Q(i1[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[2]),
        .Q(i1[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[3]),
        .Q(i1[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[4]),
        .Q(i1[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[5]),
        .Q(i1[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[6]),
        .Q(i1[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[7]),
        .Q(i1[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[0]),
        .Q(i1[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[1]),
        .Q(i1[8]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[0]),
        .Q(\n4_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[1]),
        .Q(\n4_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[2]),
        .Q(\n4_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[3]),
        .Q(\n4_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[4]),
        .Q(\n4_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[5]),
        .Q(\n4_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[6]),
        .Q(\n4_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s7_3[7]),
        .Q(\n4_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[0]),
        .Q(\n7_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[1]),
        .Q(\n7_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[2]),
        .Q(\n7_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[3]),
        .Q(\n7_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[4]),
        .Q(\n7_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[5]),
        .Q(\n7_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[6]),
        .Q(\n7_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[7]),
        .Q(\n7_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[0] ),
        .Q(\n8_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[1] ),
        .Q(\n8_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[2] ),
        .Q(\n8_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[3] ),
        .Q(\n8_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[4] ),
        .Q(\n8_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[5] ),
        .Q(\n8_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[6] ),
        .Q(\n8_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[7] ),
        .Q(\n8_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[0] ),
        .Q(\n9_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[1] ),
        .Q(\n9_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[2] ),
        .Q(\n9_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[3] ),
        .Q(\n9_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[4] ),
        .Q(\n9_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[5] ),
        .Q(\n9_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[6] ),
        .Q(\n9_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[7] ),
        .Q(\n9_reg_n_0_[7] ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_11" *) 
module switch_elements_cf_fft_512_8_11
   (\n9_reg[0] ,
    s5_3,
    rst_i,
    enable_i,
    clk_i,
    s6_3,
    D);
  output [15:0]\n9_reg[0] ;
  output [15:0]s5_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]s6_3;
  input [15:0]D;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire [15:0]n33;
  wire [15:1]n37;
  wire n4;
  wire [15:0]\n9_reg[0] ;
  wire rst_i;
  wire s29_n_0;
  wire [15:0]s5_3;
  wire [15:0]s6_3;

  switch_elements_cf_fft_512_8_31_7 s25
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i8(i8),
        .n4(n4),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_12 s26
       (.D(D),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .rst_i(rst_i),
        .s6_3(s6_3));
  switch_elements_cf_fft_512_8_26_8 s28
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .i8(i8),
        .\n1_reg[0] (s29_n_0),
        .n4(n4),
        .\n9_reg[0] (\n9_reg[0] ),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_27_9 s29
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .i8(i8),
        .\n9_reg[0]_0 (s29_n_0),
        .rst_i(rst_i),
        .s5_3(s5_3));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_12" *) 
module switch_elements_cf_fft_512_8_12
   (i1,
    rst_i,
    enable_i,
    clk_i,
    s6_3,
    D);
  output [29:0]i1;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]s6_3;
  input [15:0]D;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [7:0]n10;
  wire [7:0]n15;
  wire \n16[3]_i_10_n_0 ;
  wire \n16[3]_i_11_n_0 ;
  wire \n16[3]_i_12_n_0 ;
  wire \n16[3]_i_13_n_0 ;
  wire \n16[3]_i_14_n_0 ;
  wire \n16[3]_i_15_n_0 ;
  wire \n16[3]_i_16_n_0 ;
  wire \n16[3]_i_18_n_0 ;
  wire \n16[3]_i_19_n_0 ;
  wire \n16[3]_i_20_n_0 ;
  wire \n16[3]_i_21_n_0 ;
  wire \n16[3]_i_22_n_0 ;
  wire \n16[3]_i_23_n_0 ;
  wire \n16[3]_i_24_n_0 ;
  wire \n16[3]_i_25_n_0 ;
  wire \n16[3]_i_26_n_0 ;
  wire \n16[3]_i_27_n_0 ;
  wire \n16[3]_i_28_n_0 ;
  wire \n16[3]_i_2_n_0 ;
  wire \n16[3]_i_3_n_0 ;
  wire \n16[3]_i_4_n_0 ;
  wire \n16[3]_i_5_n_0 ;
  wire \n16[3]_i_6_n_0 ;
  wire \n16[3]_i_7_n_0 ;
  wire \n16[3]_i_8_n_0 ;
  wire \n16[3]_i_9_n_0 ;
  wire \n16[7]_i_13_n_0 ;
  wire \n16[7]_i_14_n_0 ;
  wire \n16[7]_i_15_n_0 ;
  wire \n16[7]_i_16_n_0 ;
  wire \n16[7]_i_17_n_0 ;
  wire \n16[7]_i_18_n_0 ;
  wire \n16[7]_i_19_n_0 ;
  wire \n16[7]_i_20_n_0 ;
  wire \n16[7]_i_21_n_0 ;
  wire \n16[7]_i_22_n_0 ;
  wire \n16[7]_i_23_n_0 ;
  wire \n16[7]_i_24_n_0 ;
  wire \n16[7]_i_25_n_0 ;
  wire \n16[7]_i_26_n_0 ;
  wire \n16[7]_i_27_n_0 ;
  wire \n16[7]_i_28_n_0 ;
  wire \n16[7]_i_29_n_0 ;
  wire \n16[7]_i_2_n_0 ;
  wire \n16[7]_i_30_n_0 ;
  wire \n16[7]_i_31_n_0 ;
  wire \n16[7]_i_32_n_0 ;
  wire \n16[7]_i_33_n_0 ;
  wire \n16[7]_i_34_n_0 ;
  wire \n16[7]_i_35_n_0 ;
  wire \n16[7]_i_36_n_0 ;
  wire \n16[7]_i_37_n_0 ;
  wire \n16[7]_i_38_n_0 ;
  wire \n16[7]_i_3_n_0 ;
  wire \n16[7]_i_4_n_0 ;
  wire \n16[7]_i_5_n_0 ;
  wire \n16[7]_i_6_n_0 ;
  wire \n16[7]_i_7_n_0 ;
  wire \n16[7]_i_8_n_0 ;
  wire \n16_reg[3]_i_17_n_0 ;
  wire \n16_reg[3]_i_17_n_1 ;
  wire \n16_reg[3]_i_17_n_10 ;
  wire \n16_reg[3]_i_17_n_11 ;
  wire \n16_reg[3]_i_17_n_12 ;
  wire \n16_reg[3]_i_17_n_15 ;
  wire \n16_reg[3]_i_17_n_2 ;
  wire \n16_reg[3]_i_17_n_3 ;
  wire \n16_reg[3]_i_17_n_4 ;
  wire \n16_reg[3]_i_17_n_5 ;
  wire \n16_reg[3]_i_17_n_6 ;
  wire \n16_reg[3]_i_17_n_7 ;
  wire \n16_reg[3]_i_17_n_8 ;
  wire \n16_reg[3]_i_17_n_9 ;
  wire \n16_reg[3]_i_1_n_0 ;
  wire \n16_reg[3]_i_1_n_1 ;
  wire \n16_reg[3]_i_1_n_2 ;
  wire \n16_reg[3]_i_1_n_3 ;
  wire \n16_reg[3]_i_1_n_4 ;
  wire \n16_reg[3]_i_1_n_5 ;
  wire \n16_reg[3]_i_1_n_6 ;
  wire \n16_reg[3]_i_1_n_7 ;
  wire \n16_reg[7]_i_10_n_1 ;
  wire \n16_reg[7]_i_10_n_10 ;
  wire \n16_reg[7]_i_10_n_11 ;
  wire \n16_reg[7]_i_10_n_12 ;
  wire \n16_reg[7]_i_10_n_13 ;
  wire \n16_reg[7]_i_10_n_14 ;
  wire \n16_reg[7]_i_10_n_15 ;
  wire \n16_reg[7]_i_10_n_2 ;
  wire \n16_reg[7]_i_10_n_3 ;
  wire \n16_reg[7]_i_10_n_4 ;
  wire \n16_reg[7]_i_10_n_5 ;
  wire \n16_reg[7]_i_10_n_6 ;
  wire \n16_reg[7]_i_10_n_7 ;
  wire \n16_reg[7]_i_10_n_8 ;
  wire \n16_reg[7]_i_10_n_9 ;
  wire \n16_reg[7]_i_11_n_0 ;
  wire \n16_reg[7]_i_11_n_1 ;
  wire \n16_reg[7]_i_11_n_10 ;
  wire \n16_reg[7]_i_11_n_11 ;
  wire \n16_reg[7]_i_11_n_12 ;
  wire \n16_reg[7]_i_11_n_13 ;
  wire \n16_reg[7]_i_11_n_14 ;
  wire \n16_reg[7]_i_11_n_2 ;
  wire \n16_reg[7]_i_11_n_3 ;
  wire \n16_reg[7]_i_11_n_4 ;
  wire \n16_reg[7]_i_11_n_5 ;
  wire \n16_reg[7]_i_11_n_6 ;
  wire \n16_reg[7]_i_11_n_7 ;
  wire \n16_reg[7]_i_11_n_8 ;
  wire \n16_reg[7]_i_11_n_9 ;
  wire \n16_reg[7]_i_12_n_14 ;
  wire \n16_reg[7]_i_12_n_15 ;
  wire \n16_reg[7]_i_12_n_5 ;
  wire \n16_reg[7]_i_12_n_7 ;
  wire \n16_reg[7]_i_1_n_5 ;
  wire \n16_reg[7]_i_1_n_6 ;
  wire \n16_reg[7]_i_1_n_7 ;
  wire \n16_reg[7]_i_9_n_14 ;
  wire \n16_reg[7]_i_9_n_15 ;
  wire \n16_reg[7]_i_9_n_5 ;
  wire \n16_reg[7]_i_9_n_7 ;
  wire \n16_reg_n_0_[0] ;
  wire \n16_reg_n_0_[1] ;
  wire \n16_reg_n_0_[2] ;
  wire \n16_reg_n_0_[3] ;
  wire \n16_reg_n_0_[4] ;
  wire \n16_reg_n_0_[5] ;
  wire \n16_reg_n_0_[6] ;
  wire \n16_reg_n_0_[7] ;
  wire \n1_reg_n_0_[0] ;
  wire \n1_reg_n_0_[1] ;
  wire \n1_reg_n_0_[2] ;
  wire \n1_reg_n_0_[3] ;
  wire \n1_reg_n_0_[4] ;
  wire \n1_reg_n_0_[5] ;
  wire \n1_reg_n_0_[6] ;
  wire \n1_reg_n_0_[7] ;
  wire [7:0]n2;
  wire [7:0]n202_out;
  wire [7:0]n21;
  wire \n21[7]_i_2_n_0 ;
  wire \n21[7]_i_3_n_0 ;
  wire \n21[7]_i_4_n_0 ;
  wire \n21[7]_i_5_n_0 ;
  wire \n21[7]_i_6_n_0 ;
  wire \n21[7]_i_7_n_0 ;
  wire \n21[7]_i_8_n_0 ;
  wire \n21[7]_i_9_n_0 ;
  wire \n21_reg[7]_i_1_n_1 ;
  wire \n21_reg[7]_i_1_n_2 ;
  wire \n21_reg[7]_i_1_n_3 ;
  wire \n21_reg[7]_i_1_n_4 ;
  wire \n21_reg[7]_i_1_n_5 ;
  wire \n21_reg[7]_i_1_n_6 ;
  wire \n21_reg[7]_i_1_n_7 ;
  wire n22__0_n_0;
  wire n22__1_n_0;
  wire n22__2_n_0;
  wire n22__3_n_0;
  wire n22__4_n_0;
  wire n22__5_n_0;
  wire n22__6_n_0;
  wire n22_n_0;
  wire [7:0]n26;
  wire [7:0]n27;
  wire \n27[3]_i_10_n_0 ;
  wire \n27[3]_i_11_n_0 ;
  wire \n27[3]_i_12_n_0 ;
  wire \n27[3]_i_13_n_0 ;
  wire \n27[3]_i_14_n_0 ;
  wire \n27[3]_i_15_n_0 ;
  wire \n27[3]_i_16_n_0 ;
  wire \n27[3]_i_18_n_0 ;
  wire \n27[3]_i_19_n_0 ;
  wire \n27[3]_i_20_n_0 ;
  wire \n27[3]_i_21_n_0 ;
  wire \n27[3]_i_22_n_0 ;
  wire \n27[3]_i_23_n_0 ;
  wire \n27[3]_i_24_n_0 ;
  wire \n27[3]_i_25_n_0 ;
  wire \n27[3]_i_26_n_0 ;
  wire \n27[3]_i_27_n_0 ;
  wire \n27[3]_i_28_n_0 ;
  wire \n27[3]_i_2_n_0 ;
  wire \n27[3]_i_3_n_0 ;
  wire \n27[3]_i_4_n_0 ;
  wire \n27[3]_i_5_n_0 ;
  wire \n27[3]_i_6_n_0 ;
  wire \n27[3]_i_7_n_0 ;
  wire \n27[3]_i_8_n_0 ;
  wire \n27[3]_i_9_n_0 ;
  wire \n27[7]_i_13_n_0 ;
  wire \n27[7]_i_14_n_0 ;
  wire \n27[7]_i_15_n_0 ;
  wire \n27[7]_i_16_n_0 ;
  wire \n27[7]_i_17_n_0 ;
  wire \n27[7]_i_18_n_0 ;
  wire \n27[7]_i_19_n_0 ;
  wire \n27[7]_i_20_n_0 ;
  wire \n27[7]_i_21_n_0 ;
  wire \n27[7]_i_22_n_0 ;
  wire \n27[7]_i_23_n_0 ;
  wire \n27[7]_i_24_n_0 ;
  wire \n27[7]_i_25_n_0 ;
  wire \n27[7]_i_26_n_0 ;
  wire \n27[7]_i_27_n_0 ;
  wire \n27[7]_i_28_n_0 ;
  wire \n27[7]_i_29_n_0 ;
  wire \n27[7]_i_2_n_0 ;
  wire \n27[7]_i_30_n_0 ;
  wire \n27[7]_i_31_n_0 ;
  wire \n27[7]_i_32_n_0 ;
  wire \n27[7]_i_33_n_0 ;
  wire \n27[7]_i_34_n_0 ;
  wire \n27[7]_i_35_n_0 ;
  wire \n27[7]_i_36_n_0 ;
  wire \n27[7]_i_37_n_0 ;
  wire \n27[7]_i_38_n_0 ;
  wire \n27[7]_i_3_n_0 ;
  wire \n27[7]_i_4_n_0 ;
  wire \n27[7]_i_5_n_0 ;
  wire \n27[7]_i_6_n_0 ;
  wire \n27[7]_i_7_n_0 ;
  wire \n27[7]_i_8_n_0 ;
  wire \n27_reg[3]_i_17_n_0 ;
  wire \n27_reg[3]_i_17_n_1 ;
  wire \n27_reg[3]_i_17_n_10 ;
  wire \n27_reg[3]_i_17_n_11 ;
  wire \n27_reg[3]_i_17_n_12 ;
  wire \n27_reg[3]_i_17_n_15 ;
  wire \n27_reg[3]_i_17_n_2 ;
  wire \n27_reg[3]_i_17_n_3 ;
  wire \n27_reg[3]_i_17_n_4 ;
  wire \n27_reg[3]_i_17_n_5 ;
  wire \n27_reg[3]_i_17_n_6 ;
  wire \n27_reg[3]_i_17_n_7 ;
  wire \n27_reg[3]_i_17_n_8 ;
  wire \n27_reg[3]_i_17_n_9 ;
  wire \n27_reg[3]_i_1_n_0 ;
  wire \n27_reg[3]_i_1_n_1 ;
  wire \n27_reg[3]_i_1_n_2 ;
  wire \n27_reg[3]_i_1_n_3 ;
  wire \n27_reg[3]_i_1_n_4 ;
  wire \n27_reg[3]_i_1_n_5 ;
  wire \n27_reg[3]_i_1_n_6 ;
  wire \n27_reg[3]_i_1_n_7 ;
  wire \n27_reg[7]_i_10_n_1 ;
  wire \n27_reg[7]_i_10_n_10 ;
  wire \n27_reg[7]_i_10_n_11 ;
  wire \n27_reg[7]_i_10_n_12 ;
  wire \n27_reg[7]_i_10_n_13 ;
  wire \n27_reg[7]_i_10_n_14 ;
  wire \n27_reg[7]_i_10_n_15 ;
  wire \n27_reg[7]_i_10_n_2 ;
  wire \n27_reg[7]_i_10_n_3 ;
  wire \n27_reg[7]_i_10_n_4 ;
  wire \n27_reg[7]_i_10_n_5 ;
  wire \n27_reg[7]_i_10_n_6 ;
  wire \n27_reg[7]_i_10_n_7 ;
  wire \n27_reg[7]_i_10_n_8 ;
  wire \n27_reg[7]_i_10_n_9 ;
  wire \n27_reg[7]_i_11_n_0 ;
  wire \n27_reg[7]_i_11_n_1 ;
  wire \n27_reg[7]_i_11_n_10 ;
  wire \n27_reg[7]_i_11_n_11 ;
  wire \n27_reg[7]_i_11_n_12 ;
  wire \n27_reg[7]_i_11_n_13 ;
  wire \n27_reg[7]_i_11_n_14 ;
  wire \n27_reg[7]_i_11_n_2 ;
  wire \n27_reg[7]_i_11_n_3 ;
  wire \n27_reg[7]_i_11_n_4 ;
  wire \n27_reg[7]_i_11_n_5 ;
  wire \n27_reg[7]_i_11_n_6 ;
  wire \n27_reg[7]_i_11_n_7 ;
  wire \n27_reg[7]_i_11_n_8 ;
  wire \n27_reg[7]_i_11_n_9 ;
  wire \n27_reg[7]_i_12_n_14 ;
  wire \n27_reg[7]_i_12_n_15 ;
  wire \n27_reg[7]_i_12_n_5 ;
  wire \n27_reg[7]_i_12_n_7 ;
  wire \n27_reg[7]_i_1_n_5 ;
  wire \n27_reg[7]_i_1_n_6 ;
  wire \n27_reg[7]_i_1_n_7 ;
  wire \n27_reg[7]_i_9_n_14 ;
  wire \n27_reg[7]_i_9_n_15 ;
  wire \n27_reg[7]_i_9_n_5 ;
  wire \n27_reg[7]_i_9_n_7 ;
  wire [7:0]n29;
  wire [7:7]n30;
  wire [7:0]n31;
  wire \n33[10]_i_1__3_n_0 ;
  wire \n33[11]_i_1__3_n_0 ;
  wire \n33[12]_i_1__3_n_0 ;
  wire \n33[12]_i_2__3_n_0 ;
  wire \n33[13]_i_1__3_n_0 ;
  wire \n33[14]_i_1__3_n_0 ;
  wire \n33[14]_i_2__3_n_0 ;
  wire \n33[15]_i_2__3_n_0 ;
  wire \n33[2]_i_1__3_n_0 ;
  wire \n33[3]_i_1__3_n_0 ;
  wire \n33[4]_i_1__3_n_0 ;
  wire \n33[4]_i_2__3_n_0 ;
  wire \n33[5]_i_1__3_n_0 ;
  wire \n33[6]_i_1__3_n_0 ;
  wire \n33[6]_i_2__3_n_0 ;
  wire \n33[7]_i_2__3_n_0 ;
  wire \n33[9]_i_1__3_n_0 ;
  wire [7:0]n341_out;
  wire [7:1]n350_out;
  wire \n37[12]_i_2__3_n_0 ;
  wire \n37[14]_i_2__3_n_0 ;
  wire \n37[15]_i_2__3_n_0 ;
  wire \n37[4]_i_2__3_n_0 ;
  wire \n37[6]_i_2__3_n_0 ;
  wire \n37[7]_i_2__3_n_0 ;
  wire \n4_reg_n_0_[0] ;
  wire \n4_reg_n_0_[1] ;
  wire \n4_reg_n_0_[2] ;
  wire \n4_reg_n_0_[3] ;
  wire \n4_reg_n_0_[4] ;
  wire \n4_reg_n_0_[5] ;
  wire \n4_reg_n_0_[6] ;
  wire \n4_reg_n_0_[7] ;
  wire \n7_reg_n_0_[0] ;
  wire \n7_reg_n_0_[1] ;
  wire \n7_reg_n_0_[2] ;
  wire \n7_reg_n_0_[3] ;
  wire \n7_reg_n_0_[4] ;
  wire \n7_reg_n_0_[5] ;
  wire \n7_reg_n_0_[6] ;
  wire \n7_reg_n_0_[7] ;
  wire \n8_reg_n_0_[0] ;
  wire \n8_reg_n_0_[1] ;
  wire \n8_reg_n_0_[2] ;
  wire \n8_reg_n_0_[3] ;
  wire \n8_reg_n_0_[4] ;
  wire \n8_reg_n_0_[5] ;
  wire \n8_reg_n_0_[6] ;
  wire \n8_reg_n_0_[7] ;
  wire \n9_reg_n_0_[0] ;
  wire \n9_reg_n_0_[1] ;
  wire \n9_reg_n_0_[2] ;
  wire \n9_reg_n_0_[3] ;
  wire \n9_reg_n_0_[4] ;
  wire \n9_reg_n_0_[5] ;
  wire \n9_reg_n_0_[6] ;
  wire \n9_reg_n_0_[7] ;
  wire rst_i;
  wire [15:0]s6_3;
  wire [3:0]\NLW_n16_reg[3]_i_1_O_UNCONNECTED ;
  wire [2:1]\NLW_n16_reg[3]_i_17_O_UNCONNECTED ;
  wire [7:3]\NLW_n16_reg[7]_i_1_CO_UNCONNECTED ;
  wire [7:4]\NLW_n16_reg[7]_i_1_O_UNCONNECTED ;
  wire [7:7]\NLW_n16_reg[7]_i_10_CO_UNCONNECTED ;
  wire [0:0]\NLW_n16_reg[7]_i_11_O_UNCONNECTED ;
  wire [7:1]\NLW_n16_reg[7]_i_12_CO_UNCONNECTED ;
  wire [7:2]\NLW_n16_reg[7]_i_12_O_UNCONNECTED ;
  wire [7:1]\NLW_n16_reg[7]_i_9_CO_UNCONNECTED ;
  wire [7:2]\NLW_n16_reg[7]_i_9_O_UNCONNECTED ;
  wire [7:7]\NLW_n21_reg[7]_i_1_CO_UNCONNECTED ;
  wire [3:0]\NLW_n27_reg[3]_i_1_O_UNCONNECTED ;
  wire [2:1]\NLW_n27_reg[3]_i_17_O_UNCONNECTED ;
  wire [7:3]\NLW_n27_reg[7]_i_1_CO_UNCONNECTED ;
  wire [7:4]\NLW_n27_reg[7]_i_1_O_UNCONNECTED ;
  wire [7:7]\NLW_n27_reg[7]_i_10_CO_UNCONNECTED ;
  wire [0:0]\NLW_n27_reg[7]_i_11_O_UNCONNECTED ;
  wire [7:1]\NLW_n27_reg[7]_i_12_CO_UNCONNECTED ;
  wire [7:2]\NLW_n27_reg[7]_i_12_O_UNCONNECTED ;
  wire [7:1]\NLW_n27_reg[7]_i_9_CO_UNCONNECTED ;
  wire [7:2]\NLW_n27_reg[7]_i_9_O_UNCONNECTED ;

  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[0] ),
        .Q(n10[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[1] ),
        .Q(n10[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[2] ),
        .Q(n10[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[3] ),
        .Q(n10[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[4] ),
        .Q(n10[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[5] ),
        .Q(n10[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[6] ),
        .Q(n10[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[7] ),
        .Q(n10[7]),
        .R(rst_i));
  (* HLUTNM = "lutpair47" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_10 
       (.I0(\n16_reg[7]_i_10_n_13 ),
        .I1(\n16_reg[7]_i_11_n_9 ),
        .I2(\n16_reg[7]_i_12_n_14 ),
        .I3(\n16[3]_i_3_n_0 ),
        .O(\n16[3]_i_10_n_0 ));
  (* HLUTNM = "lutpair46" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_11 
       (.I0(\n16_reg[7]_i_10_n_14 ),
        .I1(\n16_reg[7]_i_11_n_10 ),
        .I2(\n16_reg[7]_i_12_n_15 ),
        .I3(\n16[3]_i_4_n_0 ),
        .O(\n16[3]_i_11_n_0 ));
  (* HLUTNM = "lutpair45" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_12 
       (.I0(\n16_reg[7]_i_10_n_15 ),
        .I1(\n16_reg[7]_i_11_n_11 ),
        .I2(\n16_reg[3]_i_17_n_8 ),
        .I3(\n16[3]_i_5_n_0 ),
        .O(\n16[3]_i_12_n_0 ));
  (* HLUTNM = "lutpair44" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_13 
       (.I0(n22__6_n_0),
        .I1(\n16_reg[7]_i_11_n_12 ),
        .I2(\n16_reg[3]_i_17_n_9 ),
        .I3(\n16[3]_i_6_n_0 ),
        .O(\n16[3]_i_13_n_0 ));
  (* HLUTNM = "lutpair95" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n16[3]_i_14 
       (.I0(\n16_reg[7]_i_11_n_13 ),
        .I1(\n16_reg[3]_i_17_n_10 ),
        .I2(\n16_reg[3]_i_17_n_11 ),
        .I3(\n16_reg[7]_i_11_n_14 ),
        .O(\n16[3]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n16[3]_i_15 
       (.I0(\n16_reg[3]_i_17_n_12 ),
        .I1(\n16_reg[3]_i_17_n_15 ),
        .I2(\n16_reg[7]_i_11_n_14 ),
        .I3(\n16_reg[3]_i_17_n_11 ),
        .O(\n16[3]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n16[3]_i_16 
       (.I0(\n16_reg[3]_i_17_n_12 ),
        .I1(\n16_reg[3]_i_17_n_15 ),
        .O(\n16[3]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_18 
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(n22__1_n_0),
        .O(\n16[3]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_19 
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__2_n_0),
        .O(\n16[3]_i_19_n_0 ));
  (* HLUTNM = "lutpair47" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_2 
       (.I0(\n16_reg[7]_i_10_n_13 ),
        .I1(\n16_reg[7]_i_11_n_9 ),
        .I2(\n16_reg[7]_i_12_n_14 ),
        .O(\n16[3]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_20 
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(n22__3_n_0),
        .O(\n16[3]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n16[3]_i_21 
       (.I0(n22__4_n_0),
        .I1(n22__5_n_0),
        .I2(n22__3_n_0),
        .O(\n16[3]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h9669)) 
    \n16[3]_i_22 
       (.I0(\n16[7]_i_23_n_0 ),
        .I1(n22__0_n_0),
        .I2(n22__1_n_0),
        .I3(n22_n_0),
        .O(\n16[3]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[3]_i_23 
       (.I0(n22__3_n_0),
        .I1(n22__1_n_0),
        .I2(n22__2_n_0),
        .I3(n22__0_n_0),
        .O(\n16[3]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[3]_i_24 
       (.I0(n22__4_n_0),
        .I1(n22__2_n_0),
        .I2(n22__3_n_0),
        .I3(n22__1_n_0),
        .O(\n16[3]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[3]_i_25 
       (.I0(n22__5_n_0),
        .I1(n22__3_n_0),
        .I2(n22__4_n_0),
        .I3(n22__2_n_0),
        .O(\n16[3]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h6696)) 
    \n16[3]_i_26 
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__5_n_0),
        .I3(n22__6_n_0),
        .O(\n16[3]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n16[3]_i_27 
       (.I0(n22__6_n_0),
        .I1(n22__5_n_0),
        .I2(n22__4_n_0),
        .O(\n16[3]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n16[3]_i_28 
       (.I0(n22__5_n_0),
        .I1(n22__6_n_0),
        .O(\n16[3]_i_28_n_0 ));
  (* HLUTNM = "lutpair46" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_3 
       (.I0(\n16_reg[7]_i_10_n_14 ),
        .I1(\n16_reg[7]_i_11_n_10 ),
        .I2(\n16_reg[7]_i_12_n_15 ),
        .O(\n16[3]_i_3_n_0 ));
  (* HLUTNM = "lutpair45" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_4 
       (.I0(\n16_reg[7]_i_10_n_15 ),
        .I1(\n16_reg[7]_i_11_n_11 ),
        .I2(\n16_reg[3]_i_17_n_8 ),
        .O(\n16[3]_i_4_n_0 ));
  (* HLUTNM = "lutpair44" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_5 
       (.I0(n22__6_n_0),
        .I1(\n16_reg[7]_i_11_n_12 ),
        .I2(\n16_reg[3]_i_17_n_9 ),
        .O(\n16[3]_i_5_n_0 ));
  (* HLUTNM = "lutpair95" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \n16[3]_i_6 
       (.I0(\n16_reg[7]_i_11_n_13 ),
        .I1(\n16_reg[3]_i_17_n_10 ),
        .O(\n16[3]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n16[3]_i_7 
       (.I0(\n16_reg[3]_i_17_n_11 ),
        .I1(\n16_reg[7]_i_11_n_14 ),
        .O(\n16[3]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n16[3]_i_8 
       (.I0(\n16_reg[3]_i_17_n_12 ),
        .I1(\n16_reg[3]_i_17_n_15 ),
        .O(\n16[3]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_9 
       (.I0(\n16[3]_i_2_n_0 ),
        .I1(\n16_reg[7]_i_11_n_8 ),
        .I2(\n16_reg[7]_i_10_n_12 ),
        .I3(\n16_reg[7]_i_12_n_5 ),
        .O(\n16[3]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \n16[7]_i_13 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \n16[7]_i_14 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(\n16[7]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \n16[7]_i_15 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h4D)) 
    \n16[7]_i_16 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(\n16[7]_i_16_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n16[7]_i_17 
       (.I0(n22_n_0),
        .O(\n16[7]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n16[7]_i_18 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n16[7]_i_19 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .O(\n16[7]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n16[7]_i_2 
       (.I0(\n16_reg[7]_i_9_n_14 ),
        .I1(\n16_reg[7]_i_10_n_10 ),
        .O(\n16[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n16[7]_i_20 
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .O(\n16[7]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n16[7]_i_21 
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .O(\n16[7]_i_21_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n16[7]_i_22 
       (.I0(n22__5_n_0),
        .O(\n16[7]_i_22_n_0 ));
  (* HLUTNM = "lutpair94" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_23 
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .O(\n16[7]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_24 
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(n22__1_n_0),
        .O(\n16[7]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_25 
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__2_n_0),
        .O(\n16[7]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_26 
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(n22__3_n_0),
        .O(\n16[7]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n16[7]_i_27 
       (.I0(n22__4_n_0),
        .I1(n22__5_n_0),
        .I2(n22__3_n_0),
        .O(\n16[7]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h9669)) 
    \n16[7]_i_28 
       (.I0(\n16[7]_i_23_n_0 ),
        .I1(n22__0_n_0),
        .I2(n22__1_n_0),
        .I3(n22_n_0),
        .O(\n16[7]_i_28_n_0 ));
  (* HLUTNM = "lutpair94" *) 
  LUT4 #(
    .INIT(16'h781E)) 
    \n16[7]_i_29 
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(n22__3_n_0),
        .O(\n16[7]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n16[7]_i_3 
       (.I0(\n16_reg[7]_i_9_n_15 ),
        .I1(\n16_reg[7]_i_10_n_11 ),
        .O(\n16[7]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[7]_i_30 
       (.I0(n22__4_n_0),
        .I1(n22__2_n_0),
        .I2(n22__3_n_0),
        .I3(n22__1_n_0),
        .O(\n16[7]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[7]_i_31 
       (.I0(n22__5_n_0),
        .I1(n22__3_n_0),
        .I2(n22__4_n_0),
        .I3(n22__2_n_0),
        .O(\n16[7]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h6696)) 
    \n16[7]_i_32 
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__5_n_0),
        .I3(n22__6_n_0),
        .O(\n16[7]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n16[7]_i_33 
       (.I0(n22__6_n_0),
        .I1(n22__5_n_0),
        .I2(n22__4_n_0),
        .O(\n16[7]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n16[7]_i_34 
       (.I0(n22__5_n_0),
        .I1(n22__6_n_0),
        .O(\n16[7]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \n16[7]_i_35 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \n16[7]_i_36 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(\n16[7]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \n16[7]_i_37 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h4D)) 
    \n16[7]_i_38 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(\n16[7]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_4 
       (.I0(\n16_reg[7]_i_10_n_12 ),
        .I1(\n16_reg[7]_i_11_n_8 ),
        .I2(\n16_reg[7]_i_12_n_5 ),
        .O(\n16[7]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \n16[7]_i_5 
       (.I0(\n16_reg[7]_i_9_n_5 ),
        .I1(\n16_reg[7]_i_10_n_9 ),
        .I2(\n16_reg[7]_i_10_n_8 ),
        .O(\n16[7]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n16[7]_i_6 
       (.I0(\n16_reg[7]_i_9_n_14 ),
        .I1(\n16_reg[7]_i_10_n_10 ),
        .I2(\n16_reg[7]_i_10_n_9 ),
        .I3(\n16_reg[7]_i_9_n_5 ),
        .O(\n16[7]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n16[7]_i_7 
       (.I0(\n16_reg[7]_i_9_n_15 ),
        .I1(\n16_reg[7]_i_10_n_11 ),
        .I2(\n16_reg[7]_i_10_n_10 ),
        .I3(\n16_reg[7]_i_9_n_14 ),
        .O(\n16[7]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    \n16[7]_i_8 
       (.I0(\n16_reg[7]_i_12_n_5 ),
        .I1(\n16_reg[7]_i_11_n_8 ),
        .I2(\n16_reg[7]_i_10_n_12 ),
        .I3(\n16_reg[7]_i_10_n_11 ),
        .I4(\n16_reg[7]_i_9_n_15 ),
        .O(\n16[7]_i_8_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[0]),
        .Q(\n16_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[1]),
        .Q(\n16_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[2]),
        .Q(\n16_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[3]),
        .Q(\n16_reg_n_0_[3] ),
        .R(rst_i));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[3]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n16_reg[3]_i_1_n_0 ,\n16_reg[3]_i_1_n_1 ,\n16_reg[3]_i_1_n_2 ,\n16_reg[3]_i_1_n_3 ,\n16_reg[3]_i_1_n_4 ,\n16_reg[3]_i_1_n_5 ,\n16_reg[3]_i_1_n_6 ,\n16_reg[3]_i_1_n_7 }),
        .DI({\n16[3]_i_2_n_0 ,\n16[3]_i_3_n_0 ,\n16[3]_i_4_n_0 ,\n16[3]_i_5_n_0 ,\n16[3]_i_6_n_0 ,\n16[3]_i_7_n_0 ,\n16[3]_i_8_n_0 ,1'b0}),
        .O({n15[3:0],\NLW_n16_reg[3]_i_1_O_UNCONNECTED [3:0]}),
        .S({\n16[3]_i_9_n_0 ,\n16[3]_i_10_n_0 ,\n16[3]_i_11_n_0 ,\n16[3]_i_12_n_0 ,\n16[3]_i_13_n_0 ,\n16[3]_i_14_n_0 ,\n16[3]_i_15_n_0 ,\n16[3]_i_16_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[3]_i_17 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n16_reg[3]_i_17_n_0 ,\n16_reg[3]_i_17_n_1 ,\n16_reg[3]_i_17_n_2 ,\n16_reg[3]_i_17_n_3 ,\n16_reg[3]_i_17_n_4 ,\n16_reg[3]_i_17_n_5 ,\n16_reg[3]_i_17_n_6 ,\n16_reg[3]_i_17_n_7 }),
        .DI({\n16[7]_i_23_n_0 ,\n16[3]_i_18_n_0 ,\n16[3]_i_19_n_0 ,\n16[3]_i_20_n_0 ,\n16[3]_i_21_n_0 ,n22__4_n_0,n22__5_n_0,1'b0}),
        .O({\n16_reg[3]_i_17_n_8 ,\n16_reg[3]_i_17_n_9 ,\n16_reg[3]_i_17_n_10 ,\n16_reg[3]_i_17_n_11 ,\n16_reg[3]_i_17_n_12 ,\NLW_n16_reg[3]_i_17_O_UNCONNECTED [2:1],\n16_reg[3]_i_17_n_15 }),
        .S({\n16[3]_i_22_n_0 ,\n16[3]_i_23_n_0 ,\n16[3]_i_24_n_0 ,\n16[3]_i_25_n_0 ,\n16[3]_i_26_n_0 ,\n16[3]_i_27_n_0 ,\n16[3]_i_28_n_0 ,n22__6_n_0}));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[4]),
        .Q(\n16_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[5]),
        .Q(\n16_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[6]),
        .Q(\n16_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[7]),
        .Q(\n16_reg_n_0_[7] ),
        .R(rst_i));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_1 
       (.CI(\n16_reg[3]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n16_reg[7]_i_1_CO_UNCONNECTED [7:3],\n16_reg[7]_i_1_n_5 ,\n16_reg[7]_i_1_n_6 ,\n16_reg[7]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,\n16[7]_i_2_n_0 ,\n16[7]_i_3_n_0 ,\n16[7]_i_4_n_0 }),
        .O({\NLW_n16_reg[7]_i_1_O_UNCONNECTED [7:4],n15[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,\n16[7]_i_5_n_0 ,\n16[7]_i_6_n_0 ,\n16[7]_i_7_n_0 ,\n16[7]_i_8_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_10 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\NLW_n16_reg[7]_i_10_CO_UNCONNECTED [7],\n16_reg[7]_i_10_n_1 ,\n16_reg[7]_i_10_n_2 ,\n16_reg[7]_i_10_n_3 ,\n16_reg[7]_i_10_n_4 ,\n16_reg[7]_i_10_n_5 ,\n16_reg[7]_i_10_n_6 ,\n16_reg[7]_i_10_n_7 }),
        .DI({1'b0,n22__0_n_0,n22__1_n_0,n22__2_n_0,n22__3_n_0,1'b1,1'b0,1'b1}),
        .O({\n16_reg[7]_i_10_n_8 ,\n16_reg[7]_i_10_n_9 ,\n16_reg[7]_i_10_n_10 ,\n16_reg[7]_i_10_n_11 ,\n16_reg[7]_i_10_n_12 ,\n16_reg[7]_i_10_n_13 ,\n16_reg[7]_i_10_n_14 ,\n16_reg[7]_i_10_n_15 }),
        .S({\n16[7]_i_17_n_0 ,\n16[7]_i_18_n_0 ,\n16[7]_i_19_n_0 ,\n16[7]_i_20_n_0 ,\n16[7]_i_21_n_0 ,n22__3_n_0,n22__4_n_0,\n16[7]_i_22_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_11 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n16_reg[7]_i_11_n_0 ,\n16_reg[7]_i_11_n_1 ,\n16_reg[7]_i_11_n_2 ,\n16_reg[7]_i_11_n_3 ,\n16_reg[7]_i_11_n_4 ,\n16_reg[7]_i_11_n_5 ,\n16_reg[7]_i_11_n_6 ,\n16_reg[7]_i_11_n_7 }),
        .DI({\n16[7]_i_23_n_0 ,\n16[7]_i_24_n_0 ,\n16[7]_i_25_n_0 ,\n16[7]_i_26_n_0 ,\n16[7]_i_27_n_0 ,n22__4_n_0,n22__5_n_0,1'b0}),
        .O({\n16_reg[7]_i_11_n_8 ,\n16_reg[7]_i_11_n_9 ,\n16_reg[7]_i_11_n_10 ,\n16_reg[7]_i_11_n_11 ,\n16_reg[7]_i_11_n_12 ,\n16_reg[7]_i_11_n_13 ,\n16_reg[7]_i_11_n_14 ,\NLW_n16_reg[7]_i_11_O_UNCONNECTED [0]}),
        .S({\n16[7]_i_28_n_0 ,\n16[7]_i_29_n_0 ,\n16[7]_i_30_n_0 ,\n16[7]_i_31_n_0 ,\n16[7]_i_32_n_0 ,\n16[7]_i_33_n_0 ,\n16[7]_i_34_n_0 ,n22__6_n_0}));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_12 
       (.CI(\n16_reg[3]_i_17_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n16_reg[7]_i_12_CO_UNCONNECTED [7:3],\n16_reg[7]_i_12_n_5 ,\NLW_n16_reg[7]_i_12_CO_UNCONNECTED [1],\n16_reg[7]_i_12_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\n16[7]_i_35_n_0 ,\n16[7]_i_36_n_0 }),
        .O({\NLW_n16_reg[7]_i_12_O_UNCONNECTED [7:2],\n16_reg[7]_i_12_n_14 ,\n16_reg[7]_i_12_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,\n16[7]_i_37_n_0 ,\n16[7]_i_38_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_9 
       (.CI(\n16_reg[7]_i_11_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n16_reg[7]_i_9_CO_UNCONNECTED [7:3],\n16_reg[7]_i_9_n_5 ,\NLW_n16_reg[7]_i_9_CO_UNCONNECTED [1],\n16_reg[7]_i_9_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\n16[7]_i_13_n_0 ,\n16[7]_i_14_n_0 }),
        .O({\NLW_n16_reg[7]_i_9_O_UNCONNECTED [7:2],\n16_reg[7]_i_9_n_14 ,\n16_reg[7]_i_9_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,\n16[7]_i_15_n_0 ,\n16[7]_i_16_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[0]),
        .Q(\n1_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[10]),
        .Q(n2[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[11]),
        .Q(n2[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[12]),
        .Q(n2[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[13]),
        .Q(n2[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[14]),
        .Q(n2[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[15]),
        .Q(n2[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[1]),
        .Q(\n1_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[2]),
        .Q(\n1_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[3]),
        .Q(\n1_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[4]),
        .Q(\n1_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[5]),
        .Q(\n1_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[6]),
        .Q(\n1_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[7]),
        .Q(\n1_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[8]),
        .Q(n2[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[9]),
        .Q(n2[1]),
        .R(rst_i));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_2 
       (.I0(\n16_reg_n_0_[7] ),
        .O(\n21[7]_i_2_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_3 
       (.I0(\n16_reg_n_0_[6] ),
        .O(\n21[7]_i_3_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_4 
       (.I0(\n16_reg_n_0_[5] ),
        .O(\n21[7]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_5 
       (.I0(\n16_reg_n_0_[4] ),
        .O(\n21[7]_i_5_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_6 
       (.I0(\n16_reg_n_0_[3] ),
        .O(\n21[7]_i_6_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_7 
       (.I0(\n16_reg_n_0_[2] ),
        .O(\n21[7]_i_7_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_8 
       (.I0(\n16_reg_n_0_[1] ),
        .O(\n21[7]_i_8_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_9 
       (.I0(\n16_reg_n_0_[0] ),
        .O(\n21[7]_i_9_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[0]),
        .Q(n21[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[1]),
        .Q(n21[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[2]),
        .Q(n21[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[3]),
        .Q(n21[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[4]),
        .Q(n21[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[5]),
        .Q(n21[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[6]),
        .Q(n21[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[7]),
        .Q(n21[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n21_reg[7]_i_1 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\NLW_n21_reg[7]_i_1_CO_UNCONNECTED [7],\n21_reg[7]_i_1_n_1 ,\n21_reg[7]_i_1_n_2 ,\n21_reg[7]_i_1_n_3 ,\n21_reg[7]_i_1_n_4 ,\n21_reg[7]_i_1_n_5 ,\n21_reg[7]_i_1_n_6 ,\n21_reg[7]_i_1_n_7 }),
        .DI({1'b0,\n16_reg_n_0_[6] ,\n16_reg_n_0_[5] ,\n16_reg_n_0_[4] ,\n16_reg_n_0_[3] ,\n16_reg_n_0_[2] ,\n16_reg_n_0_[1] ,\n16_reg_n_0_[0] }),
        .O(n202_out),
        .S({\n21[7]_i_2_n_0 ,\n21[7]_i_3_n_0 ,\n21[7]_i_4_n_0 ,\n21[7]_i_5_n_0 ,\n21[7]_i_6_n_0 ,\n21[7]_i_7_n_0 ,\n21[7]_i_8_n_0 ,\n21[7]_i_9_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    n22
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[15]),
        .Q(n22_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__0
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[14]),
        .Q(n22__0_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__1
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[13]),
        .Q(n22__1_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__2
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[12]),
        .Q(n22__2_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__3
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[11]),
        .Q(n22__3_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__4
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[10]),
        .Q(n22__4_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__5
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[9]),
        .Q(n22__5_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__6
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[8]),
        .Q(n22__6_n_0),
        .R(rst_i));
  (* HLUTNM = "lutpair43" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_10 
       (.I0(\n27_reg[7]_i_10_n_13 ),
        .I1(\n27_reg[7]_i_11_n_9 ),
        .I2(\n27_reg[7]_i_12_n_14 ),
        .I3(\n27[3]_i_3_n_0 ),
        .O(\n27[3]_i_10_n_0 ));
  (* HLUTNM = "lutpair42" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_11 
       (.I0(\n27_reg[7]_i_10_n_14 ),
        .I1(\n27_reg[7]_i_11_n_10 ),
        .I2(\n27_reg[7]_i_12_n_15 ),
        .I3(\n27[3]_i_4_n_0 ),
        .O(\n27[3]_i_11_n_0 ));
  (* HLUTNM = "lutpair41" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_12 
       (.I0(\n27_reg[7]_i_10_n_15 ),
        .I1(\n27_reg[7]_i_11_n_11 ),
        .I2(\n27_reg[3]_i_17_n_8 ),
        .I3(\n27[3]_i_5_n_0 ),
        .O(\n27[3]_i_12_n_0 ));
  (* HLUTNM = "lutpair40" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_13 
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n27_reg[7]_i_11_n_12 ),
        .I2(\n27_reg[3]_i_17_n_9 ),
        .I3(\n27[3]_i_6_n_0 ),
        .O(\n27[3]_i_13_n_0 ));
  (* HLUTNM = "lutpair93" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n27[3]_i_14 
       (.I0(\n27_reg[7]_i_11_n_13 ),
        .I1(\n27_reg[3]_i_17_n_10 ),
        .I2(\n27_reg[3]_i_17_n_11 ),
        .I3(\n27_reg[7]_i_11_n_14 ),
        .O(\n27[3]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n27[3]_i_15 
       (.I0(\n27_reg[3]_i_17_n_12 ),
        .I1(\n27_reg[3]_i_17_n_15 ),
        .I2(\n27_reg[7]_i_11_n_14 ),
        .I3(\n27_reg[3]_i_17_n_11 ),
        .O(\n27[3]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n27[3]_i_16 
       (.I0(\n27_reg[3]_i_17_n_12 ),
        .I1(\n27_reg[3]_i_17_n_15 ),
        .O(\n27[3]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_18 
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[5] ),
        .O(\n27[3]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_19 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[4] ),
        .O(\n27[3]_i_19_n_0 ));
  (* HLUTNM = "lutpair43" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_2 
       (.I0(\n27_reg[7]_i_10_n_13 ),
        .I1(\n27_reg[7]_i_11_n_9 ),
        .I2(\n27_reg[7]_i_12_n_14 ),
        .O(\n27[3]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_20 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[2] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(\n27[3]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n27[3]_i_21 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(\n27[3]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h9669)) 
    \n27[3]_i_22 
       (.I0(\n27[7]_i_23_n_0 ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[5] ),
        .I3(\n4_reg_n_0_[7] ),
        .O(\n27[3]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[3]_i_23 
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[5] ),
        .I2(\n4_reg_n_0_[4] ),
        .I3(\n4_reg_n_0_[6] ),
        .O(\n27[3]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[3]_i_24 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[3] ),
        .I3(\n4_reg_n_0_[5] ),
        .O(\n27[3]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[3]_i_25 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[2] ),
        .I3(\n4_reg_n_0_[4] ),
        .O(\n27[3]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h6696)) 
    \n27[3]_i_26 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[1] ),
        .I3(\n4_reg_n_0_[0] ),
        .O(\n27[3]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n27[3]_i_27 
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[2] ),
        .O(\n27[3]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n27[3]_i_28 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[0] ),
        .O(\n27[3]_i_28_n_0 ));
  (* HLUTNM = "lutpair42" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_3 
       (.I0(\n27_reg[7]_i_10_n_14 ),
        .I1(\n27_reg[7]_i_11_n_10 ),
        .I2(\n27_reg[7]_i_12_n_15 ),
        .O(\n27[3]_i_3_n_0 ));
  (* HLUTNM = "lutpair41" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_4 
       (.I0(\n27_reg[7]_i_10_n_15 ),
        .I1(\n27_reg[7]_i_11_n_11 ),
        .I2(\n27_reg[3]_i_17_n_8 ),
        .O(\n27[3]_i_4_n_0 ));
  (* HLUTNM = "lutpair40" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_5 
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n27_reg[7]_i_11_n_12 ),
        .I2(\n27_reg[3]_i_17_n_9 ),
        .O(\n27[3]_i_5_n_0 ));
  (* HLUTNM = "lutpair93" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \n27[3]_i_6 
       (.I0(\n27_reg[7]_i_11_n_13 ),
        .I1(\n27_reg[3]_i_17_n_10 ),
        .O(\n27[3]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n27[3]_i_7 
       (.I0(\n27_reg[3]_i_17_n_11 ),
        .I1(\n27_reg[7]_i_11_n_14 ),
        .O(\n27[3]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n27[3]_i_8 
       (.I0(\n27_reg[3]_i_17_n_12 ),
        .I1(\n27_reg[3]_i_17_n_15 ),
        .O(\n27[3]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_9 
       (.I0(\n27[3]_i_2_n_0 ),
        .I1(\n27_reg[7]_i_11_n_8 ),
        .I2(\n27_reg[7]_i_10_n_12 ),
        .I3(\n27_reg[7]_i_12_n_5 ),
        .O(\n27[3]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \n27[7]_i_13 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \n27[7]_i_14 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \n27[7]_i_15 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h4D)) 
    \n27[7]_i_16 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_16_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n27[7]_i_17 
       (.I0(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n27[7]_i_18 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n27[7]_i_19 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .O(\n27[7]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n27[7]_i_2 
       (.I0(\n27_reg[7]_i_9_n_14 ),
        .I1(\n27_reg[7]_i_10_n_10 ),
        .O(\n27[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n27[7]_i_20 
       (.I0(\n4_reg_n_0_[4] ),
        .I1(\n4_reg_n_0_[5] ),
        .O(\n27[7]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n27[7]_i_21 
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[4] ),
        .O(\n27[7]_i_21_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n27[7]_i_22 
       (.I0(\n4_reg_n_0_[1] ),
        .O(\n27[7]_i_22_n_0 ));
  (* HLUTNM = "lutpair92" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_23 
       (.I0(\n4_reg_n_0_[4] ),
        .I1(\n4_reg_n_0_[5] ),
        .I2(\n4_reg_n_0_[6] ),
        .O(\n27[7]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_24 
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[5] ),
        .O(\n27[7]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_25 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[4] ),
        .O(\n27[7]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_26 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[2] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(\n27[7]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n27[7]_i_27 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(\n27[7]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h9669)) 
    \n27[7]_i_28 
       (.I0(\n27[7]_i_23_n_0 ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[5] ),
        .I3(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_28_n_0 ));
  (* HLUTNM = "lutpair92" *) 
  LUT4 #(
    .INIT(16'h781E)) 
    \n27[7]_i_29 
       (.I0(\n4_reg_n_0_[4] ),
        .I1(\n4_reg_n_0_[5] ),
        .I2(\n4_reg_n_0_[6] ),
        .I3(\n4_reg_n_0_[3] ),
        .O(\n27[7]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n27[7]_i_3 
       (.I0(\n27_reg[7]_i_9_n_15 ),
        .I1(\n27_reg[7]_i_10_n_11 ),
        .O(\n27[7]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[7]_i_30 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[3] ),
        .I3(\n4_reg_n_0_[5] ),
        .O(\n27[7]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[7]_i_31 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[2] ),
        .I3(\n4_reg_n_0_[4] ),
        .O(\n27[7]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h6696)) 
    \n27[7]_i_32 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[1] ),
        .I3(\n4_reg_n_0_[0] ),
        .O(\n27[7]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n27[7]_i_33 
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[2] ),
        .O(\n27[7]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n27[7]_i_34 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[0] ),
        .O(\n27[7]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \n27[7]_i_35 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \n27[7]_i_36 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \n27[7]_i_37 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h4D)) 
    \n27[7]_i_38 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_4 
       (.I0(\n27_reg[7]_i_10_n_12 ),
        .I1(\n27_reg[7]_i_11_n_8 ),
        .I2(\n27_reg[7]_i_12_n_5 ),
        .O(\n27[7]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \n27[7]_i_5 
       (.I0(\n27_reg[7]_i_9_n_5 ),
        .I1(\n27_reg[7]_i_10_n_9 ),
        .I2(\n27_reg[7]_i_10_n_8 ),
        .O(\n27[7]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n27[7]_i_6 
       (.I0(\n27_reg[7]_i_9_n_14 ),
        .I1(\n27_reg[7]_i_10_n_10 ),
        .I2(\n27_reg[7]_i_10_n_9 ),
        .I3(\n27_reg[7]_i_9_n_5 ),
        .O(\n27[7]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n27[7]_i_7 
       (.I0(\n27_reg[7]_i_9_n_15 ),
        .I1(\n27_reg[7]_i_10_n_11 ),
        .I2(\n27_reg[7]_i_10_n_10 ),
        .I3(\n27_reg[7]_i_9_n_14 ),
        .O(\n27[7]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    \n27[7]_i_8 
       (.I0(\n27_reg[7]_i_12_n_5 ),
        .I1(\n27_reg[7]_i_11_n_8 ),
        .I2(\n27_reg[7]_i_10_n_12 ),
        .I3(\n27_reg[7]_i_10_n_11 ),
        .I4(\n27_reg[7]_i_9_n_15 ),
        .O(\n27[7]_i_8_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[0]),
        .Q(n27[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[1]),
        .Q(n27[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[2]),
        .Q(n27[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[3]),
        .Q(n27[3]),
        .R(rst_i));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[3]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n27_reg[3]_i_1_n_0 ,\n27_reg[3]_i_1_n_1 ,\n27_reg[3]_i_1_n_2 ,\n27_reg[3]_i_1_n_3 ,\n27_reg[3]_i_1_n_4 ,\n27_reg[3]_i_1_n_5 ,\n27_reg[3]_i_1_n_6 ,\n27_reg[3]_i_1_n_7 }),
        .DI({\n27[3]_i_2_n_0 ,\n27[3]_i_3_n_0 ,\n27[3]_i_4_n_0 ,\n27[3]_i_5_n_0 ,\n27[3]_i_6_n_0 ,\n27[3]_i_7_n_0 ,\n27[3]_i_8_n_0 ,1'b0}),
        .O({n26[3:0],\NLW_n27_reg[3]_i_1_O_UNCONNECTED [3:0]}),
        .S({\n27[3]_i_9_n_0 ,\n27[3]_i_10_n_0 ,\n27[3]_i_11_n_0 ,\n27[3]_i_12_n_0 ,\n27[3]_i_13_n_0 ,\n27[3]_i_14_n_0 ,\n27[3]_i_15_n_0 ,\n27[3]_i_16_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[3]_i_17 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n27_reg[3]_i_17_n_0 ,\n27_reg[3]_i_17_n_1 ,\n27_reg[3]_i_17_n_2 ,\n27_reg[3]_i_17_n_3 ,\n27_reg[3]_i_17_n_4 ,\n27_reg[3]_i_17_n_5 ,\n27_reg[3]_i_17_n_6 ,\n27_reg[3]_i_17_n_7 }),
        .DI({\n27[7]_i_23_n_0 ,\n27[3]_i_18_n_0 ,\n27[3]_i_19_n_0 ,\n27[3]_i_20_n_0 ,\n27[3]_i_21_n_0 ,\n4_reg_n_0_[2] ,\n4_reg_n_0_[1] ,1'b0}),
        .O({\n27_reg[3]_i_17_n_8 ,\n27_reg[3]_i_17_n_9 ,\n27_reg[3]_i_17_n_10 ,\n27_reg[3]_i_17_n_11 ,\n27_reg[3]_i_17_n_12 ,\NLW_n27_reg[3]_i_17_O_UNCONNECTED [2:1],\n27_reg[3]_i_17_n_15 }),
        .S({\n27[3]_i_22_n_0 ,\n27[3]_i_23_n_0 ,\n27[3]_i_24_n_0 ,\n27[3]_i_25_n_0 ,\n27[3]_i_26_n_0 ,\n27[3]_i_27_n_0 ,\n27[3]_i_28_n_0 ,\n4_reg_n_0_[0] }));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[4]),
        .Q(n27[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[5]),
        .Q(n27[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[6]),
        .Q(n27[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[7]),
        .Q(n27[7]),
        .R(rst_i));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_1 
       (.CI(\n27_reg[3]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n27_reg[7]_i_1_CO_UNCONNECTED [7:3],\n27_reg[7]_i_1_n_5 ,\n27_reg[7]_i_1_n_6 ,\n27_reg[7]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,\n27[7]_i_2_n_0 ,\n27[7]_i_3_n_0 ,\n27[7]_i_4_n_0 }),
        .O({\NLW_n27_reg[7]_i_1_O_UNCONNECTED [7:4],n26[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,\n27[7]_i_5_n_0 ,\n27[7]_i_6_n_0 ,\n27[7]_i_7_n_0 ,\n27[7]_i_8_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_10 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\NLW_n27_reg[7]_i_10_CO_UNCONNECTED [7],\n27_reg[7]_i_10_n_1 ,\n27_reg[7]_i_10_n_2 ,\n27_reg[7]_i_10_n_3 ,\n27_reg[7]_i_10_n_4 ,\n27_reg[7]_i_10_n_5 ,\n27_reg[7]_i_10_n_6 ,\n27_reg[7]_i_10_n_7 }),
        .DI({1'b0,\n4_reg_n_0_[6] ,\n4_reg_n_0_[5] ,\n4_reg_n_0_[4] ,\n4_reg_n_0_[3] ,1'b1,1'b0,1'b1}),
        .O({\n27_reg[7]_i_10_n_8 ,\n27_reg[7]_i_10_n_9 ,\n27_reg[7]_i_10_n_10 ,\n27_reg[7]_i_10_n_11 ,\n27_reg[7]_i_10_n_12 ,\n27_reg[7]_i_10_n_13 ,\n27_reg[7]_i_10_n_14 ,\n27_reg[7]_i_10_n_15 }),
        .S({\n27[7]_i_17_n_0 ,\n27[7]_i_18_n_0 ,\n27[7]_i_19_n_0 ,\n27[7]_i_20_n_0 ,\n27[7]_i_21_n_0 ,\n4_reg_n_0_[3] ,\n4_reg_n_0_[2] ,\n27[7]_i_22_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_11 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n27_reg[7]_i_11_n_0 ,\n27_reg[7]_i_11_n_1 ,\n27_reg[7]_i_11_n_2 ,\n27_reg[7]_i_11_n_3 ,\n27_reg[7]_i_11_n_4 ,\n27_reg[7]_i_11_n_5 ,\n27_reg[7]_i_11_n_6 ,\n27_reg[7]_i_11_n_7 }),
        .DI({\n27[7]_i_23_n_0 ,\n27[7]_i_24_n_0 ,\n27[7]_i_25_n_0 ,\n27[7]_i_26_n_0 ,\n27[7]_i_27_n_0 ,\n4_reg_n_0_[2] ,\n4_reg_n_0_[1] ,1'b0}),
        .O({\n27_reg[7]_i_11_n_8 ,\n27_reg[7]_i_11_n_9 ,\n27_reg[7]_i_11_n_10 ,\n27_reg[7]_i_11_n_11 ,\n27_reg[7]_i_11_n_12 ,\n27_reg[7]_i_11_n_13 ,\n27_reg[7]_i_11_n_14 ,\NLW_n27_reg[7]_i_11_O_UNCONNECTED [0]}),
        .S({\n27[7]_i_28_n_0 ,\n27[7]_i_29_n_0 ,\n27[7]_i_30_n_0 ,\n27[7]_i_31_n_0 ,\n27[7]_i_32_n_0 ,\n27[7]_i_33_n_0 ,\n27[7]_i_34_n_0 ,\n4_reg_n_0_[0] }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_12 
       (.CI(\n27_reg[3]_i_17_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n27_reg[7]_i_12_CO_UNCONNECTED [7:3],\n27_reg[7]_i_12_n_5 ,\NLW_n27_reg[7]_i_12_CO_UNCONNECTED [1],\n27_reg[7]_i_12_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\n27[7]_i_35_n_0 ,\n27[7]_i_36_n_0 }),
        .O({\NLW_n27_reg[7]_i_12_O_UNCONNECTED [7:2],\n27_reg[7]_i_12_n_14 ,\n27_reg[7]_i_12_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,\n27[7]_i_37_n_0 ,\n27[7]_i_38_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_9 
       (.CI(\n27_reg[7]_i_11_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n27_reg[7]_i_9_CO_UNCONNECTED [7:3],\n27_reg[7]_i_9_n_5 ,\NLW_n27_reg[7]_i_9_CO_UNCONNECTED [1],\n27_reg[7]_i_9_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\n27[7]_i_13_n_0 ,\n27[7]_i_14_n_0 }),
        .O({\NLW_n27_reg[7]_i_9_O_UNCONNECTED [7:2],\n27_reg[7]_i_9_n_14 ,\n27_reg[7]_i_9_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,\n27[7]_i_15_n_0 ,\n27[7]_i_16_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[0]),
        .Q(n29[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[1]),
        .Q(n29[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[2]),
        .Q(n29[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[3]),
        .Q(n29[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[4]),
        .Q(n29[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[5]),
        .Q(n29[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[6]),
        .Q(n29[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[7]),
        .Q(n29[7]),
        .R(rst_i));
  LUT2 #(
    .INIT(4'h6)) 
    \n33[0]_i_1__3 
       (.I0(n29[0]),
        .I1(n10[0]),
        .O(n31[0]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[10]_i_1__3 
       (.I0(n21[2]),
        .I1(\n8_reg_n_0_[2] ),
        .I2(\n8_reg_n_0_[1] ),
        .I3(n21[1]),
        .I4(\n8_reg_n_0_[0] ),
        .I5(n21[0]),
        .O(\n33[10]_i_1__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[11]_i_1__3 
       (.I0(n21[3]),
        .I1(\n8_reg_n_0_[3] ),
        .I2(\n33[12]_i_2__3_n_0 ),
        .O(\n33[11]_i_1__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[12]_i_1__3 
       (.I0(n21[4]),
        .I1(\n8_reg_n_0_[4] ),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[3]),
        .I4(\n33[12]_i_2__3_n_0 ),
        .O(\n33[12]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[12]_i_2__3 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n33[12]_i_2__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[13]_i_1__3 
       (.I0(n21[5]),
        .I1(\n8_reg_n_0_[5] ),
        .I2(\n33[14]_i_2__3_n_0 ),
        .O(\n33[13]_i_1__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[14]_i_1__3 
       (.I0(n21[6]),
        .I1(\n8_reg_n_0_[6] ),
        .I2(\n8_reg_n_0_[5] ),
        .I3(n21[5]),
        .I4(\n33[14]_i_2__3_n_0 ),
        .O(\n33[14]_i_1__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[14]_i_2__3 
       (.I0(\n33[12]_i_2__3_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n33[14]_i_2__3_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[15]_i_1__3 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n33[15]_i_2__3_n_0 ),
        .O(n30));
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[15]_i_2__3 
       (.I0(\n33[14]_i_2__3_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n33[15]_i_2__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[1]_i_1__3 
       (.I0(n29[1]),
        .I1(n10[1]),
        .I2(n10[0]),
        .I3(n29[0]),
        .O(n31[1]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[2]_i_1__3 
       (.I0(n29[2]),
        .I1(n10[2]),
        .I2(n10[1]),
        .I3(n29[1]),
        .I4(n10[0]),
        .I5(n29[0]),
        .O(\n33[2]_i_1__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[3]_i_1__3 
       (.I0(n29[3]),
        .I1(n10[3]),
        .I2(\n33[4]_i_2__3_n_0 ),
        .O(\n33[3]_i_1__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[4]_i_1__3 
       (.I0(n29[4]),
        .I1(n10[4]),
        .I2(n10[3]),
        .I3(n29[3]),
        .I4(\n33[4]_i_2__3_n_0 ),
        .O(\n33[4]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[4]_i_2__3 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n33[4]_i_2__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[5]_i_1__3 
       (.I0(n29[5]),
        .I1(n10[5]),
        .I2(\n33[6]_i_2__3_n_0 ),
        .O(\n33[5]_i_1__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[6]_i_1__3 
       (.I0(n29[6]),
        .I1(n10[6]),
        .I2(n10[5]),
        .I3(n29[5]),
        .I4(\n33[6]_i_2__3_n_0 ),
        .O(\n33[6]_i_1__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[6]_i_2__3 
       (.I0(\n33[4]_i_2__3_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n33[6]_i_2__3_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[7]_i_1__3 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n33[7]_i_2__3_n_0 ),
        .O(n31[7]));
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[7]_i_2__3 
       (.I0(\n33[6]_i_2__3_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n33[7]_i_2__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[9]_i_1__3 
       (.I0(n21[1]),
        .I1(\n8_reg_n_0_[1] ),
        .I2(\n8_reg_n_0_[0] ),
        .I3(n21[0]),
        .O(\n33[9]_i_1__3_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[0]),
        .Q(i1[15]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[10]_i_1__3_n_0 ),
        .Q(i1[24]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[11]_i_1__3_n_0 ),
        .Q(i1[25]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[12]_i_1__3_n_0 ),
        .Q(i1[26]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[13]_i_1__3_n_0 ),
        .Q(i1[27]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[14]_i_1__3_n_0 ),
        .Q(i1[28]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n30),
        .Q(i1[29]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[1]),
        .Q(i1[16]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[2]_i_1__3_n_0 ),
        .Q(i1[17]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[3]_i_1__3_n_0 ),
        .Q(i1[18]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[4]_i_1__3_n_0 ),
        .Q(i1[19]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[5]_i_1__3_n_0 ),
        .Q(i1[20]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[6]_i_1__3_n_0 ),
        .Q(i1[21]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[7]),
        .Q(i1[22]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[9]_i_1__3_n_0 ),
        .Q(i1[23]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[10]_i_1__3 
       (.I0(\n8_reg_n_0_[1] ),
        .I1(n21[1]),
        .I2(n21[0]),
        .I3(\n8_reg_n_0_[0] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(n341_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[11]_i_1__3 
       (.I0(\n37[12]_i_2__3_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .O(n341_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[12]_i_1__3 
       (.I0(\n8_reg_n_0_[3] ),
        .I1(n21[3]),
        .I2(\n37[12]_i_2__3_n_0 ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(n341_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[12]_i_2__3 
       (.I0(\n8_reg_n_0_[0] ),
        .I1(n21[0]),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n37[12]_i_2__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[13]_i_1__3 
       (.I0(\n37[14]_i_2__3_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(n341_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[14]_i_1__3 
       (.I0(\n8_reg_n_0_[5] ),
        .I1(n21[5]),
        .I2(\n37[14]_i_2__3_n_0 ),
        .I3(n21[6]),
        .I4(\n8_reg_n_0_[6] ),
        .O(n341_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[14]_i_2__3 
       (.I0(\n37[12]_i_2__3_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n37[14]_i_2__3_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[15]_i_1__3 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n37[15]_i_2__3_n_0 ),
        .O(n341_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[15]_i_2__3 
       (.I0(\n37[14]_i_2__3_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n37[15]_i_2__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[1]_i_1__3 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .O(n350_out[1]));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[2]_i_1__3 
       (.I0(n10[1]),
        .I1(n29[1]),
        .I2(n29[0]),
        .I3(n10[0]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(n350_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[3]_i_1__3 
       (.I0(\n37[4]_i_2__3_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .O(n350_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[4]_i_1__3 
       (.I0(n10[3]),
        .I1(n29[3]),
        .I2(\n37[4]_i_2__3_n_0 ),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(n350_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[4]_i_2__3 
       (.I0(n10[0]),
        .I1(n29[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n37[4]_i_2__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[5]_i_1__3 
       (.I0(\n37[6]_i_2__3_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(n350_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[6]_i_1__3 
       (.I0(n10[5]),
        .I1(n29[5]),
        .I2(\n37[6]_i_2__3_n_0 ),
        .I3(n29[6]),
        .I4(n10[6]),
        .O(n350_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[6]_i_2__3 
       (.I0(\n37[4]_i_2__3_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n37[6]_i_2__3_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[7]_i_1__3 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n37[7]_i_2__3_n_0 ),
        .O(n350_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[7]_i_2__3 
       (.I0(\n37[6]_i_2__3_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n37[7]_i_2__3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n37[8]_i_1__0 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .O(n341_out[0]));
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[9]_i_1__3 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .O(n341_out[1]));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[2]),
        .Q(i1[9]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[3]),
        .Q(i1[10]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[4]),
        .Q(i1[11]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[5]),
        .Q(i1[12]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[6]),
        .Q(i1[13]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[7]),
        .Q(i1[14]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[1]),
        .Q(i1[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[2]),
        .Q(i1[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[3]),
        .Q(i1[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[4]),
        .Q(i1[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[5]),
        .Q(i1[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[6]),
        .Q(i1[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[7]),
        .Q(i1[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[0]),
        .Q(i1[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[1]),
        .Q(i1[8]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[0]),
        .Q(\n4_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[1]),
        .Q(\n4_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[2]),
        .Q(\n4_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[3]),
        .Q(\n4_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[4]),
        .Q(\n4_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[5]),
        .Q(\n4_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[6]),
        .Q(\n4_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s6_3[7]),
        .Q(\n4_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[0]),
        .Q(\n7_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[1]),
        .Q(\n7_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[2]),
        .Q(\n7_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[3]),
        .Q(\n7_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[4]),
        .Q(\n7_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[5]),
        .Q(\n7_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[6]),
        .Q(\n7_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[7]),
        .Q(\n7_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[0] ),
        .Q(\n8_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[1] ),
        .Q(\n8_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[2] ),
        .Q(\n8_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[3] ),
        .Q(\n8_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[4] ),
        .Q(\n8_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[5] ),
        .Q(\n8_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[6] ),
        .Q(\n8_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[7] ),
        .Q(\n8_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[0] ),
        .Q(\n9_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[1] ),
        .Q(\n9_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[2] ),
        .Q(\n9_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[3] ),
        .Q(\n9_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[4] ),
        .Q(\n9_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[5] ),
        .Q(\n9_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[6] ),
        .Q(\n9_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[7] ),
        .Q(\n9_reg_n_0_[7] ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_13" *) 
module switch_elements_cf_fft_512_8_13
   (\n9_reg[0] ,
    s4_3,
    rst_i,
    enable_i,
    clk_i,
    s5_3,
    D);
  output [15:0]\n9_reg[0] ;
  output [15:0]s4_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]s5_3;
  input [15:0]D;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire [15:0]n33;
  wire [15:1]n37;
  wire n4;
  wire [15:0]\n9_reg[0] ;
  wire rst_i;
  wire s29_n_0;
  wire [15:0]s4_3;
  wire [15:0]s5_3;

  switch_elements_cf_fft_512_8_31_10 s25
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i8(i8),
        .n4(n4),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_14 s26
       (.D(D),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:1],n37[15:9],n37[7:1],n33[0]}),
        .rst_i(rst_i),
        .s5_3(s5_3));
  switch_elements_cf_fft_512_8_26_11 s28
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:1],n37[15:9],n37[7:1],n33[0]}),
        .i8(i8),
        .\n1_reg[0] (s29_n_0),
        .n4(n4),
        .\n9_reg[0] (\n9_reg[0] ),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_27_12 s29
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:1],n37[15:9],n37[7:1],n33[0]}),
        .i8(i8),
        .\n9_reg[0]_0 (s29_n_0),
        .rst_i(rst_i),
        .s4_3(s4_3));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_14" *) 
module switch_elements_cf_fft_512_8_14
   (i1,
    rst_i,
    enable_i,
    clk_i,
    s5_3,
    D);
  output [29:0]i1;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]s5_3;
  input [15:0]D;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [7:0]n10;
  wire n14__21_carry__0_i_1__1_n_0;
  wire n14__21_carry__0_i_2_n_0;
  wire n14__21_carry__0_i_3__1_n_0;
  wire n14__21_carry__0_i_4_n_0;
  wire n14__21_carry__0_n_14;
  wire n14__21_carry__0_n_15;
  wire n14__21_carry__0_n_5;
  wire n14__21_carry__0_n_7;
  wire n14__21_carry_i_10_n_0;
  wire n14__21_carry_i_11__1_n_0;
  wire n14__21_carry_i_1_n_0;
  wire n14__21_carry_i_2_n_0;
  wire n14__21_carry_i_3_n_0;
  wire n14__21_carry_i_4_n_0;
  wire n14__21_carry_i_5_n_0;
  wire n14__21_carry_i_6__1_n_0;
  wire n14__21_carry_i_7__1_n_0;
  wire n14__21_carry_i_8_n_0;
  wire n14__21_carry_i_9__1_n_0;
  wire n14__21_carry_n_0;
  wire n14__21_carry_n_1;
  wire n14__21_carry_n_10;
  wire n14__21_carry_n_11;
  wire n14__21_carry_n_12;
  wire n14__21_carry_n_13;
  wire n14__21_carry_n_14;
  wire n14__21_carry_n_2;
  wire n14__21_carry_n_3;
  wire n14__21_carry_n_4;
  wire n14__21_carry_n_5;
  wire n14__21_carry_n_6;
  wire n14__21_carry_n_7;
  wire n14__21_carry_n_8;
  wire n14__21_carry_n_9;
  wire n14__47_carry_i_1_n_0;
  wire n14__47_carry_i_2_n_0;
  wire n14__47_carry_i_3__1_n_0;
  wire n14__47_carry_i_4__1_n_0;
  wire n14__47_carry_i_5__1_n_0;
  wire n14__47_carry_i_6_n_0;
  wire n14__47_carry_n_1;
  wire n14__47_carry_n_10;
  wire n14__47_carry_n_11;
  wire n14__47_carry_n_12;
  wire n14__47_carry_n_13;
  wire n14__47_carry_n_14;
  wire n14__47_carry_n_15;
  wire n14__47_carry_n_2;
  wire n14__47_carry_n_3;
  wire n14__47_carry_n_4;
  wire n14__47_carry_n_5;
  wire n14__47_carry_n_6;
  wire n14__47_carry_n_7;
  wire n14__47_carry_n_8;
  wire n14__47_carry_n_9;
  wire n14__67_carry__0_i_1_n_0;
  wire n14__67_carry__0_i_2_n_0;
  wire n14__67_carry__0_i_3_n_0;
  wire n14__67_carry__0_i_4_n_0;
  wire n14__67_carry__0_i_5_n_0;
  wire n14__67_carry__0_i_6_n_0;
  wire n14__67_carry__0_i_7_n_0;
  wire n14__67_carry__0_n_5;
  wire n14__67_carry__0_n_6;
  wire n14__67_carry__0_n_7;
  wire n14__67_carry_i_10_n_0;
  wire n14__67_carry_i_11_n_0;
  wire n14__67_carry_i_12_n_0;
  wire n14__67_carry_i_13_n_0;
  wire n14__67_carry_i_14_n_0;
  wire n14__67_carry_i_15_n_0;
  wire n14__67_carry_i_1_n_0;
  wire n14__67_carry_i_2_n_0;
  wire n14__67_carry_i_3_n_0;
  wire n14__67_carry_i_4_n_0;
  wire n14__67_carry_i_5_n_0;
  wire n14__67_carry_i_6_n_0;
  wire n14__67_carry_i_7_n_0;
  wire n14__67_carry_i_8_n_0;
  wire n14__67_carry_i_9_n_0;
  wire n14__67_carry_n_0;
  wire n14__67_carry_n_1;
  wire n14__67_carry_n_2;
  wire n14__67_carry_n_3;
  wire n14__67_carry_n_4;
  wire n14__67_carry_n_5;
  wire n14__67_carry_n_6;
  wire n14__67_carry_n_7;
  wire n14_carry__0_i_1_n_0;
  wire n14_carry__0_i_2_n_0;
  wire n14_carry__0_i_3__1_n_0;
  wire n14_carry__0_i_4_n_0;
  wire n14_carry__0_n_14;
  wire n14_carry__0_n_15;
  wire n14_carry__0_n_5;
  wire n14_carry__0_n_7;
  wire n14_carry_i_10_n_0;
  wire n14_carry_i_11_n_0;
  wire n14_carry_i_12_n_0;
  wire n14_carry_i_1_n_0;
  wire n14_carry_i_2_n_0;
  wire n14_carry_i_3_n_0;
  wire n14_carry_i_4_n_0;
  wire n14_carry_i_5_n_0;
  wire n14_carry_i_6_n_0;
  wire n14_carry_i_7__1_n_0;
  wire n14_carry_i_8__1_n_0;
  wire n14_carry_i_9_n_0;
  wire n14_carry_n_0;
  wire n14_carry_n_1;
  wire n14_carry_n_10;
  wire n14_carry_n_11;
  wire n14_carry_n_12;
  wire n14_carry_n_15;
  wire n14_carry_n_2;
  wire n14_carry_n_3;
  wire n14_carry_n_4;
  wire n14_carry_n_5;
  wire n14_carry_n_6;
  wire n14_carry_n_7;
  wire n14_carry_n_8;
  wire n14_carry_n_9;
  wire [7:0]n15;
  wire \n16_reg_n_0_[0] ;
  wire \n16_reg_n_0_[1] ;
  wire \n16_reg_n_0_[2] ;
  wire \n16_reg_n_0_[3] ;
  wire \n16_reg_n_0_[4] ;
  wire \n16_reg_n_0_[5] ;
  wire \n16_reg_n_0_[6] ;
  wire \n16_reg_n_0_[7] ;
  wire \n1_reg_n_0_[0] ;
  wire \n1_reg_n_0_[1] ;
  wire \n1_reg_n_0_[2] ;
  wire \n1_reg_n_0_[3] ;
  wire \n1_reg_n_0_[4] ;
  wire \n1_reg_n_0_[5] ;
  wire \n1_reg_n_0_[6] ;
  wire \n1_reg_n_0_[7] ;
  wire [7:0]n2;
  wire [7:0]n202_out;
  wire n20_carry_i_1_n_0;
  wire n20_carry_i_2_n_0;
  wire n20_carry_i_3_n_0;
  wire n20_carry_i_4_n_0;
  wire n20_carry_i_5_n_0;
  wire n20_carry_i_6_n_0;
  wire n20_carry_i_7_n_0;
  wire n20_carry_i_8_n_0;
  wire n20_carry_n_1;
  wire n20_carry_n_2;
  wire n20_carry_n_3;
  wire n20_carry_n_4;
  wire n20_carry_n_5;
  wire n20_carry_n_6;
  wire n20_carry_n_7;
  wire [7:0]n21;
  wire n22__0_n_0;
  wire n22__1_n_0;
  wire n22__2_n_0;
  wire n22__3_n_0;
  wire n22__4_n_0;
  wire n22__5_n_0;
  wire n22__6_n_0;
  wire n22_n_0;
  wire n25__17_carry__0_i_1__1_n_0;
  wire n25__17_carry__0_i_2_n_0;
  wire n25__17_carry__0_i_3__1_n_0;
  wire n25__17_carry__0_i_4_n_0;
  wire n25__17_carry__0_n_14;
  wire n25__17_carry__0_n_15;
  wire n25__17_carry__0_n_5;
  wire n25__17_carry__0_n_7;
  wire n25__17_carry_i_10_n_0;
  wire n25__17_carry_i_11__1_n_0;
  wire n25__17_carry_i_1_n_0;
  wire n25__17_carry_i_2_n_0;
  wire n25__17_carry_i_3_n_0;
  wire n25__17_carry_i_4_n_0;
  wire n25__17_carry_i_5_n_0;
  wire n25__17_carry_i_6__1_n_0;
  wire n25__17_carry_i_7__1_n_0;
  wire n25__17_carry_i_8_n_0;
  wire n25__17_carry_i_9__1_n_0;
  wire n25__17_carry_n_0;
  wire n25__17_carry_n_1;
  wire n25__17_carry_n_10;
  wire n25__17_carry_n_11;
  wire n25__17_carry_n_12;
  wire n25__17_carry_n_13;
  wire n25__17_carry_n_14;
  wire n25__17_carry_n_2;
  wire n25__17_carry_n_3;
  wire n25__17_carry_n_4;
  wire n25__17_carry_n_5;
  wire n25__17_carry_n_6;
  wire n25__17_carry_n_7;
  wire n25__17_carry_n_8;
  wire n25__17_carry_n_9;
  wire n25__47_carry_i_1_n_0;
  wire n25__47_carry_i_2_n_0;
  wire n25__47_carry_i_3__1_n_0;
  wire n25__47_carry_i_4__1_n_0;
  wire n25__47_carry_i_5__1_n_0;
  wire n25__47_carry_i_6_n_0;
  wire n25__47_carry_n_1;
  wire n25__47_carry_n_10;
  wire n25__47_carry_n_11;
  wire n25__47_carry_n_12;
  wire n25__47_carry_n_13;
  wire n25__47_carry_n_14;
  wire n25__47_carry_n_15;
  wire n25__47_carry_n_2;
  wire n25__47_carry_n_3;
  wire n25__47_carry_n_4;
  wire n25__47_carry_n_5;
  wire n25__47_carry_n_6;
  wire n25__47_carry_n_7;
  wire n25__47_carry_n_8;
  wire n25__47_carry_n_9;
  wire n25__67_carry__0_i_1_n_0;
  wire n25__67_carry__0_i_2_n_0;
  wire n25__67_carry__0_i_3_n_0;
  wire n25__67_carry__0_i_4_n_0;
  wire n25__67_carry__0_i_5_n_0;
  wire n25__67_carry__0_i_6_n_0;
  wire n25__67_carry__0_i_7_n_0;
  wire n25__67_carry__0_n_5;
  wire n25__67_carry__0_n_6;
  wire n25__67_carry__0_n_7;
  wire n25__67_carry_i_10_n_0;
  wire n25__67_carry_i_11_n_0;
  wire n25__67_carry_i_12_n_0;
  wire n25__67_carry_i_13_n_0;
  wire n25__67_carry_i_14_n_0;
  wire n25__67_carry_i_15_n_0;
  wire n25__67_carry_i_1_n_0;
  wire n25__67_carry_i_2_n_0;
  wire n25__67_carry_i_3_n_0;
  wire n25__67_carry_i_4_n_0;
  wire n25__67_carry_i_5_n_0;
  wire n25__67_carry_i_6_n_0;
  wire n25__67_carry_i_7_n_0;
  wire n25__67_carry_i_8_n_0;
  wire n25__67_carry_i_9_n_0;
  wire n25__67_carry_n_0;
  wire n25__67_carry_n_1;
  wire n25__67_carry_n_2;
  wire n25__67_carry_n_3;
  wire n25__67_carry_n_4;
  wire n25__67_carry_n_5;
  wire n25__67_carry_n_6;
  wire n25__67_carry_n_7;
  wire n25_carry__0_i_1_n_0;
  wire n25_carry__0_i_2_n_0;
  wire n25_carry__0_i_3__1_n_0;
  wire n25_carry__0_i_4_n_0;
  wire n25_carry__0_n_14;
  wire n25_carry__0_n_15;
  wire n25_carry__0_n_5;
  wire n25_carry__0_n_7;
  wire n25_carry_i_10_n_0;
  wire n25_carry_i_11_n_0;
  wire n25_carry_i_12_n_0;
  wire n25_carry_i_1_n_0;
  wire n25_carry_i_2_n_0;
  wire n25_carry_i_3_n_0;
  wire n25_carry_i_4_n_0;
  wire n25_carry_i_5_n_0;
  wire n25_carry_i_6_n_0;
  wire n25_carry_i_7__1_n_0;
  wire n25_carry_i_8__1_n_0;
  wire n25_carry_i_9_n_0;
  wire n25_carry_n_0;
  wire n25_carry_n_1;
  wire n25_carry_n_10;
  wire n25_carry_n_11;
  wire n25_carry_n_12;
  wire n25_carry_n_15;
  wire n25_carry_n_2;
  wire n25_carry_n_3;
  wire n25_carry_n_4;
  wire n25_carry_n_5;
  wire n25_carry_n_6;
  wire n25_carry_n_7;
  wire n25_carry_n_8;
  wire n25_carry_n_9;
  wire [7:0]n26;
  wire [7:0]n27;
  wire [7:0]n29;
  wire [7:0]n30;
  wire [7:0]n31;
  wire \n33[10]_i_1__2_n_0 ;
  wire \n33[11]_i_1__2_n_0 ;
  wire \n33[12]_i_1__2_n_0 ;
  wire \n33[12]_i_2__2_n_0 ;
  wire \n33[13]_i_1__2_n_0 ;
  wire \n33[14]_i_1__2_n_0 ;
  wire \n33[14]_i_2__2_n_0 ;
  wire \n33[15]_i_2__2_n_0 ;
  wire \n33[2]_i_1__2_n_0 ;
  wire \n33[3]_i_1__2_n_0 ;
  wire \n33[4]_i_1__2_n_0 ;
  wire \n33[4]_i_2__2_n_0 ;
  wire \n33[5]_i_1__2_n_0 ;
  wire \n33[6]_i_1__2_n_0 ;
  wire \n33[6]_i_2__2_n_0 ;
  wire \n33[7]_i_2__2_n_0 ;
  wire \n33[9]_i_1__2_n_0 ;
  wire [7:1]n341_out;
  wire [7:1]n350_out;
  wire \n37[12]_i_2__2_n_0 ;
  wire \n37[14]_i_2__2_n_0 ;
  wire \n37[15]_i_2__2_n_0 ;
  wire \n37[4]_i_2__2_n_0 ;
  wire \n37[6]_i_2__2_n_0 ;
  wire \n37[7]_i_2__2_n_0 ;
  wire \n4_reg_n_0_[0] ;
  wire \n4_reg_n_0_[1] ;
  wire \n4_reg_n_0_[2] ;
  wire \n4_reg_n_0_[3] ;
  wire \n4_reg_n_0_[4] ;
  wire \n4_reg_n_0_[5] ;
  wire \n4_reg_n_0_[6] ;
  wire \n4_reg_n_0_[7] ;
  wire \n7_reg_n_0_[0] ;
  wire \n7_reg_n_0_[1] ;
  wire \n7_reg_n_0_[2] ;
  wire \n7_reg_n_0_[3] ;
  wire \n7_reg_n_0_[4] ;
  wire \n7_reg_n_0_[5] ;
  wire \n7_reg_n_0_[6] ;
  wire \n7_reg_n_0_[7] ;
  wire \n8_reg_n_0_[0] ;
  wire \n8_reg_n_0_[1] ;
  wire \n8_reg_n_0_[2] ;
  wire \n8_reg_n_0_[3] ;
  wire \n8_reg_n_0_[4] ;
  wire \n8_reg_n_0_[5] ;
  wire \n8_reg_n_0_[6] ;
  wire \n8_reg_n_0_[7] ;
  wire \n9_reg_n_0_[0] ;
  wire \n9_reg_n_0_[1] ;
  wire \n9_reg_n_0_[2] ;
  wire \n9_reg_n_0_[3] ;
  wire \n9_reg_n_0_[4] ;
  wire \n9_reg_n_0_[5] ;
  wire \n9_reg_n_0_[6] ;
  wire \n9_reg_n_0_[7] ;
  wire rst_i;
  wire [15:0]s5_3;
  wire [0:0]NLW_n14__21_carry_O_UNCONNECTED;
  wire [7:1]NLW_n14__21_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n14__21_carry__0_O_UNCONNECTED;
  wire [7:7]NLW_n14__47_carry_CO_UNCONNECTED;
  wire [3:0]NLW_n14__67_carry_O_UNCONNECTED;
  wire [7:3]NLW_n14__67_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n14__67_carry__0_O_UNCONNECTED;
  wire [2:1]NLW_n14_carry_O_UNCONNECTED;
  wire [7:1]NLW_n14_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n14_carry__0_O_UNCONNECTED;
  wire [7:7]NLW_n20_carry_CO_UNCONNECTED;
  wire [0:0]NLW_n25__17_carry_O_UNCONNECTED;
  wire [7:1]NLW_n25__17_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n25__17_carry__0_O_UNCONNECTED;
  wire [7:7]NLW_n25__47_carry_CO_UNCONNECTED;
  wire [3:0]NLW_n25__67_carry_O_UNCONNECTED;
  wire [7:3]NLW_n25__67_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n25__67_carry__0_O_UNCONNECTED;
  wire [2:1]NLW_n25_carry_O_UNCONNECTED;
  wire [7:1]NLW_n25_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n25_carry__0_O_UNCONNECTED;

  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[0] ),
        .Q(n10[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[1] ),
        .Q(n10[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[2] ),
        .Q(n10[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[3] ),
        .Q(n10[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[4] ),
        .Q(n10[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[5] ),
        .Q(n10[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[6] ),
        .Q(n10[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[7] ),
        .Q(n10[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__21_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__21_carry_n_0,n14__21_carry_n_1,n14__21_carry_n_2,n14__21_carry_n_3,n14__21_carry_n_4,n14__21_carry_n_5,n14__21_carry_n_6,n14__21_carry_n_7}),
        .DI({n14_carry_i_1_n_0,n14__21_carry_i_1_n_0,n14__21_carry_i_2_n_0,n14__21_carry_i_3_n_0,n14__21_carry_i_4_n_0,n22__4_n_0,n22__5_n_0,1'b0}),
        .O({n14__21_carry_n_8,n14__21_carry_n_9,n14__21_carry_n_10,n14__21_carry_n_11,n14__21_carry_n_12,n14__21_carry_n_13,n14__21_carry_n_14,NLW_n14__21_carry_O_UNCONNECTED[0]}),
        .S({n14__21_carry_i_5_n_0,n14__21_carry_i_6__1_n_0,n14__21_carry_i_7__1_n_0,n14__21_carry_i_8_n_0,n14__21_carry_i_9__1_n_0,n14__21_carry_i_10_n_0,n14__21_carry_i_11__1_n_0,n22__6_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__21_carry__0
       (.CI(n14__21_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__21_carry__0_CO_UNCONNECTED[7:3],n14__21_carry__0_n_5,NLW_n14__21_carry__0_CO_UNCONNECTED[1],n14__21_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14__21_carry__0_i_1__1_n_0,n14__21_carry__0_i_2_n_0}),
        .O({NLW_n14__21_carry__0_O_UNCONNECTED[7:2],n14__21_carry__0_n_14,n14__21_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n14__21_carry__0_i_3__1_n_0,n14__21_carry__0_i_4_n_0}));
  LUT2 #(
    .INIT(4'h2)) 
    n14__21_carry__0_i_1__1
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(n14__21_carry__0_i_1__1_n_0));
  LUT3 #(
    .INIT(8'h8E)) 
    n14__21_carry__0_i_2
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(n14__21_carry__0_i_2_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    n14__21_carry__0_i_3__1
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(n14__21_carry__0_i_3__1_n_0));
  LUT3 #(
    .INIT(8'h4D)) 
    n14__21_carry__0_i_4
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(n14__21_carry__0_i_4_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14__21_carry_i_1
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(n22__1_n_0),
        .O(n14__21_carry_i_1_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    n14__21_carry_i_10
       (.I0(n22__6_n_0),
        .I1(n22__5_n_0),
        .I2(n22__4_n_0),
        .O(n14__21_carry_i_10_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n14__21_carry_i_11__1
       (.I0(n22__5_n_0),
        .I1(n22__6_n_0),
        .O(n14__21_carry_i_11__1_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14__21_carry_i_2
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__2_n_0),
        .O(n14__21_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14__21_carry_i_3
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(n22__3_n_0),
        .O(n14__21_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    n14__21_carry_i_4
       (.I0(n22__4_n_0),
        .I1(n22__5_n_0),
        .I2(n22__3_n_0),
        .O(n14__21_carry_i_4_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    n14__21_carry_i_5
       (.I0(n14_carry_i_1_n_0),
        .I1(n22__0_n_0),
        .I2(n22__1_n_0),
        .I3(n22_n_0),
        .O(n14__21_carry_i_5_n_0));
  (* HLUTNM = "lutpair90" *) 
  LUT4 #(
    .INIT(16'h781E)) 
    n14__21_carry_i_6__1
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(n22__3_n_0),
        .O(n14__21_carry_i_6__1_n_0));
  LUT4 #(
    .INIT(16'h2BD4)) 
    n14__21_carry_i_7__1
       (.I0(n22__4_n_0),
        .I1(n22__2_n_0),
        .I2(n22__3_n_0),
        .I3(n22__1_n_0),
        .O(n14__21_carry_i_7__1_n_0));
  LUT4 #(
    .INIT(16'h2BD4)) 
    n14__21_carry_i_8
       (.I0(n22__5_n_0),
        .I1(n22__3_n_0),
        .I2(n22__4_n_0),
        .I3(n22__2_n_0),
        .O(n14__21_carry_i_8_n_0));
  LUT4 #(
    .INIT(16'h6696)) 
    n14__21_carry_i_9__1
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__5_n_0),
        .I3(n22__6_n_0),
        .O(n14__21_carry_i_9__1_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__47_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__47_carry_CO_UNCONNECTED[7],n14__47_carry_n_1,n14__47_carry_n_2,n14__47_carry_n_3,n14__47_carry_n_4,n14__47_carry_n_5,n14__47_carry_n_6,n14__47_carry_n_7}),
        .DI({1'b0,n22__0_n_0,n22__1_n_0,n22__2_n_0,n22__3_n_0,1'b1,1'b0,1'b1}),
        .O({n14__47_carry_n_8,n14__47_carry_n_9,n14__47_carry_n_10,n14__47_carry_n_11,n14__47_carry_n_12,n14__47_carry_n_13,n14__47_carry_n_14,n14__47_carry_n_15}),
        .S({n14__47_carry_i_1_n_0,n14__47_carry_i_2_n_0,n14__47_carry_i_3__1_n_0,n14__47_carry_i_4__1_n_0,n14__47_carry_i_5__1_n_0,n22__3_n_0,n22__4_n_0,n14__47_carry_i_6_n_0}));
  LUT1 #(
    .INIT(2'h1)) 
    n14__47_carry_i_1
       (.I0(n22_n_0),
        .O(n14__47_carry_i_1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n14__47_carry_i_2
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(n14__47_carry_i_2_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n14__47_carry_i_3__1
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .O(n14__47_carry_i_3__1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n14__47_carry_i_4__1
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .O(n14__47_carry_i_4__1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n14__47_carry_i_5__1
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .O(n14__47_carry_i_5__1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    n14__47_carry_i_6
       (.I0(n22__5_n_0),
        .O(n14__47_carry_i_6_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__67_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__67_carry_n_0,n14__67_carry_n_1,n14__67_carry_n_2,n14__67_carry_n_3,n14__67_carry_n_4,n14__67_carry_n_5,n14__67_carry_n_6,n14__67_carry_n_7}),
        .DI({n14__67_carry_i_1_n_0,n14__67_carry_i_2_n_0,n14__67_carry_i_3_n_0,n14__67_carry_i_4_n_0,n14__67_carry_i_5_n_0,n14__67_carry_i_6_n_0,n14__67_carry_i_7_n_0,1'b0}),
        .O({n15[3:0],NLW_n14__67_carry_O_UNCONNECTED[3:0]}),
        .S({n14__67_carry_i_8_n_0,n14__67_carry_i_9_n_0,n14__67_carry_i_10_n_0,n14__67_carry_i_11_n_0,n14__67_carry_i_12_n_0,n14__67_carry_i_13_n_0,n14__67_carry_i_14_n_0,n14__67_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__67_carry__0
       (.CI(n14__67_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__67_carry__0_CO_UNCONNECTED[7:3],n14__67_carry__0_n_5,n14__67_carry__0_n_6,n14__67_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n14__67_carry__0_i_1_n_0,n14__67_carry__0_i_2_n_0,n14__67_carry__0_i_3_n_0}),
        .O({NLW_n14__67_carry__0_O_UNCONNECTED[7:4],n15[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n14__67_carry__0_i_4_n_0,n14__67_carry__0_i_5_n_0,n14__67_carry__0_i_6_n_0,n14__67_carry__0_i_7_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry__0_i_1
       (.I0(n14__21_carry__0_n_14),
        .I1(n14__47_carry_n_10),
        .O(n14__67_carry__0_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry__0_i_2
       (.I0(n14__21_carry__0_n_15),
        .I1(n14__47_carry_n_11),
        .O(n14__67_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14__67_carry__0_i_3
       (.I0(n14__47_carry_n_12),
        .I1(n14__21_carry_n_8),
        .I2(n14_carry__0_n_5),
        .O(n14__67_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n14__67_carry__0_i_4
       (.I0(n14__21_carry__0_n_5),
        .I1(n14__47_carry_n_9),
        .I2(n14__47_carry_n_8),
        .O(n14__67_carry__0_i_4_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__67_carry__0_i_5
       (.I0(n14__21_carry__0_n_14),
        .I1(n14__47_carry_n_10),
        .I2(n14__47_carry_n_9),
        .I3(n14__21_carry__0_n_5),
        .O(n14__67_carry__0_i_5_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__67_carry__0_i_6
       (.I0(n14__21_carry__0_n_15),
        .I1(n14__47_carry_n_11),
        .I2(n14__47_carry_n_10),
        .I3(n14__21_carry__0_n_14),
        .O(n14__67_carry__0_i_6_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n14__67_carry__0_i_7
       (.I0(n14_carry__0_n_5),
        .I1(n14__21_carry_n_8),
        .I2(n14__47_carry_n_12),
        .I3(n14__47_carry_n_11),
        .I4(n14__21_carry__0_n_15),
        .O(n14__67_carry__0_i_7_n_0));
  (* HLUTNM = "lutpair39" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__67_carry_i_1
       (.I0(n14__47_carry_n_13),
        .I1(n14__21_carry_n_9),
        .I2(n14_carry__0_n_14),
        .O(n14__67_carry_i_1_n_0));
  (* HLUTNM = "lutpair38" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__67_carry_i_10
       (.I0(n14__47_carry_n_14),
        .I1(n14__21_carry_n_10),
        .I2(n14_carry__0_n_15),
        .I3(n14__67_carry_i_3_n_0),
        .O(n14__67_carry_i_10_n_0));
  (* HLUTNM = "lutpair37" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__67_carry_i_11
       (.I0(n14__47_carry_n_15),
        .I1(n14__21_carry_n_11),
        .I2(n14_carry_n_8),
        .I3(n14__67_carry_i_4_n_0),
        .O(n14__67_carry_i_11_n_0));
  (* HLUTNM = "lutpair36" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__67_carry_i_12
       (.I0(n14_carry_n_15),
        .I1(n14__21_carry_n_12),
        .I2(n14_carry_n_9),
        .I3(n14__67_carry_i_5_n_0),
        .O(n14__67_carry_i_12_n_0));
  (* HLUTNM = "lutpair91" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n14__67_carry_i_13
       (.I0(n14__21_carry_n_13),
        .I1(n14_carry_n_10),
        .I2(n14_carry_n_11),
        .I3(n14__21_carry_n_14),
        .O(n14__67_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__67_carry_i_14
       (.I0(n14_carry_n_12),
        .I1(n22__6_n_0),
        .I2(n14__21_carry_n_14),
        .I3(n14_carry_n_11),
        .O(n14__67_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n14__67_carry_i_15
       (.I0(n14_carry_n_12),
        .I1(n22__6_n_0),
        .O(n14__67_carry_i_15_n_0));
  (* HLUTNM = "lutpair38" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__67_carry_i_2
       (.I0(n14__47_carry_n_14),
        .I1(n14__21_carry_n_10),
        .I2(n14_carry__0_n_15),
        .O(n14__67_carry_i_2_n_0));
  (* HLUTNM = "lutpair37" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__67_carry_i_3
       (.I0(n14__47_carry_n_15),
        .I1(n14__21_carry_n_11),
        .I2(n14_carry_n_8),
        .O(n14__67_carry_i_3_n_0));
  (* HLUTNM = "lutpair36" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__67_carry_i_4
       (.I0(n14_carry_n_15),
        .I1(n14__21_carry_n_12),
        .I2(n14_carry_n_9),
        .O(n14__67_carry_i_4_n_0));
  (* HLUTNM = "lutpair91" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry_i_5
       (.I0(n14__21_carry_n_13),
        .I1(n14_carry_n_10),
        .O(n14__67_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry_i_6
       (.I0(n14_carry_n_11),
        .I1(n14__21_carry_n_14),
        .O(n14__67_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry_i_7
       (.I0(n14_carry_n_12),
        .I1(n22__6_n_0),
        .O(n14__67_carry_i_7_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n14__67_carry_i_8
       (.I0(n14__67_carry_i_1_n_0),
        .I1(n14__21_carry_n_8),
        .I2(n14__47_carry_n_12),
        .I3(n14_carry__0_n_5),
        .O(n14__67_carry_i_8_n_0));
  (* HLUTNM = "lutpair39" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__67_carry_i_9
       (.I0(n14__47_carry_n_13),
        .I1(n14__21_carry_n_9),
        .I2(n14_carry__0_n_14),
        .I3(n14__67_carry_i_2_n_0),
        .O(n14__67_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14_carry_n_0,n14_carry_n_1,n14_carry_n_2,n14_carry_n_3,n14_carry_n_4,n14_carry_n_5,n14_carry_n_6,n14_carry_n_7}),
        .DI({n14_carry_i_1_n_0,n14_carry_i_2_n_0,n14_carry_i_3_n_0,n14_carry_i_4_n_0,n14_carry_i_5_n_0,n22__4_n_0,n22__5_n_0,1'b0}),
        .O({n14_carry_n_8,n14_carry_n_9,n14_carry_n_10,n14_carry_n_11,n14_carry_n_12,NLW_n14_carry_O_UNCONNECTED[2:1],n14_carry_n_15}),
        .S({n14_carry_i_6_n_0,n14_carry_i_7__1_n_0,n14_carry_i_8__1_n_0,n14_carry_i_9_n_0,n14_carry_i_10_n_0,n14_carry_i_11_n_0,n14_carry_i_12_n_0,n22__6_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14_carry__0
       (.CI(n14_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14_carry__0_CO_UNCONNECTED[7:3],n14_carry__0_n_5,NLW_n14_carry__0_CO_UNCONNECTED[1],n14_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14_carry__0_i_1_n_0,n14_carry__0_i_2_n_0}),
        .O({NLW_n14_carry__0_O_UNCONNECTED[7:2],n14_carry__0_n_14,n14_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n14_carry__0_i_3__1_n_0,n14_carry__0_i_4_n_0}));
  LUT2 #(
    .INIT(4'h2)) 
    n14_carry__0_i_1
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(n14_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h8E)) 
    n14_carry__0_i_2
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(n14_carry__0_i_2_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    n14_carry__0_i_3__1
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(n14_carry__0_i_3__1_n_0));
  LUT3 #(
    .INIT(8'h4D)) 
    n14_carry__0_i_4
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(n14_carry__0_i_4_n_0));
  (* HLUTNM = "lutpair90" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14_carry_i_1
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .O(n14_carry_i_1_n_0));
  LUT4 #(
    .INIT(16'h6696)) 
    n14_carry_i_10
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__5_n_0),
        .I3(n22__6_n_0),
        .O(n14_carry_i_10_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    n14_carry_i_11
       (.I0(n22__6_n_0),
        .I1(n22__5_n_0),
        .I2(n22__4_n_0),
        .O(n14_carry_i_11_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n14_carry_i_12
       (.I0(n22__5_n_0),
        .I1(n22__6_n_0),
        .O(n14_carry_i_12_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14_carry_i_2
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(n22__1_n_0),
        .O(n14_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14_carry_i_3
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__2_n_0),
        .O(n14_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14_carry_i_4
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(n22__3_n_0),
        .O(n14_carry_i_4_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    n14_carry_i_5
       (.I0(n22__4_n_0),
        .I1(n22__5_n_0),
        .I2(n22__3_n_0),
        .O(n14_carry_i_5_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    n14_carry_i_6
       (.I0(n14_carry_i_1_n_0),
        .I1(n22__0_n_0),
        .I2(n22__1_n_0),
        .I3(n22_n_0),
        .O(n14_carry_i_6_n_0));
  LUT4 #(
    .INIT(16'h2BD4)) 
    n14_carry_i_7__1
       (.I0(n22__3_n_0),
        .I1(n22__1_n_0),
        .I2(n22__2_n_0),
        .I3(n22__0_n_0),
        .O(n14_carry_i_7__1_n_0));
  LUT4 #(
    .INIT(16'h2BD4)) 
    n14_carry_i_8__1
       (.I0(n22__4_n_0),
        .I1(n22__2_n_0),
        .I2(n22__3_n_0),
        .I3(n22__1_n_0),
        .O(n14_carry_i_8__1_n_0));
  LUT4 #(
    .INIT(16'h2BD4)) 
    n14_carry_i_9
       (.I0(n22__5_n_0),
        .I1(n22__3_n_0),
        .I2(n22__4_n_0),
        .I3(n22__2_n_0),
        .O(n14_carry_i_9_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[0]),
        .Q(\n16_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[1]),
        .Q(\n16_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[2]),
        .Q(\n16_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[3]),
        .Q(\n16_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[4]),
        .Q(\n16_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[5]),
        .Q(\n16_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[6]),
        .Q(\n16_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[7]),
        .Q(\n16_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[0]),
        .Q(\n1_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[10]),
        .Q(n2[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[11]),
        .Q(n2[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[12]),
        .Q(n2[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[13]),
        .Q(n2[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[14]),
        .Q(n2[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[15]),
        .Q(n2[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[1]),
        .Q(\n1_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[2]),
        .Q(\n1_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[3]),
        .Q(\n1_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[4]),
        .Q(\n1_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[5]),
        .Q(\n1_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[6]),
        .Q(\n1_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[7]),
        .Q(\n1_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[8]),
        .Q(n2[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[9]),
        .Q(n2[1]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n20_carry
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({NLW_n20_carry_CO_UNCONNECTED[7],n20_carry_n_1,n20_carry_n_2,n20_carry_n_3,n20_carry_n_4,n20_carry_n_5,n20_carry_n_6,n20_carry_n_7}),
        .DI({1'b0,\n16_reg_n_0_[6] ,\n16_reg_n_0_[5] ,\n16_reg_n_0_[4] ,\n16_reg_n_0_[3] ,\n16_reg_n_0_[2] ,\n16_reg_n_0_[1] ,\n16_reg_n_0_[0] }),
        .O(n202_out),
        .S({n20_carry_i_1_n_0,n20_carry_i_2_n_0,n20_carry_i_3_n_0,n20_carry_i_4_n_0,n20_carry_i_5_n_0,n20_carry_i_6_n_0,n20_carry_i_7_n_0,n20_carry_i_8_n_0}));
  LUT1 #(
    .INIT(2'h1)) 
    n20_carry_i_1
       (.I0(\n16_reg_n_0_[7] ),
        .O(n20_carry_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    n20_carry_i_2
       (.I0(\n16_reg_n_0_[6] ),
        .O(n20_carry_i_2_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    n20_carry_i_3
       (.I0(\n16_reg_n_0_[5] ),
        .O(n20_carry_i_3_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    n20_carry_i_4
       (.I0(\n16_reg_n_0_[4] ),
        .O(n20_carry_i_4_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    n20_carry_i_5
       (.I0(\n16_reg_n_0_[3] ),
        .O(n20_carry_i_5_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    n20_carry_i_6
       (.I0(\n16_reg_n_0_[2] ),
        .O(n20_carry_i_6_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    n20_carry_i_7
       (.I0(\n16_reg_n_0_[1] ),
        .O(n20_carry_i_7_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    n20_carry_i_8
       (.I0(\n16_reg_n_0_[0] ),
        .O(n20_carry_i_8_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[0]),
        .Q(n21[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[1]),
        .Q(n21[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[2]),
        .Q(n21[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[3]),
        .Q(n21[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[4]),
        .Q(n21[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[5]),
        .Q(n21[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[6]),
        .Q(n21[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[7]),
        .Q(n21[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[15]),
        .Q(n22_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__0
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[14]),
        .Q(n22__0_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__1
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[13]),
        .Q(n22__1_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__2
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[12]),
        .Q(n22__2_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__3
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[11]),
        .Q(n22__3_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__4
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[10]),
        .Q(n22__4_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__5
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[9]),
        .Q(n22__5_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__6
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[8]),
        .Q(n22__6_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__17_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__17_carry_n_0,n25__17_carry_n_1,n25__17_carry_n_2,n25__17_carry_n_3,n25__17_carry_n_4,n25__17_carry_n_5,n25__17_carry_n_6,n25__17_carry_n_7}),
        .DI({n25_carry_i_1_n_0,n25__17_carry_i_1_n_0,n25__17_carry_i_2_n_0,n25__17_carry_i_3_n_0,n25__17_carry_i_4_n_0,\n4_reg_n_0_[2] ,\n4_reg_n_0_[1] ,1'b0}),
        .O({n25__17_carry_n_8,n25__17_carry_n_9,n25__17_carry_n_10,n25__17_carry_n_11,n25__17_carry_n_12,n25__17_carry_n_13,n25__17_carry_n_14,NLW_n25__17_carry_O_UNCONNECTED[0]}),
        .S({n25__17_carry_i_5_n_0,n25__17_carry_i_6__1_n_0,n25__17_carry_i_7__1_n_0,n25__17_carry_i_8_n_0,n25__17_carry_i_9__1_n_0,n25__17_carry_i_10_n_0,n25__17_carry_i_11__1_n_0,\n4_reg_n_0_[0] }));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__17_carry__0
       (.CI(n25__17_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__17_carry__0_CO_UNCONNECTED[7:3],n25__17_carry__0_n_5,NLW_n25__17_carry__0_CO_UNCONNECTED[1],n25__17_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25__17_carry__0_i_1__1_n_0,n25__17_carry__0_i_2_n_0}),
        .O({NLW_n25__17_carry__0_O_UNCONNECTED[7:2],n25__17_carry__0_n_14,n25__17_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n25__17_carry__0_i_3__1_n_0,n25__17_carry__0_i_4_n_0}));
  LUT2 #(
    .INIT(4'h2)) 
    n25__17_carry__0_i_1__1
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(n25__17_carry__0_i_1__1_n_0));
  LUT3 #(
    .INIT(8'h8E)) 
    n25__17_carry__0_i_2
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(n25__17_carry__0_i_2_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    n25__17_carry__0_i_3__1
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(n25__17_carry__0_i_3__1_n_0));
  LUT3 #(
    .INIT(8'h4D)) 
    n25__17_carry__0_i_4
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(n25__17_carry__0_i_4_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25__17_carry_i_1
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[5] ),
        .O(n25__17_carry_i_1_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    n25__17_carry_i_10
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[2] ),
        .O(n25__17_carry_i_10_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n25__17_carry_i_11__1
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[0] ),
        .O(n25__17_carry_i_11__1_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25__17_carry_i_2
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[4] ),
        .O(n25__17_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25__17_carry_i_3
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[2] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(n25__17_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    n25__17_carry_i_4
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(n25__17_carry_i_4_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    n25__17_carry_i_5
       (.I0(n25_carry_i_1_n_0),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[5] ),
        .I3(\n4_reg_n_0_[7] ),
        .O(n25__17_carry_i_5_n_0));
  (* HLUTNM = "lutpair88" *) 
  LUT4 #(
    .INIT(16'h781E)) 
    n25__17_carry_i_6__1
       (.I0(\n4_reg_n_0_[4] ),
        .I1(\n4_reg_n_0_[5] ),
        .I2(\n4_reg_n_0_[6] ),
        .I3(\n4_reg_n_0_[3] ),
        .O(n25__17_carry_i_6__1_n_0));
  LUT4 #(
    .INIT(16'h2BD4)) 
    n25__17_carry_i_7__1
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[3] ),
        .I3(\n4_reg_n_0_[5] ),
        .O(n25__17_carry_i_7__1_n_0));
  LUT4 #(
    .INIT(16'h2BD4)) 
    n25__17_carry_i_8
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[2] ),
        .I3(\n4_reg_n_0_[4] ),
        .O(n25__17_carry_i_8_n_0));
  LUT4 #(
    .INIT(16'h6696)) 
    n25__17_carry_i_9__1
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[1] ),
        .I3(\n4_reg_n_0_[0] ),
        .O(n25__17_carry_i_9__1_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__47_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__47_carry_CO_UNCONNECTED[7],n25__47_carry_n_1,n25__47_carry_n_2,n25__47_carry_n_3,n25__47_carry_n_4,n25__47_carry_n_5,n25__47_carry_n_6,n25__47_carry_n_7}),
        .DI({1'b0,\n4_reg_n_0_[6] ,\n4_reg_n_0_[5] ,\n4_reg_n_0_[4] ,\n4_reg_n_0_[3] ,1'b1,1'b0,1'b1}),
        .O({n25__47_carry_n_8,n25__47_carry_n_9,n25__47_carry_n_10,n25__47_carry_n_11,n25__47_carry_n_12,n25__47_carry_n_13,n25__47_carry_n_14,n25__47_carry_n_15}),
        .S({n25__47_carry_i_1_n_0,n25__47_carry_i_2_n_0,n25__47_carry_i_3__1_n_0,n25__47_carry_i_4__1_n_0,n25__47_carry_i_5__1_n_0,\n4_reg_n_0_[3] ,\n4_reg_n_0_[2] ,n25__47_carry_i_6_n_0}));
  LUT1 #(
    .INIT(2'h1)) 
    n25__47_carry_i_1
       (.I0(\n4_reg_n_0_[7] ),
        .O(n25__47_carry_i_1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n25__47_carry_i_2
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(n25__47_carry_i_2_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n25__47_carry_i_3__1
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .O(n25__47_carry_i_3__1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n25__47_carry_i_4__1
       (.I0(\n4_reg_n_0_[4] ),
        .I1(\n4_reg_n_0_[5] ),
        .O(n25__47_carry_i_4__1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n25__47_carry_i_5__1
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[4] ),
        .O(n25__47_carry_i_5__1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    n25__47_carry_i_6
       (.I0(\n4_reg_n_0_[1] ),
        .O(n25__47_carry_i_6_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__67_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__67_carry_n_0,n25__67_carry_n_1,n25__67_carry_n_2,n25__67_carry_n_3,n25__67_carry_n_4,n25__67_carry_n_5,n25__67_carry_n_6,n25__67_carry_n_7}),
        .DI({n25__67_carry_i_1_n_0,n25__67_carry_i_2_n_0,n25__67_carry_i_3_n_0,n25__67_carry_i_4_n_0,n25__67_carry_i_5_n_0,n25__67_carry_i_6_n_0,n25__67_carry_i_7_n_0,1'b0}),
        .O({n26[3:0],NLW_n25__67_carry_O_UNCONNECTED[3:0]}),
        .S({n25__67_carry_i_8_n_0,n25__67_carry_i_9_n_0,n25__67_carry_i_10_n_0,n25__67_carry_i_11_n_0,n25__67_carry_i_12_n_0,n25__67_carry_i_13_n_0,n25__67_carry_i_14_n_0,n25__67_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__67_carry__0
       (.CI(n25__67_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__67_carry__0_CO_UNCONNECTED[7:3],n25__67_carry__0_n_5,n25__67_carry__0_n_6,n25__67_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n25__67_carry__0_i_1_n_0,n25__67_carry__0_i_2_n_0,n25__67_carry__0_i_3_n_0}),
        .O({NLW_n25__67_carry__0_O_UNCONNECTED[7:4],n26[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n25__67_carry__0_i_4_n_0,n25__67_carry__0_i_5_n_0,n25__67_carry__0_i_6_n_0,n25__67_carry__0_i_7_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry__0_i_1
       (.I0(n25__17_carry__0_n_14),
        .I1(n25__47_carry_n_10),
        .O(n25__67_carry__0_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry__0_i_2
       (.I0(n25__17_carry__0_n_15),
        .I1(n25__47_carry_n_11),
        .O(n25__67_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25__67_carry__0_i_3
       (.I0(n25__47_carry_n_12),
        .I1(n25__17_carry_n_8),
        .I2(n25_carry__0_n_5),
        .O(n25__67_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n25__67_carry__0_i_4
       (.I0(n25__17_carry__0_n_5),
        .I1(n25__47_carry_n_9),
        .I2(n25__47_carry_n_8),
        .O(n25__67_carry__0_i_4_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__67_carry__0_i_5
       (.I0(n25__17_carry__0_n_14),
        .I1(n25__47_carry_n_10),
        .I2(n25__47_carry_n_9),
        .I3(n25__17_carry__0_n_5),
        .O(n25__67_carry__0_i_5_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__67_carry__0_i_6
       (.I0(n25__17_carry__0_n_15),
        .I1(n25__47_carry_n_11),
        .I2(n25__47_carry_n_10),
        .I3(n25__17_carry__0_n_14),
        .O(n25__67_carry__0_i_6_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n25__67_carry__0_i_7
       (.I0(n25_carry__0_n_5),
        .I1(n25__17_carry_n_8),
        .I2(n25__47_carry_n_12),
        .I3(n25__47_carry_n_11),
        .I4(n25__17_carry__0_n_15),
        .O(n25__67_carry__0_i_7_n_0));
  (* HLUTNM = "lutpair35" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__67_carry_i_1
       (.I0(n25__47_carry_n_13),
        .I1(n25__17_carry_n_9),
        .I2(n25_carry__0_n_14),
        .O(n25__67_carry_i_1_n_0));
  (* HLUTNM = "lutpair34" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__67_carry_i_10
       (.I0(n25__47_carry_n_14),
        .I1(n25__17_carry_n_10),
        .I2(n25_carry__0_n_15),
        .I3(n25__67_carry_i_3_n_0),
        .O(n25__67_carry_i_10_n_0));
  (* HLUTNM = "lutpair33" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__67_carry_i_11
       (.I0(n25__47_carry_n_15),
        .I1(n25__17_carry_n_11),
        .I2(n25_carry_n_8),
        .I3(n25__67_carry_i_4_n_0),
        .O(n25__67_carry_i_11_n_0));
  (* HLUTNM = "lutpair32" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__67_carry_i_12
       (.I0(n25_carry_n_15),
        .I1(n25__17_carry_n_12),
        .I2(n25_carry_n_9),
        .I3(n25__67_carry_i_5_n_0),
        .O(n25__67_carry_i_12_n_0));
  (* HLUTNM = "lutpair89" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n25__67_carry_i_13
       (.I0(n25__17_carry_n_13),
        .I1(n25_carry_n_10),
        .I2(n25_carry_n_11),
        .I3(n25__17_carry_n_14),
        .O(n25__67_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__67_carry_i_14
       (.I0(n25_carry_n_12),
        .I1(\n4_reg_n_0_[0] ),
        .I2(n25__17_carry_n_14),
        .I3(n25_carry_n_11),
        .O(n25__67_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n25__67_carry_i_15
       (.I0(n25_carry_n_12),
        .I1(\n4_reg_n_0_[0] ),
        .O(n25__67_carry_i_15_n_0));
  (* HLUTNM = "lutpair34" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__67_carry_i_2
       (.I0(n25__47_carry_n_14),
        .I1(n25__17_carry_n_10),
        .I2(n25_carry__0_n_15),
        .O(n25__67_carry_i_2_n_0));
  (* HLUTNM = "lutpair33" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__67_carry_i_3
       (.I0(n25__47_carry_n_15),
        .I1(n25__17_carry_n_11),
        .I2(n25_carry_n_8),
        .O(n25__67_carry_i_3_n_0));
  (* HLUTNM = "lutpair32" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__67_carry_i_4
       (.I0(n25_carry_n_15),
        .I1(n25__17_carry_n_12),
        .I2(n25_carry_n_9),
        .O(n25__67_carry_i_4_n_0));
  (* HLUTNM = "lutpair89" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry_i_5
       (.I0(n25__17_carry_n_13),
        .I1(n25_carry_n_10),
        .O(n25__67_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry_i_6
       (.I0(n25_carry_n_11),
        .I1(n25__17_carry_n_14),
        .O(n25__67_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry_i_7
       (.I0(n25_carry_n_12),
        .I1(\n4_reg_n_0_[0] ),
        .O(n25__67_carry_i_7_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n25__67_carry_i_8
       (.I0(n25__67_carry_i_1_n_0),
        .I1(n25__17_carry_n_8),
        .I2(n25__47_carry_n_12),
        .I3(n25_carry__0_n_5),
        .O(n25__67_carry_i_8_n_0));
  (* HLUTNM = "lutpair35" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__67_carry_i_9
       (.I0(n25__47_carry_n_13),
        .I1(n25__17_carry_n_9),
        .I2(n25_carry__0_n_14),
        .I3(n25__67_carry_i_2_n_0),
        .O(n25__67_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25_carry_n_0,n25_carry_n_1,n25_carry_n_2,n25_carry_n_3,n25_carry_n_4,n25_carry_n_5,n25_carry_n_6,n25_carry_n_7}),
        .DI({n25_carry_i_1_n_0,n25_carry_i_2_n_0,n25_carry_i_3_n_0,n25_carry_i_4_n_0,n25_carry_i_5_n_0,\n4_reg_n_0_[2] ,\n4_reg_n_0_[1] ,1'b0}),
        .O({n25_carry_n_8,n25_carry_n_9,n25_carry_n_10,n25_carry_n_11,n25_carry_n_12,NLW_n25_carry_O_UNCONNECTED[2:1],n25_carry_n_15}),
        .S({n25_carry_i_6_n_0,n25_carry_i_7__1_n_0,n25_carry_i_8__1_n_0,n25_carry_i_9_n_0,n25_carry_i_10_n_0,n25_carry_i_11_n_0,n25_carry_i_12_n_0,\n4_reg_n_0_[0] }));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25_carry__0
       (.CI(n25_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25_carry__0_CO_UNCONNECTED[7:3],n25_carry__0_n_5,NLW_n25_carry__0_CO_UNCONNECTED[1],n25_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25_carry__0_i_1_n_0,n25_carry__0_i_2_n_0}),
        .O({NLW_n25_carry__0_O_UNCONNECTED[7:2],n25_carry__0_n_14,n25_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n25_carry__0_i_3__1_n_0,n25_carry__0_i_4_n_0}));
  LUT2 #(
    .INIT(4'h2)) 
    n25_carry__0_i_1
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(n25_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h8E)) 
    n25_carry__0_i_2
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(n25_carry__0_i_2_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    n25_carry__0_i_3__1
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(n25_carry__0_i_3__1_n_0));
  LUT3 #(
    .INIT(8'h4D)) 
    n25_carry__0_i_4
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(n25_carry__0_i_4_n_0));
  (* HLUTNM = "lutpair88" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25_carry_i_1
       (.I0(\n4_reg_n_0_[4] ),
        .I1(\n4_reg_n_0_[5] ),
        .I2(\n4_reg_n_0_[6] ),
        .O(n25_carry_i_1_n_0));
  LUT4 #(
    .INIT(16'h6696)) 
    n25_carry_i_10
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[1] ),
        .I3(\n4_reg_n_0_[0] ),
        .O(n25_carry_i_10_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    n25_carry_i_11
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[2] ),
        .O(n25_carry_i_11_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n25_carry_i_12
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[0] ),
        .O(n25_carry_i_12_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25_carry_i_2
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[5] ),
        .O(n25_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25_carry_i_3
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[4] ),
        .O(n25_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25_carry_i_4
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[2] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(n25_carry_i_4_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    n25_carry_i_5
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(n25_carry_i_5_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    n25_carry_i_6
       (.I0(n25_carry_i_1_n_0),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[5] ),
        .I3(\n4_reg_n_0_[7] ),
        .O(n25_carry_i_6_n_0));
  LUT4 #(
    .INIT(16'h2BD4)) 
    n25_carry_i_7__1
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[5] ),
        .I2(\n4_reg_n_0_[4] ),
        .I3(\n4_reg_n_0_[6] ),
        .O(n25_carry_i_7__1_n_0));
  LUT4 #(
    .INIT(16'h2BD4)) 
    n25_carry_i_8__1
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[3] ),
        .I3(\n4_reg_n_0_[5] ),
        .O(n25_carry_i_8__1_n_0));
  LUT4 #(
    .INIT(16'h2BD4)) 
    n25_carry_i_9
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[2] ),
        .I3(\n4_reg_n_0_[4] ),
        .O(n25_carry_i_9_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[0]),
        .Q(n27[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[1]),
        .Q(n27[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[2]),
        .Q(n27[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[3]),
        .Q(n27[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[4]),
        .Q(n27[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[5]),
        .Q(n27[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[6]),
        .Q(n27[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[7]),
        .Q(n27[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[0]),
        .Q(n29[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[1]),
        .Q(n29[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[2]),
        .Q(n29[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[3]),
        .Q(n29[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[4]),
        .Q(n29[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[5]),
        .Q(n29[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[6]),
        .Q(n29[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[7]),
        .Q(n29[7]),
        .R(rst_i));
  LUT2 #(
    .INIT(4'h6)) 
    \n33[0]_i_1__2 
       (.I0(n29[0]),
        .I1(n10[0]),
        .O(n31[0]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[10]_i_1__2 
       (.I0(n21[2]),
        .I1(\n8_reg_n_0_[2] ),
        .I2(\n8_reg_n_0_[1] ),
        .I3(n21[1]),
        .I4(\n8_reg_n_0_[0] ),
        .I5(n21[0]),
        .O(\n33[10]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[11]_i_1__2 
       (.I0(n21[3]),
        .I1(\n8_reg_n_0_[3] ),
        .I2(\n33[12]_i_2__2_n_0 ),
        .O(\n33[11]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[12]_i_1__2 
       (.I0(n21[4]),
        .I1(\n8_reg_n_0_[4] ),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[3]),
        .I4(\n33[12]_i_2__2_n_0 ),
        .O(\n33[12]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[12]_i_2__2 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n33[12]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[13]_i_1__2 
       (.I0(n21[5]),
        .I1(\n8_reg_n_0_[5] ),
        .I2(\n33[14]_i_2__2_n_0 ),
        .O(\n33[13]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[14]_i_1__2 
       (.I0(n21[6]),
        .I1(\n8_reg_n_0_[6] ),
        .I2(\n8_reg_n_0_[5] ),
        .I3(n21[5]),
        .I4(\n33[14]_i_2__2_n_0 ),
        .O(\n33[14]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[14]_i_2__2 
       (.I0(\n33[12]_i_2__2_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n33[14]_i_2__2_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[15]_i_1__2 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n33[15]_i_2__2_n_0 ),
        .O(n30[7]));
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[15]_i_2__2 
       (.I0(\n33[14]_i_2__2_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n33[15]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[1]_i_1__2 
       (.I0(n29[1]),
        .I1(n10[1]),
        .I2(n10[0]),
        .I3(n29[0]),
        .O(n31[1]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[2]_i_1__2 
       (.I0(n29[2]),
        .I1(n10[2]),
        .I2(n10[1]),
        .I3(n29[1]),
        .I4(n10[0]),
        .I5(n29[0]),
        .O(\n33[2]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[3]_i_1__2 
       (.I0(n29[3]),
        .I1(n10[3]),
        .I2(\n33[4]_i_2__2_n_0 ),
        .O(\n33[3]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[4]_i_1__2 
       (.I0(n29[4]),
        .I1(n10[4]),
        .I2(n10[3]),
        .I3(n29[3]),
        .I4(\n33[4]_i_2__2_n_0 ),
        .O(\n33[4]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[4]_i_2__2 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n33[4]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[5]_i_1__2 
       (.I0(n29[5]),
        .I1(n10[5]),
        .I2(\n33[6]_i_2__2_n_0 ),
        .O(\n33[5]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[6]_i_1__2 
       (.I0(n29[6]),
        .I1(n10[6]),
        .I2(n10[5]),
        .I3(n29[5]),
        .I4(\n33[6]_i_2__2_n_0 ),
        .O(\n33[6]_i_1__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[6]_i_2__2 
       (.I0(\n33[4]_i_2__2_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n33[6]_i_2__2_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[7]_i_1__2 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n33[7]_i_2__2_n_0 ),
        .O(n31[7]));
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[7]_i_2__2 
       (.I0(\n33[6]_i_2__2_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n33[7]_i_2__2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n33[8]_i_1__1 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .O(n30[0]));
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[9]_i_1__2 
       (.I0(n21[1]),
        .I1(\n8_reg_n_0_[1] ),
        .I2(\n8_reg_n_0_[0] ),
        .I3(n21[0]),
        .O(\n33[9]_i_1__2_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[0]),
        .Q(i1[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[10]_i_1__2_n_0 ),
        .Q(i1[24]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[11]_i_1__2_n_0 ),
        .Q(i1[25]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[12]_i_1__2_n_0 ),
        .Q(i1[26]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[13]_i_1__2_n_0 ),
        .Q(i1[27]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[14]_i_1__2_n_0 ),
        .Q(i1[28]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n30[7]),
        .Q(i1[29]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[1]),
        .Q(i1[15]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[2]_i_1__2_n_0 ),
        .Q(i1[16]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[3]_i_1__2_n_0 ),
        .Q(i1[17]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[4]_i_1__2_n_0 ),
        .Q(i1[18]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[5]_i_1__2_n_0 ),
        .Q(i1[19]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[6]_i_1__2_n_0 ),
        .Q(i1[20]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[7]),
        .Q(i1[21]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n30[0]),
        .Q(i1[22]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[9]_i_1__2_n_0 ),
        .Q(i1[23]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[10]_i_1__2 
       (.I0(\n8_reg_n_0_[1] ),
        .I1(n21[1]),
        .I2(n21[0]),
        .I3(\n8_reg_n_0_[0] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(n341_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[11]_i_1__2 
       (.I0(\n37[12]_i_2__2_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .O(n341_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[12]_i_1__2 
       (.I0(\n8_reg_n_0_[3] ),
        .I1(n21[3]),
        .I2(\n37[12]_i_2__2_n_0 ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(n341_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[12]_i_2__2 
       (.I0(\n8_reg_n_0_[0] ),
        .I1(n21[0]),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n37[12]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[13]_i_1__2 
       (.I0(\n37[14]_i_2__2_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(n341_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[14]_i_1__2 
       (.I0(\n8_reg_n_0_[5] ),
        .I1(n21[5]),
        .I2(\n37[14]_i_2__2_n_0 ),
        .I3(n21[6]),
        .I4(\n8_reg_n_0_[6] ),
        .O(n341_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[14]_i_2__2 
       (.I0(\n37[12]_i_2__2_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n37[14]_i_2__2_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[15]_i_1__2 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n37[15]_i_2__2_n_0 ),
        .O(n341_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[15]_i_2__2 
       (.I0(\n37[14]_i_2__2_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n37[15]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[1]_i_1__2 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .O(n350_out[1]));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[2]_i_1__2 
       (.I0(n10[1]),
        .I1(n29[1]),
        .I2(n29[0]),
        .I3(n10[0]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(n350_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[3]_i_1__2 
       (.I0(\n37[4]_i_2__2_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .O(n350_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[4]_i_1__2 
       (.I0(n10[3]),
        .I1(n29[3]),
        .I2(\n37[4]_i_2__2_n_0 ),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(n350_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[4]_i_2__2 
       (.I0(n10[0]),
        .I1(n29[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n37[4]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[5]_i_1__2 
       (.I0(\n37[6]_i_2__2_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(n350_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[6]_i_1__2 
       (.I0(n10[5]),
        .I1(n29[5]),
        .I2(\n37[6]_i_2__2_n_0 ),
        .I3(n29[6]),
        .I4(n10[6]),
        .O(n350_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[6]_i_2__2 
       (.I0(\n37[4]_i_2__2_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n37[6]_i_2__2_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[7]_i_1__2 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n37[7]_i_2__2_n_0 ),
        .O(n350_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[7]_i_2__2 
       (.I0(\n37[6]_i_2__2_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n37[7]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[9]_i_1__2 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .O(n341_out[1]));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[2]),
        .Q(i1[9]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[3]),
        .Q(i1[10]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[4]),
        .Q(i1[11]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[5]),
        .Q(i1[12]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[6]),
        .Q(i1[13]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[7]),
        .Q(i1[14]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[1]),
        .Q(i1[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[2]),
        .Q(i1[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[3]),
        .Q(i1[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[4]),
        .Q(i1[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[5]),
        .Q(i1[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[6]),
        .Q(i1[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[7]),
        .Q(i1[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[1]),
        .Q(i1[8]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[0]),
        .Q(\n4_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[1]),
        .Q(\n4_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[2]),
        .Q(\n4_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[3]),
        .Q(\n4_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[4]),
        .Q(\n4_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[5]),
        .Q(\n4_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[6]),
        .Q(\n4_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s5_3[7]),
        .Q(\n4_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[0]),
        .Q(\n7_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[1]),
        .Q(\n7_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[2]),
        .Q(\n7_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[3]),
        .Q(\n7_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[4]),
        .Q(\n7_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[5]),
        .Q(\n7_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[6]),
        .Q(\n7_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[7]),
        .Q(\n7_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[0] ),
        .Q(\n8_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[1] ),
        .Q(\n8_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[2] ),
        .Q(\n8_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[3] ),
        .Q(\n8_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[4] ),
        .Q(\n8_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[5] ),
        .Q(\n8_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[6] ),
        .Q(\n8_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[7] ),
        .Q(\n8_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[0] ),
        .Q(\n9_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[1] ),
        .Q(\n9_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[2] ),
        .Q(\n9_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[3] ),
        .Q(\n9_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[4] ),
        .Q(\n9_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[5] ),
        .Q(\n9_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[6] ),
        .Q(\n9_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[7] ),
        .Q(\n9_reg_n_0_[7] ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_15" *) 
module switch_elements_cf_fft_512_8_15
   (\n9_reg[0] ,
    s3_3,
    rst_i,
    enable_i,
    clk_i,
    n14__56_carry,
    s4_3,
    D);
  output [15:0]\n9_reg[0] ;
  output [15:0]s3_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]n14__56_carry;
  input [15:0]s4_3;
  input [15:0]D;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire [15:0]n14__56_carry;
  wire [15:0]n33;
  wire [15:1]n37;
  wire n4;
  wire [15:0]\n9_reg[0] ;
  wire rst_i;
  wire s29_n_0;
  wire [15:0]s3_3;
  wire [15:0]s4_3;

  switch_elements_cf_fft_512_8_31_13 s25
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i8(i8),
        .n4(n4),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_16 s26
       (.D(D),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:1],n37[15:9],n37[7:1],n33[0]}),
        .n14__56_carry_0(n14__56_carry),
        .rst_i(rst_i),
        .s4_3(s4_3));
  switch_elements_cf_fft_512_8_26_14 s28
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:1],n37[15:9],n37[7:1],n33[0]}),
        .i8(i8),
        .\n1_reg[0] (s29_n_0),
        .n4(n4),
        .\n9_reg[0] (\n9_reg[0] ),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_27_15 s29
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:1],n37[15:9],n37[7:1],n33[0]}),
        .i8(i8),
        .\n9_reg[0]_0 (s29_n_0),
        .rst_i(rst_i),
        .s3_3(s3_3));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_16" *) 
module switch_elements_cf_fft_512_8_16
   (i1,
    rst_i,
    enable_i,
    clk_i,
    n14__56_carry_0,
    s4_3,
    D);
  output [29:0]i1;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]n14__56_carry_0;
  input [15:0]s4_3;
  input [15:0]D;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [7:0]n10;
  wire n14__0_carry__0_i_1__1_n_0;
  wire n14__0_carry__0_i_2__1_n_0;
  wire n14__0_carry__0_i_3__1_n_0;
  wire n14__0_carry__0_i_4__1_n_0;
  wire n14__0_carry__0_n_14;
  wire n14__0_carry__0_n_15;
  wire n14__0_carry__0_n_5;
  wire n14__0_carry__0_n_7;
  wire n14__0_carry_i_10__1_n_0;
  wire n14__0_carry_i_11__1_n_0;
  wire n14__0_carry_i_12__1_n_0;
  wire n14__0_carry_i_13__1_n_0;
  wire n14__0_carry_i_14__1_n_0;
  wire n14__0_carry_i_15__1_n_0;
  wire n14__0_carry_i_16__1_n_0;
  wire n14__0_carry_i_17__1_n_0;
  wire n14__0_carry_i_18__1_n_0;
  wire n14__0_carry_i_19__1_n_0;
  wire n14__0_carry_i_1__1_n_0;
  wire n14__0_carry_i_20__1_n_0;
  wire n14__0_carry_i_2__1_n_0;
  wire n14__0_carry_i_3__1_n_0;
  wire n14__0_carry_i_4__1_n_0;
  wire n14__0_carry_i_5__1_n_0;
  wire n14__0_carry_i_6__1_n_0;
  wire n14__0_carry_i_7__1_n_0;
  wire n14__0_carry_i_8__1_n_0;
  wire n14__0_carry_i_9__1_n_0;
  wire n14__0_carry_n_0;
  wire n14__0_carry_n_1;
  wire n14__0_carry_n_10;
  wire n14__0_carry_n_11;
  wire n14__0_carry_n_12;
  wire n14__0_carry_n_2;
  wire n14__0_carry_n_3;
  wire n14__0_carry_n_4;
  wire n14__0_carry_n_5;
  wire n14__0_carry_n_6;
  wire n14__0_carry_n_7;
  wire n14__0_carry_n_8;
  wire n14__0_carry_n_9;
  wire n14__27_carry__0_i_1__1_n_0;
  wire n14__27_carry__0_i_2__1_n_0;
  wire n14__27_carry__0_i_3__1_n_0;
  wire n14__27_carry__0_i_4__1_n_0;
  wire n14__27_carry__0_n_14;
  wire n14__27_carry__0_n_15;
  wire n14__27_carry__0_n_5;
  wire n14__27_carry__0_n_7;
  wire n14__27_carry_i_10__1_n_0;
  wire n14__27_carry_i_11__1_n_0;
  wire n14__27_carry_i_12__1_n_0;
  wire n14__27_carry_i_13__1_n_0;
  wire n14__27_carry_i_14__1_n_0;
  wire n14__27_carry_i_15__1_n_0;
  wire n14__27_carry_i_16__1_n_0;
  wire n14__27_carry_i_17__1_n_0;
  wire n14__27_carry_i_18__1_n_0;
  wire n14__27_carry_i_19__1_n_0;
  wire n14__27_carry_i_1__1_n_0;
  wire n14__27_carry_i_20__1_n_0;
  wire n14__27_carry_i_2__1_n_0;
  wire n14__27_carry_i_3__1_n_0;
  wire n14__27_carry_i_4__1_n_0;
  wire n14__27_carry_i_5__1_n_0;
  wire n14__27_carry_i_6__1_n_0;
  wire n14__27_carry_i_7__1_n_0;
  wire n14__27_carry_i_8__1_n_0;
  wire n14__27_carry_i_9__1_n_0;
  wire n14__27_carry_n_0;
  wire n14__27_carry_n_1;
  wire n14__27_carry_n_10;
  wire n14__27_carry_n_11;
  wire n14__27_carry_n_12;
  wire n14__27_carry_n_13;
  wire n14__27_carry_n_14;
  wire n14__27_carry_n_15;
  wire n14__27_carry_n_2;
  wire n14__27_carry_n_3;
  wire n14__27_carry_n_4;
  wire n14__27_carry_n_5;
  wire n14__27_carry_n_6;
  wire n14__27_carry_n_7;
  wire n14__27_carry_n_8;
  wire n14__27_carry_n_9;
  wire [15:0]n14__56_carry_0;
  wire n14__56_carry__0_i_1__1_n_0;
  wire n14__56_carry__0_n_15;
  wire n14__56_carry_i_10__1_n_0;
  wire n14__56_carry_i_11__1_n_0;
  wire n14__56_carry_i_12__1_n_0;
  wire n14__56_carry_i_13__1_n_0;
  wire n14__56_carry_i_14__1_n_0;
  wire n14__56_carry_i_15__1_n_0;
  wire n14__56_carry_i_1__1_n_0;
  wire n14__56_carry_i_2__1_n_0;
  wire n14__56_carry_i_3__1_n_0;
  wire n14__56_carry_i_4__1_n_0;
  wire n14__56_carry_i_5__1_n_0;
  wire n14__56_carry_i_6__1_n_0;
  wire n14__56_carry_i_7__1_n_0;
  wire n14__56_carry_i_8__1_n_0;
  wire n14__56_carry_i_9__1_n_0;
  wire n14__56_carry_n_0;
  wire n14__56_carry_n_1;
  wire n14__56_carry_n_10;
  wire n14__56_carry_n_11;
  wire n14__56_carry_n_12;
  wire n14__56_carry_n_13;
  wire n14__56_carry_n_14;
  wire n14__56_carry_n_15;
  wire n14__56_carry_n_2;
  wire n14__56_carry_n_3;
  wire n14__56_carry_n_4;
  wire n14__56_carry_n_5;
  wire n14__56_carry_n_6;
  wire n14__56_carry_n_7;
  wire n14__56_carry_n_8;
  wire n14__56_carry_n_9;
  wire n14__81_carry__0_i_1__1_n_0;
  wire n14__81_carry__0_i_2__1_n_0;
  wire n14__81_carry__0_i_3__1_n_0;
  wire n14__81_carry__0_i_4__1_n_0;
  wire n14__81_carry__0_i_5__1_n_0;
  wire n14__81_carry__0_i_6__1_n_0;
  wire n14__81_carry__0_i_7__1_n_0;
  wire n14__81_carry__0_n_5;
  wire n14__81_carry__0_n_6;
  wire n14__81_carry__0_n_7;
  wire n14__81_carry_i_10__1_n_0;
  wire n14__81_carry_i_11__1_n_0;
  wire n14__81_carry_i_12__1_n_0;
  wire n14__81_carry_i_13__1_n_0;
  wire n14__81_carry_i_14__1_n_0;
  wire n14__81_carry_i_15__1_n_0;
  wire n14__81_carry_i_1__1_n_0;
  wire n14__81_carry_i_2__1_n_0;
  wire n14__81_carry_i_3__1_n_0;
  wire n14__81_carry_i_4__1_n_0;
  wire n14__81_carry_i_5__1_n_0;
  wire n14__81_carry_i_6__1_n_0;
  wire n14__81_carry_i_7__1_n_0;
  wire n14__81_carry_i_8__1_n_0;
  wire n14__81_carry_i_9__1_n_0;
  wire n14__81_carry_n_0;
  wire n14__81_carry_n_1;
  wire n14__81_carry_n_2;
  wire n14__81_carry_n_3;
  wire n14__81_carry_n_4;
  wire n14__81_carry_n_5;
  wire n14__81_carry_n_6;
  wire n14__81_carry_n_7;
  wire [7:0]n15;
  wire \n16_reg_n_0_[0] ;
  wire \n16_reg_n_0_[1] ;
  wire \n16_reg_n_0_[2] ;
  wire \n16_reg_n_0_[3] ;
  wire \n16_reg_n_0_[4] ;
  wire \n16_reg_n_0_[5] ;
  wire \n16_reg_n_0_[6] ;
  wire \n16_reg_n_0_[7] ;
  wire [14:7]n17;
  wire n17__0_carry__0_i_1__1_n_0;
  wire n17__0_carry__0_i_2__1_n_0;
  wire n17__0_carry__0_i_3__1_n_0;
  wire n17__0_carry__0_i_4__1_n_0;
  wire n17__0_carry__0_n_14;
  wire n17__0_carry__0_n_15;
  wire n17__0_carry__0_n_5;
  wire n17__0_carry__0_n_7;
  wire n17__0_carry_i_10__1_n_0;
  wire n17__0_carry_i_11__1_n_0;
  wire n17__0_carry_i_12__1_n_0;
  wire n17__0_carry_i_13__1_n_0;
  wire n17__0_carry_i_14__1_n_0;
  wire n17__0_carry_i_15__1_n_0;
  wire n17__0_carry_i_16__1_n_0;
  wire n17__0_carry_i_17__1_n_0;
  wire n17__0_carry_i_18__1_n_0;
  wire n17__0_carry_i_19__1_n_0;
  wire n17__0_carry_i_1__1_n_0;
  wire n17__0_carry_i_20__1_n_0;
  wire n17__0_carry_i_2__1_n_0;
  wire n17__0_carry_i_3__1_n_0;
  wire n17__0_carry_i_4__1_n_0;
  wire n17__0_carry_i_5__1_n_0;
  wire n17__0_carry_i_6__1_n_0;
  wire n17__0_carry_i_7__1_n_0;
  wire n17__0_carry_i_8__1_n_0;
  wire n17__0_carry_i_9__1_n_0;
  wire n17__0_carry_n_0;
  wire n17__0_carry_n_1;
  wire n17__0_carry_n_10;
  wire n17__0_carry_n_11;
  wire n17__0_carry_n_12;
  wire n17__0_carry_n_2;
  wire n17__0_carry_n_3;
  wire n17__0_carry_n_4;
  wire n17__0_carry_n_5;
  wire n17__0_carry_n_6;
  wire n17__0_carry_n_7;
  wire n17__0_carry_n_8;
  wire n17__0_carry_n_9;
  wire n17__27_carry__0_i_1__1_n_0;
  wire n17__27_carry__0_i_2__1_n_0;
  wire n17__27_carry__0_i_3__1_n_0;
  wire n17__27_carry__0_i_4__1_n_0;
  wire n17__27_carry__0_n_14;
  wire n17__27_carry__0_n_15;
  wire n17__27_carry__0_n_5;
  wire n17__27_carry__0_n_7;
  wire n17__27_carry_i_10__1_n_0;
  wire n17__27_carry_i_11__1_n_0;
  wire n17__27_carry_i_12__1_n_0;
  wire n17__27_carry_i_13__1_n_0;
  wire n17__27_carry_i_14__1_n_0;
  wire n17__27_carry_i_15__1_n_0;
  wire n17__27_carry_i_16__1_n_0;
  wire n17__27_carry_i_17__1_n_0;
  wire n17__27_carry_i_18__1_n_0;
  wire n17__27_carry_i_19__1_n_0;
  wire n17__27_carry_i_1__1_n_0;
  wire n17__27_carry_i_20__1_n_0;
  wire n17__27_carry_i_2__1_n_0;
  wire n17__27_carry_i_3__1_n_0;
  wire n17__27_carry_i_4__1_n_0;
  wire n17__27_carry_i_5__1_n_0;
  wire n17__27_carry_i_6__1_n_0;
  wire n17__27_carry_i_7__1_n_0;
  wire n17__27_carry_i_8__1_n_0;
  wire n17__27_carry_i_9__1_n_0;
  wire n17__27_carry_n_0;
  wire n17__27_carry_n_1;
  wire n17__27_carry_n_10;
  wire n17__27_carry_n_11;
  wire n17__27_carry_n_12;
  wire n17__27_carry_n_13;
  wire n17__27_carry_n_14;
  wire n17__27_carry_n_15;
  wire n17__27_carry_n_2;
  wire n17__27_carry_n_3;
  wire n17__27_carry_n_4;
  wire n17__27_carry_n_5;
  wire n17__27_carry_n_6;
  wire n17__27_carry_n_7;
  wire n17__27_carry_n_8;
  wire n17__27_carry_n_9;
  wire n17__56_carry__0_i_1__1_n_0;
  wire n17__56_carry__0_n_15;
  wire n17__56_carry_i_10__1_n_0;
  wire n17__56_carry_i_11__1_n_0;
  wire n17__56_carry_i_12__1_n_0;
  wire n17__56_carry_i_13__1_n_0;
  wire n17__56_carry_i_14__1_n_0;
  wire n17__56_carry_i_15__1_n_0;
  wire n17__56_carry_i_1__1_n_0;
  wire n17__56_carry_i_2__1_n_0;
  wire n17__56_carry_i_3__1_n_0;
  wire n17__56_carry_i_4__1_n_0;
  wire n17__56_carry_i_5__1_n_0;
  wire n17__56_carry_i_6__1_n_0;
  wire n17__56_carry_i_7__1_n_0;
  wire n17__56_carry_i_8__1_n_0;
  wire n17__56_carry_i_9__1_n_0;
  wire n17__56_carry_n_0;
  wire n17__56_carry_n_1;
  wire n17__56_carry_n_10;
  wire n17__56_carry_n_11;
  wire n17__56_carry_n_12;
  wire n17__56_carry_n_13;
  wire n17__56_carry_n_14;
  wire n17__56_carry_n_15;
  wire n17__56_carry_n_2;
  wire n17__56_carry_n_3;
  wire n17__56_carry_n_4;
  wire n17__56_carry_n_5;
  wire n17__56_carry_n_6;
  wire n17__56_carry_n_7;
  wire n17__56_carry_n_8;
  wire n17__56_carry_n_9;
  wire n17__81_carry__0_i_1__1_n_0;
  wire n17__81_carry__0_i_2__1_n_0;
  wire n17__81_carry__0_i_3__1_n_0;
  wire n17__81_carry__0_i_4__1_n_0;
  wire n17__81_carry__0_i_5__1_n_0;
  wire n17__81_carry__0_i_6__1_n_0;
  wire n17__81_carry__0_i_7__1_n_0;
  wire n17__81_carry__0_n_5;
  wire n17__81_carry__0_n_6;
  wire n17__81_carry__0_n_7;
  wire n17__81_carry_i_10__1_n_0;
  wire n17__81_carry_i_11__1_n_0;
  wire n17__81_carry_i_12__1_n_0;
  wire n17__81_carry_i_13__1_n_0;
  wire n17__81_carry_i_14__1_n_0;
  wire n17__81_carry_i_15__1_n_0;
  wire n17__81_carry_i_1__1_n_0;
  wire n17__81_carry_i_2__1_n_0;
  wire n17__81_carry_i_3__1_n_0;
  wire n17__81_carry_i_4__1_n_0;
  wire n17__81_carry_i_5__1_n_0;
  wire n17__81_carry_i_6__1_n_0;
  wire n17__81_carry_i_7__1_n_0;
  wire n17__81_carry_i_8__1_n_0;
  wire n17__81_carry_i_9__1_n_0;
  wire n17__81_carry_n_0;
  wire n17__81_carry_n_1;
  wire n17__81_carry_n_2;
  wire n17__81_carry_n_3;
  wire n17__81_carry_n_4;
  wire n17__81_carry_n_5;
  wire n17__81_carry_n_6;
  wire n17__81_carry_n_7;
  wire n19_reg__0_n_0;
  wire n19_reg__1_n_0;
  wire n19_reg__2_n_0;
  wire n19_reg__3_n_0;
  wire n19_reg__4_n_0;
  wire n19_reg__5_n_0;
  wire n19_reg__6_n_0;
  wire n19_reg_n_0;
  wire \n1_reg_n_0_[0] ;
  wire \n1_reg_n_0_[1] ;
  wire \n1_reg_n_0_[2] ;
  wire \n1_reg_n_0_[3] ;
  wire \n1_reg_n_0_[4] ;
  wire \n1_reg_n_0_[5] ;
  wire \n1_reg_n_0_[6] ;
  wire \n1_reg_n_0_[7] ;
  wire [7:0]n2;
  wire [7:0]n202_out;
  wire n20_carry_i_1__2_n_0;
  wire n20_carry_i_2__2_n_0;
  wire n20_carry_i_3__2_n_0;
  wire n20_carry_i_4__2_n_0;
  wire n20_carry_i_5__2_n_0;
  wire n20_carry_i_6__2_n_0;
  wire n20_carry_i_7__2_n_0;
  wire n20_carry_i_8__2_n_0;
  wire n20_carry_n_1;
  wire n20_carry_n_2;
  wire n20_carry_n_3;
  wire n20_carry_n_4;
  wire n20_carry_n_5;
  wire n20_carry_n_6;
  wire n20_carry_n_7;
  wire [7:0]n21;
  wire n22__0_carry__0_i_1__1_n_0;
  wire n22__0_carry__0_i_2__1_n_0;
  wire n22__0_carry__0_i_3__1_n_0;
  wire n22__0_carry__0_i_4__1_n_0;
  wire n22__0_carry__0_n_14;
  wire n22__0_carry__0_n_15;
  wire n22__0_carry__0_n_5;
  wire n22__0_carry__0_n_7;
  wire n22__0_carry_i_10__1_n_0;
  wire n22__0_carry_i_11__1_n_0;
  wire n22__0_carry_i_12__1_n_0;
  wire n22__0_carry_i_13__1_n_0;
  wire n22__0_carry_i_14__1_n_0;
  wire n22__0_carry_i_15__1_n_0;
  wire n22__0_carry_i_16__1_n_0;
  wire n22__0_carry_i_17__1_n_0;
  wire n22__0_carry_i_18__1_n_0;
  wire n22__0_carry_i_19__1_n_0;
  wire n22__0_carry_i_1__1_n_0;
  wire n22__0_carry_i_20__1_n_0;
  wire n22__0_carry_i_2__1_n_0;
  wire n22__0_carry_i_3__1_n_0;
  wire n22__0_carry_i_4__1_n_0;
  wire n22__0_carry_i_5__1_n_0;
  wire n22__0_carry_i_6__1_n_0;
  wire n22__0_carry_i_7__1_n_0;
  wire n22__0_carry_i_8__1_n_0;
  wire n22__0_carry_i_9__1_n_0;
  wire n22__0_carry_n_0;
  wire n22__0_carry_n_1;
  wire n22__0_carry_n_10;
  wire n22__0_carry_n_11;
  wire n22__0_carry_n_12;
  wire n22__0_carry_n_2;
  wire n22__0_carry_n_3;
  wire n22__0_carry_n_4;
  wire n22__0_carry_n_5;
  wire n22__0_carry_n_6;
  wire n22__0_carry_n_7;
  wire n22__0_carry_n_8;
  wire n22__0_carry_n_9;
  wire n22__0_n_0;
  wire n22__1_n_0;
  wire n22__27_carry__0_i_1__1_n_0;
  wire n22__27_carry__0_i_2__1_n_0;
  wire n22__27_carry__0_i_3__1_n_0;
  wire n22__27_carry__0_i_4__1_n_0;
  wire n22__27_carry__0_n_14;
  wire n22__27_carry__0_n_15;
  wire n22__27_carry__0_n_5;
  wire n22__27_carry__0_n_7;
  wire n22__27_carry_i_10__1_n_0;
  wire n22__27_carry_i_11__1_n_0;
  wire n22__27_carry_i_12__1_n_0;
  wire n22__27_carry_i_13__1_n_0;
  wire n22__27_carry_i_14__1_n_0;
  wire n22__27_carry_i_15__1_n_0;
  wire n22__27_carry_i_16__1_n_0;
  wire n22__27_carry_i_17__1_n_0;
  wire n22__27_carry_i_18__1_n_0;
  wire n22__27_carry_i_19__1_n_0;
  wire n22__27_carry_i_1__1_n_0;
  wire n22__27_carry_i_20__1_n_0;
  wire n22__27_carry_i_2__1_n_0;
  wire n22__27_carry_i_3__1_n_0;
  wire n22__27_carry_i_4__1_n_0;
  wire n22__27_carry_i_5__1_n_0;
  wire n22__27_carry_i_6__1_n_0;
  wire n22__27_carry_i_7__1_n_0;
  wire n22__27_carry_i_8__1_n_0;
  wire n22__27_carry_i_9__1_n_0;
  wire n22__27_carry_n_0;
  wire n22__27_carry_n_1;
  wire n22__27_carry_n_10;
  wire n22__27_carry_n_11;
  wire n22__27_carry_n_12;
  wire n22__27_carry_n_13;
  wire n22__27_carry_n_14;
  wire n22__27_carry_n_15;
  wire n22__27_carry_n_2;
  wire n22__27_carry_n_3;
  wire n22__27_carry_n_4;
  wire n22__27_carry_n_5;
  wire n22__27_carry_n_6;
  wire n22__27_carry_n_7;
  wire n22__27_carry_n_8;
  wire n22__27_carry_n_9;
  wire n22__2_n_0;
  wire n22__3_n_0;
  wire n22__4_n_0;
  wire n22__56_carry__0_i_1__1_n_0;
  wire n22__56_carry__0_n_15;
  wire n22__56_carry_i_10__1_n_0;
  wire n22__56_carry_i_11__1_n_0;
  wire n22__56_carry_i_12__1_n_0;
  wire n22__56_carry_i_13__1_n_0;
  wire n22__56_carry_i_14__1_n_0;
  wire n22__56_carry_i_15__1_n_0;
  wire n22__56_carry_i_1__1_n_0;
  wire n22__56_carry_i_2__1_n_0;
  wire n22__56_carry_i_3__1_n_0;
  wire n22__56_carry_i_4__1_n_0;
  wire n22__56_carry_i_5__1_n_0;
  wire n22__56_carry_i_6__1_n_0;
  wire n22__56_carry_i_7__1_n_0;
  wire n22__56_carry_i_8__1_n_0;
  wire n22__56_carry_i_9__1_n_0;
  wire n22__56_carry_n_0;
  wire n22__56_carry_n_1;
  wire n22__56_carry_n_10;
  wire n22__56_carry_n_11;
  wire n22__56_carry_n_12;
  wire n22__56_carry_n_13;
  wire n22__56_carry_n_14;
  wire n22__56_carry_n_15;
  wire n22__56_carry_n_2;
  wire n22__56_carry_n_3;
  wire n22__56_carry_n_4;
  wire n22__56_carry_n_5;
  wire n22__56_carry_n_6;
  wire n22__56_carry_n_7;
  wire n22__56_carry_n_8;
  wire n22__56_carry_n_9;
  wire n22__5_n_0;
  wire n22__6_n_0;
  wire n22__81_carry__0_i_1__1_n_0;
  wire n22__81_carry__0_i_2__1_n_0;
  wire n22__81_carry__0_i_3__1_n_0;
  wire n22__81_carry__0_i_4__1_n_0;
  wire n22__81_carry__0_i_5__1_n_0;
  wire n22__81_carry__0_i_6__1_n_0;
  wire n22__81_carry__0_i_7__1_n_0;
  wire n22__81_carry__0_n_5;
  wire n22__81_carry__0_n_6;
  wire n22__81_carry__0_n_7;
  wire n22__81_carry_i_10__1_n_0;
  wire n22__81_carry_i_11__1_n_0;
  wire n22__81_carry_i_12__1_n_0;
  wire n22__81_carry_i_13__1_n_0;
  wire n22__81_carry_i_14__1_n_0;
  wire n22__81_carry_i_15__1_n_0;
  wire n22__81_carry_i_1__1_n_0;
  wire n22__81_carry_i_2__1_n_0;
  wire n22__81_carry_i_3__1_n_0;
  wire n22__81_carry_i_4__1_n_0;
  wire n22__81_carry_i_5__1_n_0;
  wire n22__81_carry_i_6__1_n_0;
  wire n22__81_carry_i_7__1_n_0;
  wire n22__81_carry_i_8__1_n_0;
  wire n22__81_carry_i_9__1_n_0;
  wire n22__81_carry_n_0;
  wire n22__81_carry_n_1;
  wire n22__81_carry_n_2;
  wire n22__81_carry_n_3;
  wire n22__81_carry_n_4;
  wire n22__81_carry_n_5;
  wire n22__81_carry_n_6;
  wire n22__81_carry_n_7;
  wire n22_n_0;
  wire [7:0]n23;
  wire [7:0]n24;
  wire n25__0_carry__0_i_1__1_n_0;
  wire n25__0_carry__0_i_2__1_n_0;
  wire n25__0_carry__0_i_3__1_n_0;
  wire n25__0_carry__0_i_4__1_n_0;
  wire n25__0_carry__0_n_14;
  wire n25__0_carry__0_n_15;
  wire n25__0_carry__0_n_5;
  wire n25__0_carry__0_n_7;
  wire n25__0_carry_i_10__1_n_0;
  wire n25__0_carry_i_11__1_n_0;
  wire n25__0_carry_i_12__1_n_0;
  wire n25__0_carry_i_13__1_n_0;
  wire n25__0_carry_i_14__1_n_0;
  wire n25__0_carry_i_15__1_n_0;
  wire n25__0_carry_i_17__1_n_0;
  wire n25__0_carry_i_18__1_n_0;
  wire n25__0_carry_i_19__1_n_0;
  wire n25__0_carry_i_1__1_n_0;
  wire n25__0_carry_i_20__1_n_0;
  wire n25__0_carry_i_21__0_n_0;
  wire n25__0_carry_i_2__1_n_0;
  wire n25__0_carry_i_3__1_n_0;
  wire n25__0_carry_i_4__1_n_0;
  wire n25__0_carry_i_5__1_n_0;
  wire n25__0_carry_i_6__1_n_0;
  wire n25__0_carry_i_7__1_n_0;
  wire n25__0_carry_i_8__1_n_0;
  wire n25__0_carry_i_9__1_n_0;
  wire n25__0_carry_n_0;
  wire n25__0_carry_n_1;
  wire n25__0_carry_n_10;
  wire n25__0_carry_n_11;
  wire n25__0_carry_n_12;
  wire n25__0_carry_n_2;
  wire n25__0_carry_n_3;
  wire n25__0_carry_n_4;
  wire n25__0_carry_n_5;
  wire n25__0_carry_n_6;
  wire n25__0_carry_n_7;
  wire n25__0_carry_n_8;
  wire n25__0_carry_n_9;
  wire n25__27_carry__0_i_1__1_n_0;
  wire n25__27_carry__0_i_2__1_n_0;
  wire n25__27_carry__0_i_3__1_n_0;
  wire n25__27_carry__0_i_4__1_n_0;
  wire n25__27_carry__0_n_14;
  wire n25__27_carry__0_n_15;
  wire n25__27_carry__0_n_5;
  wire n25__27_carry__0_n_7;
  wire n25__27_carry_i_10__1_n_0;
  wire n25__27_carry_i_11__1_n_0;
  wire n25__27_carry_i_12__1_n_0;
  wire n25__27_carry_i_13__1_n_0;
  wire n25__27_carry_i_14__1_n_0;
  wire n25__27_carry_i_15__1_n_0;
  wire n25__27_carry_i_16__1_n_0;
  wire n25__27_carry_i_17__1_n_0;
  wire n25__27_carry_i_18__1_n_0;
  wire n25__27_carry_i_19__1_n_0;
  wire n25__27_carry_i_1__1_n_0;
  wire n25__27_carry_i_20__1_n_0;
  wire n25__27_carry_i_2__1_n_0;
  wire n25__27_carry_i_3__1_n_0;
  wire n25__27_carry_i_4__1_n_0;
  wire n25__27_carry_i_5__1_n_0;
  wire n25__27_carry_i_6__1_n_0;
  wire n25__27_carry_i_7__1_n_0;
  wire n25__27_carry_i_8__1_n_0;
  wire n25__27_carry_i_9__1_n_0;
  wire n25__27_carry_n_0;
  wire n25__27_carry_n_1;
  wire n25__27_carry_n_10;
  wire n25__27_carry_n_11;
  wire n25__27_carry_n_12;
  wire n25__27_carry_n_13;
  wire n25__27_carry_n_14;
  wire n25__27_carry_n_15;
  wire n25__27_carry_n_2;
  wire n25__27_carry_n_3;
  wire n25__27_carry_n_4;
  wire n25__27_carry_n_5;
  wire n25__27_carry_n_6;
  wire n25__27_carry_n_7;
  wire n25__27_carry_n_8;
  wire n25__27_carry_n_9;
  wire n25__56_carry__0_i_1__1_n_0;
  wire n25__56_carry__0_n_15;
  wire n25__56_carry_i_10__1_n_0;
  wire n25__56_carry_i_11__1_n_0;
  wire n25__56_carry_i_12__1_n_0;
  wire n25__56_carry_i_13__1_n_0;
  wire n25__56_carry_i_14__1_n_0;
  wire n25__56_carry_i_15__1_n_0;
  wire n25__56_carry_i_1__1_n_0;
  wire n25__56_carry_i_2__1_n_0;
  wire n25__56_carry_i_3__1_n_0;
  wire n25__56_carry_i_4__1_n_0;
  wire n25__56_carry_i_5__1_n_0;
  wire n25__56_carry_i_6__1_n_0;
  wire n25__56_carry_i_7__1_n_0;
  wire n25__56_carry_i_8__1_n_0;
  wire n25__56_carry_i_9__1_n_0;
  wire n25__56_carry_n_0;
  wire n25__56_carry_n_1;
  wire n25__56_carry_n_10;
  wire n25__56_carry_n_11;
  wire n25__56_carry_n_12;
  wire n25__56_carry_n_13;
  wire n25__56_carry_n_14;
  wire n25__56_carry_n_15;
  wire n25__56_carry_n_2;
  wire n25__56_carry_n_3;
  wire n25__56_carry_n_4;
  wire n25__56_carry_n_5;
  wire n25__56_carry_n_6;
  wire n25__56_carry_n_7;
  wire n25__56_carry_n_8;
  wire n25__56_carry_n_9;
  wire n25__81_carry__0_i_1__1_n_0;
  wire n25__81_carry__0_i_2__1_n_0;
  wire n25__81_carry__0_i_3__1_n_0;
  wire n25__81_carry__0_i_4__1_n_0;
  wire n25__81_carry__0_i_5__1_n_0;
  wire n25__81_carry__0_i_6__1_n_0;
  wire n25__81_carry__0_i_7__1_n_0;
  wire n25__81_carry__0_n_5;
  wire n25__81_carry__0_n_6;
  wire n25__81_carry__0_n_7;
  wire n25__81_carry_i_10__1_n_0;
  wire n25__81_carry_i_11__1_n_0;
  wire n25__81_carry_i_12__1_n_0;
  wire n25__81_carry_i_13__1_n_0;
  wire n25__81_carry_i_14__1_n_0;
  wire n25__81_carry_i_15__1_n_0;
  wire n25__81_carry_i_1__1_n_0;
  wire n25__81_carry_i_2__1_n_0;
  wire n25__81_carry_i_3__1_n_0;
  wire n25__81_carry_i_4__1_n_0;
  wire n25__81_carry_i_5__1_n_0;
  wire n25__81_carry_i_6__1_n_0;
  wire n25__81_carry_i_7__1_n_0;
  wire n25__81_carry_i_8__1_n_0;
  wire n25__81_carry_i_9__1_n_0;
  wire n25__81_carry_n_0;
  wire n25__81_carry_n_1;
  wire n25__81_carry_n_2;
  wire n25__81_carry_n_3;
  wire n25__81_carry_n_4;
  wire n25__81_carry_n_5;
  wire n25__81_carry_n_6;
  wire n25__81_carry_n_7;
  wire [7:0]n26;
  wire [7:0]n27;
  wire [7:0]n28;
  wire [7:0]n29;
  wire \n29[7]_i_2_n_0 ;
  wire \n29[7]_i_3_n_0 ;
  wire \n29[7]_i_4_n_0 ;
  wire \n29[7]_i_5_n_0 ;
  wire \n29[7]_i_6_n_0 ;
  wire \n29[7]_i_7_n_0 ;
  wire \n29[7]_i_8_n_0 ;
  wire \n29[7]_i_9_n_0 ;
  wire \n29_reg[7]_i_1_n_1 ;
  wire \n29_reg[7]_i_1_n_2 ;
  wire \n29_reg[7]_i_1_n_3 ;
  wire \n29_reg[7]_i_1_n_4 ;
  wire \n29_reg[7]_i_1_n_5 ;
  wire \n29_reg[7]_i_1_n_6 ;
  wire \n29_reg[7]_i_1_n_7 ;
  wire [7:0]n30;
  wire [7:0]n31;
  wire \n33[10]_i_1__1_n_0 ;
  wire \n33[11]_i_1__1_n_0 ;
  wire \n33[12]_i_1__1_n_0 ;
  wire \n33[12]_i_2__1_n_0 ;
  wire \n33[13]_i_1__1_n_0 ;
  wire \n33[14]_i_1__1_n_0 ;
  wire \n33[14]_i_2__1_n_0 ;
  wire \n33[15]_i_2__1_n_0 ;
  wire \n33[2]_i_1__1_n_0 ;
  wire \n33[3]_i_1__1_n_0 ;
  wire \n33[4]_i_1__1_n_0 ;
  wire \n33[4]_i_2__1_n_0 ;
  wire \n33[5]_i_1__1_n_0 ;
  wire \n33[6]_i_1__1_n_0 ;
  wire \n33[6]_i_2__1_n_0 ;
  wire \n33[7]_i_2__1_n_0 ;
  wire \n33[9]_i_1__1_n_0 ;
  wire [7:1]n341_out;
  wire [7:1]n350_out;
  wire \n37[12]_i_2__1_n_0 ;
  wire \n37[14]_i_2__1_n_0 ;
  wire \n37[15]_i_2__1_n_0 ;
  wire \n37[4]_i_2__1_n_0 ;
  wire \n37[6]_i_2__1_n_0 ;
  wire \n37[7]_i_2__1_n_0 ;
  wire [7:0]n4;
  wire \n7_reg_n_0_[0] ;
  wire \n7_reg_n_0_[1] ;
  wire \n7_reg_n_0_[2] ;
  wire \n7_reg_n_0_[3] ;
  wire \n7_reg_n_0_[4] ;
  wire \n7_reg_n_0_[5] ;
  wire \n7_reg_n_0_[6] ;
  wire \n7_reg_n_0_[7] ;
  wire \n8_reg_n_0_[0] ;
  wire \n8_reg_n_0_[1] ;
  wire \n8_reg_n_0_[2] ;
  wire \n8_reg_n_0_[3] ;
  wire \n8_reg_n_0_[4] ;
  wire \n8_reg_n_0_[5] ;
  wire \n8_reg_n_0_[6] ;
  wire \n8_reg_n_0_[7] ;
  wire \n9_reg_n_0_[0] ;
  wire \n9_reg_n_0_[1] ;
  wire \n9_reg_n_0_[2] ;
  wire \n9_reg_n_0_[3] ;
  wire \n9_reg_n_0_[4] ;
  wire \n9_reg_n_0_[5] ;
  wire \n9_reg_n_0_[6] ;
  wire \n9_reg_n_0_[7] ;
  wire rst_i;
  wire [15:0]s4_3;
  wire [2:0]NLW_n14__0_carry_O_UNCONNECTED;
  wire [7:1]NLW_n14__0_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n14__0_carry__0_O_UNCONNECTED;
  wire [7:1]NLW_n14__27_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n14__27_carry__0_O_UNCONNECTED;
  wire [7:0]NLW_n14__56_carry__0_CO_UNCONNECTED;
  wire [7:1]NLW_n14__56_carry__0_O_UNCONNECTED;
  wire [3:0]NLW_n14__81_carry_O_UNCONNECTED;
  wire [7:3]NLW_n14__81_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n14__81_carry__0_O_UNCONNECTED;
  wire [2:0]NLW_n17__0_carry_O_UNCONNECTED;
  wire [7:1]NLW_n17__0_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n17__0_carry__0_O_UNCONNECTED;
  wire [7:1]NLW_n17__27_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n17__27_carry__0_O_UNCONNECTED;
  wire [7:0]NLW_n17__56_carry__0_CO_UNCONNECTED;
  wire [7:1]NLW_n17__56_carry__0_O_UNCONNECTED;
  wire [3:0]NLW_n17__81_carry_O_UNCONNECTED;
  wire [7:3]NLW_n17__81_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n17__81_carry__0_O_UNCONNECTED;
  wire [7:7]NLW_n20_carry_CO_UNCONNECTED;
  wire [2:0]NLW_n22__0_carry_O_UNCONNECTED;
  wire [7:1]NLW_n22__0_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n22__0_carry__0_O_UNCONNECTED;
  wire [7:1]NLW_n22__27_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n22__27_carry__0_O_UNCONNECTED;
  wire [7:0]NLW_n22__56_carry__0_CO_UNCONNECTED;
  wire [7:1]NLW_n22__56_carry__0_O_UNCONNECTED;
  wire [3:0]NLW_n22__81_carry_O_UNCONNECTED;
  wire [7:3]NLW_n22__81_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n22__81_carry__0_O_UNCONNECTED;
  wire [2:0]NLW_n25__0_carry_O_UNCONNECTED;
  wire [7:1]NLW_n25__0_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n25__0_carry__0_O_UNCONNECTED;
  wire [7:1]NLW_n25__27_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n25__27_carry__0_O_UNCONNECTED;
  wire [7:0]NLW_n25__56_carry__0_CO_UNCONNECTED;
  wire [7:1]NLW_n25__56_carry__0_O_UNCONNECTED;
  wire [3:0]NLW_n25__81_carry_O_UNCONNECTED;
  wire [7:3]NLW_n25__81_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n25__81_carry__0_O_UNCONNECTED;
  wire [7:7]\NLW_n29_reg[7]_i_1_CO_UNCONNECTED ;

  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[0] ),
        .Q(n10[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[1] ),
        .Q(n10[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[2] ),
        .Q(n10[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[3] ),
        .Q(n10[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[4] ),
        .Q(n10[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[5] ),
        .Q(n10[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[6] ),
        .Q(n10[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[7] ),
        .Q(n10[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__0_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__0_carry_n_0,n14__0_carry_n_1,n14__0_carry_n_2,n14__0_carry_n_3,n14__0_carry_n_4,n14__0_carry_n_5,n14__0_carry_n_6,n14__0_carry_n_7}),
        .DI({n14__0_carry_i_1__1_n_0,n14__0_carry_i_2__1_n_0,n14__0_carry_i_3__1_n_0,n14__0_carry_i_4__1_n_0,n14__0_carry_i_5__1_n_0,n14__0_carry_i_6__1_n_0,n14__0_carry_i_7__1_n_0,1'b0}),
        .O({n14__0_carry_n_8,n14__0_carry_n_9,n14__0_carry_n_10,n14__0_carry_n_11,n14__0_carry_n_12,NLW_n14__0_carry_O_UNCONNECTED[2:0]}),
        .S({n14__0_carry_i_8__1_n_0,n14__0_carry_i_9__1_n_0,n14__0_carry_i_10__1_n_0,n14__0_carry_i_11__1_n_0,n14__0_carry_i_12__1_n_0,n14__0_carry_i_13__1_n_0,n14__0_carry_i_14__1_n_0,n14__0_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__0_carry__0
       (.CI(n14__0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__0_carry__0_CO_UNCONNECTED[7:3],n14__0_carry__0_n_5,NLW_n14__0_carry__0_CO_UNCONNECTED[1],n14__0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14__0_carry__0_i_1__1_n_0,n14__0_carry__0_i_2__1_n_0}),
        .O({NLW_n14__0_carry__0_O_UNCONNECTED[7:2],n14__0_carry__0_n_14,n14__0_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n14__0_carry__0_i_3__1_n_0,n14__0_carry__0_i_4__1_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__0_carry__0_i_1__1
       (.I0(n14__56_carry_0[9]),
        .I1(n22_n_0),
        .I2(n14__56_carry_0[10]),
        .I3(n22__0_n_0),
        .O(n14__0_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n14__0_carry__0_i_2__1
       (.I0(n14__56_carry_0[10]),
        .I1(n22__1_n_0),
        .I2(n14__56_carry_0[9]),
        .I3(n22__0_n_0),
        .I4(n14__56_carry_0[8]),
        .I5(n22_n_0),
        .O(n14__0_carry__0_i_2__1_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n14__0_carry__0_i_3__1
       (.I0(n22__0_n_0),
        .I1(n14__56_carry_0[9]),
        .I2(n14__56_carry_0[10]),
        .I3(n22_n_0),
        .O(n14__0_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n14__0_carry__0_i_4__1
       (.I0(n14__56_carry_0[8]),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(n14__56_carry_0[10]),
        .I4(n22_n_0),
        .I5(n14__56_carry_0[9]),
        .O(n14__0_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__0_carry_i_10__1
       (.I0(n14__0_carry_i_3__1_n_0),
        .I1(n14__56_carry_0[9]),
        .I2(n22__2_n_0),
        .I3(n14__0_carry_i_18__1_n_0),
        .I4(n22__1_n_0),
        .I5(n14__56_carry_0[8]),
        .O(n14__0_carry_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__0_carry_i_11__1
       (.I0(n14__0_carry_i_4__1_n_0),
        .I1(n14__56_carry_0[9]),
        .I2(n22__3_n_0),
        .I3(n14__0_carry_i_19__1_n_0),
        .I4(n22__2_n_0),
        .I5(n14__56_carry_0[8]),
        .O(n14__0_carry_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n14__0_carry_i_12__1
       (.I0(n22__4_n_0),
        .I1(n14__0_carry_i_20__1_n_0),
        .I2(n22__5_n_0),
        .I3(n14__56_carry_0[9]),
        .I4(n22__6_n_0),
        .I5(n14__56_carry_0[10]),
        .O(n14__0_carry_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n14__0_carry_i_13__1
       (.I0(n22__6_n_0),
        .I1(n14__56_carry_0[10]),
        .I2(n22__5_n_0),
        .I3(n14__56_carry_0[9]),
        .I4(n14__56_carry_0[8]),
        .I5(n22__4_n_0),
        .O(n14__0_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__0_carry_i_14__1
       (.I0(n14__56_carry_0[8]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[9]),
        .I3(n22__6_n_0),
        .O(n14__0_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__0_carry_i_15__1
       (.I0(n22__6_n_0),
        .I1(n14__56_carry_0[8]),
        .O(n14__0_carry_i_15__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_16__1
       (.I0(n22__1_n_0),
        .I1(n14__56_carry_0[10]),
        .O(n14__0_carry_i_16__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_17__1
       (.I0(n22__2_n_0),
        .I1(n14__56_carry_0[10]),
        .O(n14__0_carry_i_17__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_18__1
       (.I0(n22__3_n_0),
        .I1(n14__56_carry_0[10]),
        .O(n14__0_carry_i_18__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_19__1
       (.I0(n22__4_n_0),
        .I1(n14__56_carry_0[10]),
        .O(n14__0_carry_i_19__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__0_carry_i_1__1
       (.I0(n14__56_carry_0[10]),
        .I1(n22__2_n_0),
        .I2(n14__56_carry_0[9]),
        .I3(n22__1_n_0),
        .I4(n14__56_carry_0[8]),
        .I5(n22__0_n_0),
        .O(n14__0_carry_i_1__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_20__1
       (.I0(n22__3_n_0),
        .I1(n14__56_carry_0[8]),
        .O(n14__0_carry_i_20__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__0_carry_i_2__1
       (.I0(n14__56_carry_0[10]),
        .I1(n22__3_n_0),
        .I2(n14__56_carry_0[9]),
        .I3(n22__2_n_0),
        .I4(n14__56_carry_0[8]),
        .I5(n22__1_n_0),
        .O(n14__0_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__0_carry_i_3__1
       (.I0(n14__56_carry_0[10]),
        .I1(n22__4_n_0),
        .I2(n14__56_carry_0[9]),
        .I3(n22__3_n_0),
        .I4(n14__56_carry_0[8]),
        .I5(n22__2_n_0),
        .O(n14__0_carry_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__0_carry_i_4__1
       (.I0(n14__56_carry_0[10]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[9]),
        .I3(n22__4_n_0),
        .I4(n14__56_carry_0[8]),
        .I5(n22__3_n_0),
        .O(n14__0_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n14__0_carry_i_5__1
       (.I0(n14__56_carry_0[9]),
        .I1(n22__4_n_0),
        .I2(n14__56_carry_0[10]),
        .I3(n22__5_n_0),
        .I4(n22__3_n_0),
        .I5(n14__56_carry_0[8]),
        .O(n14__0_carry_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__0_carry_i_6__1
       (.I0(n14__56_carry_0[9]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[10]),
        .I3(n22__6_n_0),
        .O(n14__0_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__0_carry_i_7__1
       (.I0(n14__56_carry_0[8]),
        .I1(n22__5_n_0),
        .O(n14__0_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n14__0_carry_i_8__1
       (.I0(n14__0_carry_i_1__1_n_0),
        .I1(n14__56_carry_0[9]),
        .I2(n22__0_n_0),
        .I3(n14__0_carry_i_16__1_n_0),
        .I4(n22_n_0),
        .I5(n14__56_carry_0[8]),
        .O(n14__0_carry_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__0_carry_i_9__1
       (.I0(n14__0_carry_i_2__1_n_0),
        .I1(n14__56_carry_0[9]),
        .I2(n22__1_n_0),
        .I3(n14__0_carry_i_17__1_n_0),
        .I4(n22__0_n_0),
        .I5(n14__56_carry_0[8]),
        .O(n14__0_carry_i_9__1_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__27_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__27_carry_n_0,n14__27_carry_n_1,n14__27_carry_n_2,n14__27_carry_n_3,n14__27_carry_n_4,n14__27_carry_n_5,n14__27_carry_n_6,n14__27_carry_n_7}),
        .DI({n14__27_carry_i_1__1_n_0,n14__27_carry_i_2__1_n_0,n14__27_carry_i_3__1_n_0,n14__27_carry_i_4__1_n_0,n14__27_carry_i_5__1_n_0,n14__27_carry_i_6__1_n_0,n14__27_carry_i_7__1_n_0,1'b0}),
        .O({n14__27_carry_n_8,n14__27_carry_n_9,n14__27_carry_n_10,n14__27_carry_n_11,n14__27_carry_n_12,n14__27_carry_n_13,n14__27_carry_n_14,n14__27_carry_n_15}),
        .S({n14__27_carry_i_8__1_n_0,n14__27_carry_i_9__1_n_0,n14__27_carry_i_10__1_n_0,n14__27_carry_i_11__1_n_0,n14__27_carry_i_12__1_n_0,n14__27_carry_i_13__1_n_0,n14__27_carry_i_14__1_n_0,n14__27_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__27_carry__0
       (.CI(n14__27_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__27_carry__0_CO_UNCONNECTED[7:3],n14__27_carry__0_n_5,NLW_n14__27_carry__0_CO_UNCONNECTED[1],n14__27_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14__27_carry__0_i_1__1_n_0,n14__27_carry__0_i_2__1_n_0}),
        .O({NLW_n14__27_carry__0_O_UNCONNECTED[7:2],n14__27_carry__0_n_14,n14__27_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n14__27_carry__0_i_3__1_n_0,n14__27_carry__0_i_4__1_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__27_carry__0_i_1__1
       (.I0(n14__56_carry_0[12]),
        .I1(n22_n_0),
        .I2(n14__56_carry_0[13]),
        .I3(n22__0_n_0),
        .O(n14__27_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n14__27_carry__0_i_2__1
       (.I0(n14__56_carry_0[13]),
        .I1(n22__1_n_0),
        .I2(n14__56_carry_0[12]),
        .I3(n22__0_n_0),
        .I4(n14__56_carry_0[11]),
        .I5(n22_n_0),
        .O(n14__27_carry__0_i_2__1_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n14__27_carry__0_i_3__1
       (.I0(n22__0_n_0),
        .I1(n14__56_carry_0[12]),
        .I2(n14__56_carry_0[13]),
        .I3(n22_n_0),
        .O(n14__27_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n14__27_carry__0_i_4__1
       (.I0(n14__56_carry_0[11]),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(n14__56_carry_0[13]),
        .I4(n22_n_0),
        .I5(n14__56_carry_0[12]),
        .O(n14__27_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__27_carry_i_10__1
       (.I0(n14__27_carry_i_3__1_n_0),
        .I1(n14__56_carry_0[12]),
        .I2(n22__2_n_0),
        .I3(n14__27_carry_i_18__1_n_0),
        .I4(n22__1_n_0),
        .I5(n14__56_carry_0[11]),
        .O(n14__27_carry_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__27_carry_i_11__1
       (.I0(n14__27_carry_i_4__1_n_0),
        .I1(n14__56_carry_0[12]),
        .I2(n22__3_n_0),
        .I3(n14__27_carry_i_19__1_n_0),
        .I4(n22__2_n_0),
        .I5(n14__56_carry_0[11]),
        .O(n14__27_carry_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n14__27_carry_i_12__1
       (.I0(n22__4_n_0),
        .I1(n14__27_carry_i_20__1_n_0),
        .I2(n22__5_n_0),
        .I3(n14__56_carry_0[12]),
        .I4(n22__6_n_0),
        .I5(n14__56_carry_0[13]),
        .O(n14__27_carry_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n14__27_carry_i_13__1
       (.I0(n22__6_n_0),
        .I1(n14__56_carry_0[13]),
        .I2(n22__5_n_0),
        .I3(n14__56_carry_0[12]),
        .I4(n14__56_carry_0[11]),
        .I5(n22__4_n_0),
        .O(n14__27_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__27_carry_i_14__1
       (.I0(n14__56_carry_0[11]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[12]),
        .I3(n22__6_n_0),
        .O(n14__27_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__27_carry_i_15__1
       (.I0(n22__6_n_0),
        .I1(n14__56_carry_0[11]),
        .O(n14__27_carry_i_15__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_16__1
       (.I0(n22__1_n_0),
        .I1(n14__56_carry_0[13]),
        .O(n14__27_carry_i_16__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_17__1
       (.I0(n22__2_n_0),
        .I1(n14__56_carry_0[13]),
        .O(n14__27_carry_i_17__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_18__1
       (.I0(n22__3_n_0),
        .I1(n14__56_carry_0[13]),
        .O(n14__27_carry_i_18__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_19__1
       (.I0(n22__4_n_0),
        .I1(n14__56_carry_0[13]),
        .O(n14__27_carry_i_19__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__27_carry_i_1__1
       (.I0(n14__56_carry_0[13]),
        .I1(n22__2_n_0),
        .I2(n14__56_carry_0[12]),
        .I3(n22__1_n_0),
        .I4(n14__56_carry_0[11]),
        .I5(n22__0_n_0),
        .O(n14__27_carry_i_1__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_20__1
       (.I0(n22__3_n_0),
        .I1(n14__56_carry_0[11]),
        .O(n14__27_carry_i_20__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__27_carry_i_2__1
       (.I0(n14__56_carry_0[13]),
        .I1(n22__3_n_0),
        .I2(n14__56_carry_0[12]),
        .I3(n22__2_n_0),
        .I4(n14__56_carry_0[11]),
        .I5(n22__1_n_0),
        .O(n14__27_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__27_carry_i_3__1
       (.I0(n14__56_carry_0[13]),
        .I1(n22__4_n_0),
        .I2(n14__56_carry_0[12]),
        .I3(n22__3_n_0),
        .I4(n14__56_carry_0[11]),
        .I5(n22__2_n_0),
        .O(n14__27_carry_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__27_carry_i_4__1
       (.I0(n14__56_carry_0[13]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[12]),
        .I3(n22__4_n_0),
        .I4(n14__56_carry_0[11]),
        .I5(n22__3_n_0),
        .O(n14__27_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n14__27_carry_i_5__1
       (.I0(n14__56_carry_0[12]),
        .I1(n22__4_n_0),
        .I2(n14__56_carry_0[13]),
        .I3(n22__5_n_0),
        .I4(n22__3_n_0),
        .I5(n14__56_carry_0[11]),
        .O(n14__27_carry_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__27_carry_i_6__1
       (.I0(n14__56_carry_0[12]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[13]),
        .I3(n22__6_n_0),
        .O(n14__27_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__27_carry_i_7__1
       (.I0(n14__56_carry_0[11]),
        .I1(n22__5_n_0),
        .O(n14__27_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n14__27_carry_i_8__1
       (.I0(n14__27_carry_i_1__1_n_0),
        .I1(n14__56_carry_0[12]),
        .I2(n22__0_n_0),
        .I3(n14__27_carry_i_16__1_n_0),
        .I4(n22_n_0),
        .I5(n14__56_carry_0[11]),
        .O(n14__27_carry_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__27_carry_i_9__1
       (.I0(n14__27_carry_i_2__1_n_0),
        .I1(n14__56_carry_0[12]),
        .I2(n22__1_n_0),
        .I3(n14__27_carry_i_17__1_n_0),
        .I4(n22__0_n_0),
        .I5(n14__56_carry_0[11]),
        .O(n14__27_carry_i_9__1_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__56_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__56_carry_n_0,n14__56_carry_n_1,n14__56_carry_n_2,n14__56_carry_n_3,n14__56_carry_n_4,n14__56_carry_n_5,n14__56_carry_n_6,n14__56_carry_n_7}),
        .DI({n14__56_carry_i_1__1_n_0,n14__56_carry_i_2__1_n_0,n14__56_carry_i_3__1_n_0,n14__56_carry_i_4__1_n_0,n14__56_carry_i_5__1_n_0,n14__56_carry_i_6__1_n_0,n14__56_carry_i_7__1_n_0,1'b0}),
        .O({n14__56_carry_n_8,n14__56_carry_n_9,n14__56_carry_n_10,n14__56_carry_n_11,n14__56_carry_n_12,n14__56_carry_n_13,n14__56_carry_n_14,n14__56_carry_n_15}),
        .S({n14__56_carry_i_8__1_n_0,n14__56_carry_i_9__1_n_0,n14__56_carry_i_10__1_n_0,n14__56_carry_i_11__1_n_0,n14__56_carry_i_12__1_n_0,n14__56_carry_i_13__1_n_0,n14__56_carry_i_14__1_n_0,n14__56_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__56_carry__0
       (.CI(n14__56_carry_n_0),
        .CI_TOP(1'b0),
        .CO(NLW_n14__56_carry__0_CO_UNCONNECTED[7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_n14__56_carry__0_O_UNCONNECTED[7:1],n14__56_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14__56_carry__0_i_1__1_n_0}));
  LUT4 #(
    .INIT(16'hE53F)) 
    n14__56_carry__0_i_1__1
       (.I0(n14__56_carry_0[14]),
        .I1(n22__0_n_0),
        .I2(n14__56_carry_0[15]),
        .I3(n22_n_0),
        .O(n14__56_carry__0_i_1__1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n14__56_carry_i_10__1
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(n14__56_carry_0[15]),
        .I3(n22__1_n_0),
        .I4(n14__56_carry_0[14]),
        .O(n14__56_carry_i_10__1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n14__56_carry_i_11__1
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n14__56_carry_0[15]),
        .I3(n22__2_n_0),
        .I4(n14__56_carry_0[14]),
        .O(n14__56_carry_i_11__1_n_0));
  LUT5 #(
    .INIT(32'h9F606060)) 
    n14__56_carry_i_12__1
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(n14__56_carry_0[15]),
        .I3(n22__3_n_0),
        .I4(n14__56_carry_0[14]),
        .O(n14__56_carry_i_12__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__56_carry_i_13__1
       (.I0(n14__56_carry_0[15]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[14]),
        .I3(n22__4_n_0),
        .O(n14__56_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h8777)) 
    n14__56_carry_i_14__1
       (.I0(n14__56_carry_0[15]),
        .I1(n22__6_n_0),
        .I2(n14__56_carry_0[14]),
        .I3(n22__5_n_0),
        .O(n14__56_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__56_carry_i_15__1
       (.I0(n22__6_n_0),
        .I1(n14__56_carry_0[14]),
        .O(n14__56_carry_i_15__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__56_carry_i_1__1
       (.I0(n14__56_carry_0[15]),
        .I1(n22__1_n_0),
        .I2(n14__56_carry_0[14]),
        .I3(n22__0_n_0),
        .O(n14__56_carry_i_1__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__56_carry_i_2__1
       (.I0(n14__56_carry_0[15]),
        .I1(n22__2_n_0),
        .I2(n14__56_carry_0[14]),
        .I3(n22__1_n_0),
        .O(n14__56_carry_i_2__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__56_carry_i_3__1
       (.I0(n14__56_carry_0[15]),
        .I1(n22__3_n_0),
        .I2(n14__56_carry_0[14]),
        .I3(n22__2_n_0),
        .O(n14__56_carry_i_3__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__56_carry_i_4__1
       (.I0(n14__56_carry_0[15]),
        .I1(n22__4_n_0),
        .I2(n14__56_carry_0[14]),
        .I3(n22__3_n_0),
        .O(n14__56_carry_i_4__1_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n14__56_carry_i_5__1
       (.I0(n22__5_n_0),
        .I1(n14__56_carry_0[15]),
        .O(n14__56_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__56_carry_i_6__1
       (.I0(n14__56_carry_0[15]),
        .I1(n22__5_n_0),
        .O(n14__56_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n14__56_carry_i_7__1
       (.I0(n22__6_n_0),
        .I1(n14__56_carry_0[15]),
        .O(n14__56_carry_i_7__1_n_0));
  LUT5 #(
    .INIT(32'h738CC0C0)) 
    n14__56_carry_i_8__1
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n14__56_carry_0[15]),
        .I3(n22_n_0),
        .I4(n14__56_carry_0[14]),
        .O(n14__56_carry_i_8__1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n14__56_carry_i_9__1
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(n14__56_carry_0[15]),
        .I3(n22__0_n_0),
        .I4(n14__56_carry_0[14]),
        .O(n14__56_carry_i_9__1_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__81_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__81_carry_n_0,n14__81_carry_n_1,n14__81_carry_n_2,n14__81_carry_n_3,n14__81_carry_n_4,n14__81_carry_n_5,n14__81_carry_n_6,n14__81_carry_n_7}),
        .DI({n14__81_carry_i_1__1_n_0,n14__81_carry_i_2__1_n_0,n14__81_carry_i_3__1_n_0,n14__81_carry_i_4__1_n_0,n14__81_carry_i_5__1_n_0,n14__81_carry_i_6__1_n_0,n14__81_carry_i_7__1_n_0,1'b0}),
        .O({n15[3:0],NLW_n14__81_carry_O_UNCONNECTED[3:0]}),
        .S({n14__81_carry_i_8__1_n_0,n14__81_carry_i_9__1_n_0,n14__81_carry_i_10__1_n_0,n14__81_carry_i_11__1_n_0,n14__81_carry_i_12__1_n_0,n14__81_carry_i_13__1_n_0,n14__81_carry_i_14__1_n_0,n14__81_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__81_carry__0
       (.CI(n14__81_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__81_carry__0_CO_UNCONNECTED[7:3],n14__81_carry__0_n_5,n14__81_carry__0_n_6,n14__81_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n14__81_carry__0_i_1__1_n_0,n14__81_carry__0_i_2__1_n_0,n14__81_carry__0_i_3__1_n_0}),
        .O({NLW_n14__81_carry__0_O_UNCONNECTED[7:4],n15[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n14__81_carry__0_i_4__1_n_0,n14__81_carry__0_i_5__1_n_0,n14__81_carry__0_i_6__1_n_0,n14__81_carry__0_i_7__1_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry__0_i_1__1
       (.I0(n14__27_carry__0_n_14),
        .I1(n14__56_carry_n_9),
        .O(n14__81_carry__0_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry__0_i_2__1
       (.I0(n14__27_carry__0_n_15),
        .I1(n14__56_carry_n_10),
        .O(n14__81_carry__0_i_2__1_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry__0_i_3__1
       (.I0(n14__56_carry_n_11),
        .I1(n14__27_carry_n_8),
        .I2(n14__0_carry__0_n_5),
        .O(n14__81_carry__0_i_3__1_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n14__81_carry__0_i_4__1
       (.I0(n14__27_carry__0_n_5),
        .I1(n14__56_carry_n_8),
        .I2(n14__56_carry__0_n_15),
        .O(n14__81_carry__0_i_4__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__81_carry__0_i_5__1
       (.I0(n14__27_carry__0_n_14),
        .I1(n14__56_carry_n_9),
        .I2(n14__56_carry_n_8),
        .I3(n14__27_carry__0_n_5),
        .O(n14__81_carry__0_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__81_carry__0_i_6__1
       (.I0(n14__27_carry__0_n_15),
        .I1(n14__56_carry_n_10),
        .I2(n14__56_carry_n_9),
        .I3(n14__27_carry__0_n_14),
        .O(n14__81_carry__0_i_6__1_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n14__81_carry__0_i_7__1
       (.I0(n14__0_carry__0_n_5),
        .I1(n14__27_carry_n_8),
        .I2(n14__56_carry_n_11),
        .I3(n14__56_carry_n_10),
        .I4(n14__27_carry__0_n_15),
        .O(n14__81_carry__0_i_7__1_n_0));
  (* HLUTNM = "lutpair30" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_10__1
       (.I0(n14__56_carry_n_13),
        .I1(n14__27_carry_n_10),
        .I2(n14__0_carry__0_n_15),
        .I3(n14__81_carry_i_3__1_n_0),
        .O(n14__81_carry_i_10__1_n_0));
  (* HLUTNM = "lutpair29" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_11__1
       (.I0(n14__56_carry_n_14),
        .I1(n14__27_carry_n_11),
        .I2(n14__0_carry_n_8),
        .I3(n14__81_carry_i_4__1_n_0),
        .O(n14__81_carry_i_11__1_n_0));
  (* HLUTNM = "lutpair28" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_12__1
       (.I0(n14__56_carry_n_15),
        .I1(n14__27_carry_n_12),
        .I2(n14__0_carry_n_9),
        .I3(n14__81_carry_i_5__1_n_0),
        .O(n14__81_carry_i_12__1_n_0));
  (* HLUTNM = "lutpair87" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n14__81_carry_i_13__1
       (.I0(n14__27_carry_n_13),
        .I1(n14__0_carry_n_10),
        .I2(n14__0_carry_n_11),
        .I3(n14__27_carry_n_14),
        .O(n14__81_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__81_carry_i_14__1
       (.I0(n14__0_carry_n_12),
        .I1(n14__27_carry_n_15),
        .I2(n14__27_carry_n_14),
        .I3(n14__0_carry_n_11),
        .O(n14__81_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n14__81_carry_i_15__1
       (.I0(n14__0_carry_n_12),
        .I1(n14__27_carry_n_15),
        .O(n14__81_carry_i_15__1_n_0));
  (* HLUTNM = "lutpair31" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry_i_1__1
       (.I0(n14__56_carry_n_12),
        .I1(n14__27_carry_n_9),
        .I2(n14__0_carry__0_n_14),
        .O(n14__81_carry_i_1__1_n_0));
  (* HLUTNM = "lutpair30" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry_i_2__1
       (.I0(n14__56_carry_n_13),
        .I1(n14__27_carry_n_10),
        .I2(n14__0_carry__0_n_15),
        .O(n14__81_carry_i_2__1_n_0));
  (* HLUTNM = "lutpair29" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry_i_3__1
       (.I0(n14__56_carry_n_14),
        .I1(n14__27_carry_n_11),
        .I2(n14__0_carry_n_8),
        .O(n14__81_carry_i_3__1_n_0));
  (* HLUTNM = "lutpair28" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry_i_4__1
       (.I0(n14__56_carry_n_15),
        .I1(n14__27_carry_n_12),
        .I2(n14__0_carry_n_9),
        .O(n14__81_carry_i_4__1_n_0));
  (* HLUTNM = "lutpair87" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry_i_5__1
       (.I0(n14__27_carry_n_13),
        .I1(n14__0_carry_n_10),
        .O(n14__81_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry_i_6__1
       (.I0(n14__0_carry_n_11),
        .I1(n14__27_carry_n_14),
        .O(n14__81_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry_i_7__1
       (.I0(n14__0_carry_n_12),
        .I1(n14__27_carry_n_15),
        .O(n14__81_carry_i_7__1_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_8__1
       (.I0(n14__81_carry_i_1__1_n_0),
        .I1(n14__27_carry_n_8),
        .I2(n14__56_carry_n_11),
        .I3(n14__0_carry__0_n_5),
        .O(n14__81_carry_i_8__1_n_0));
  (* HLUTNM = "lutpair31" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_9__1
       (.I0(n14__56_carry_n_12),
        .I1(n14__27_carry_n_9),
        .I2(n14__0_carry__0_n_14),
        .I3(n14__81_carry_i_2__1_n_0),
        .O(n14__81_carry_i_9__1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[0]),
        .Q(\n16_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[1]),
        .Q(\n16_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[2]),
        .Q(\n16_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[3]),
        .Q(\n16_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[4]),
        .Q(\n16_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[5]),
        .Q(\n16_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[6]),
        .Q(\n16_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[7]),
        .Q(\n16_reg_n_0_[7] ),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__0_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n17__0_carry_n_0,n17__0_carry_n_1,n17__0_carry_n_2,n17__0_carry_n_3,n17__0_carry_n_4,n17__0_carry_n_5,n17__0_carry_n_6,n17__0_carry_n_7}),
        .DI({n17__0_carry_i_1__1_n_0,n17__0_carry_i_2__1_n_0,n17__0_carry_i_3__1_n_0,n17__0_carry_i_4__1_n_0,n17__0_carry_i_5__1_n_0,n17__0_carry_i_6__1_n_0,n17__0_carry_i_7__1_n_0,1'b0}),
        .O({n17__0_carry_n_8,n17__0_carry_n_9,n17__0_carry_n_10,n17__0_carry_n_11,n17__0_carry_n_12,NLW_n17__0_carry_O_UNCONNECTED[2:0]}),
        .S({n17__0_carry_i_8__1_n_0,n17__0_carry_i_9__1_n_0,n17__0_carry_i_10__1_n_0,n17__0_carry_i_11__1_n_0,n17__0_carry_i_12__1_n_0,n17__0_carry_i_13__1_n_0,n17__0_carry_i_14__1_n_0,n17__0_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__0_carry__0
       (.CI(n17__0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n17__0_carry__0_CO_UNCONNECTED[7:3],n17__0_carry__0_n_5,NLW_n17__0_carry__0_CO_UNCONNECTED[1],n17__0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n17__0_carry__0_i_1__1_n_0,n17__0_carry__0_i_2__1_n_0}),
        .O({NLW_n17__0_carry__0_O_UNCONNECTED[7:2],n17__0_carry__0_n_14,n17__0_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n17__0_carry__0_i_3__1_n_0,n17__0_carry__0_i_4__1_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__0_carry__0_i_1__1
       (.I0(n14__56_carry_0[1]),
        .I1(n4[7]),
        .I2(n14__56_carry_0[2]),
        .I3(n4[6]),
        .O(n17__0_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n17__0_carry__0_i_2__1
       (.I0(n14__56_carry_0[2]),
        .I1(n4[5]),
        .I2(n14__56_carry_0[1]),
        .I3(n4[6]),
        .I4(n14__56_carry_0[0]),
        .I5(n4[7]),
        .O(n17__0_carry__0_i_2__1_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n17__0_carry__0_i_3__1
       (.I0(n4[6]),
        .I1(n14__56_carry_0[1]),
        .I2(n14__56_carry_0[2]),
        .I3(n4[7]),
        .O(n17__0_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n17__0_carry__0_i_4__1
       (.I0(n14__56_carry_0[0]),
        .I1(n4[5]),
        .I2(n4[6]),
        .I3(n14__56_carry_0[2]),
        .I4(n4[7]),
        .I5(n14__56_carry_0[1]),
        .O(n17__0_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__0_carry_i_10__1
       (.I0(n17__0_carry_i_3__1_n_0),
        .I1(n14__56_carry_0[1]),
        .I2(n4[4]),
        .I3(n17__0_carry_i_18__1_n_0),
        .I4(n4[5]),
        .I5(n14__56_carry_0[0]),
        .O(n17__0_carry_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__0_carry_i_11__1
       (.I0(n17__0_carry_i_4__1_n_0),
        .I1(n14__56_carry_0[1]),
        .I2(n4[3]),
        .I3(n17__0_carry_i_19__1_n_0),
        .I4(n4[4]),
        .I5(n14__56_carry_0[0]),
        .O(n17__0_carry_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n17__0_carry_i_12__1
       (.I0(n4[2]),
        .I1(n17__0_carry_i_20__1_n_0),
        .I2(n4[1]),
        .I3(n14__56_carry_0[1]),
        .I4(n4[0]),
        .I5(n14__56_carry_0[2]),
        .O(n17__0_carry_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n17__0_carry_i_13__1
       (.I0(n4[0]),
        .I1(n14__56_carry_0[2]),
        .I2(n4[1]),
        .I3(n14__56_carry_0[1]),
        .I4(n14__56_carry_0[0]),
        .I5(n4[2]),
        .O(n17__0_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__0_carry_i_14__1
       (.I0(n14__56_carry_0[0]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[1]),
        .I3(n4[0]),
        .O(n17__0_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__0_carry_i_15__1
       (.I0(n4[0]),
        .I1(n14__56_carry_0[0]),
        .O(n17__0_carry_i_15__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_16__1
       (.I0(n4[5]),
        .I1(n14__56_carry_0[2]),
        .O(n17__0_carry_i_16__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_17__1
       (.I0(n4[4]),
        .I1(n14__56_carry_0[2]),
        .O(n17__0_carry_i_17__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_18__1
       (.I0(n4[3]),
        .I1(n14__56_carry_0[2]),
        .O(n17__0_carry_i_18__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_19__1
       (.I0(n4[2]),
        .I1(n14__56_carry_0[2]),
        .O(n17__0_carry_i_19__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__0_carry_i_1__1
       (.I0(n14__56_carry_0[2]),
        .I1(n4[4]),
        .I2(n14__56_carry_0[1]),
        .I3(n4[5]),
        .I4(n14__56_carry_0[0]),
        .I5(n4[6]),
        .O(n17__0_carry_i_1__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_20__1
       (.I0(n4[3]),
        .I1(n14__56_carry_0[0]),
        .O(n17__0_carry_i_20__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__0_carry_i_2__1
       (.I0(n14__56_carry_0[2]),
        .I1(n4[3]),
        .I2(n14__56_carry_0[1]),
        .I3(n4[4]),
        .I4(n14__56_carry_0[0]),
        .I5(n4[5]),
        .O(n17__0_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__0_carry_i_3__1
       (.I0(n14__56_carry_0[2]),
        .I1(n4[2]),
        .I2(n14__56_carry_0[1]),
        .I3(n4[3]),
        .I4(n14__56_carry_0[0]),
        .I5(n4[4]),
        .O(n17__0_carry_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__0_carry_i_4__1
       (.I0(n14__56_carry_0[2]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[1]),
        .I3(n4[2]),
        .I4(n14__56_carry_0[0]),
        .I5(n4[3]),
        .O(n17__0_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n17__0_carry_i_5__1
       (.I0(n14__56_carry_0[1]),
        .I1(n4[2]),
        .I2(n14__56_carry_0[2]),
        .I3(n4[1]),
        .I4(n4[3]),
        .I5(n14__56_carry_0[0]),
        .O(n17__0_carry_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__0_carry_i_6__1
       (.I0(n14__56_carry_0[1]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[2]),
        .I3(n4[0]),
        .O(n17__0_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__0_carry_i_7__1
       (.I0(n14__56_carry_0[0]),
        .I1(n4[1]),
        .O(n17__0_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n17__0_carry_i_8__1
       (.I0(n17__0_carry_i_1__1_n_0),
        .I1(n14__56_carry_0[1]),
        .I2(n4[6]),
        .I3(n17__0_carry_i_16__1_n_0),
        .I4(n4[7]),
        .I5(n14__56_carry_0[0]),
        .O(n17__0_carry_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__0_carry_i_9__1
       (.I0(n17__0_carry_i_2__1_n_0),
        .I1(n14__56_carry_0[1]),
        .I2(n4[5]),
        .I3(n17__0_carry_i_17__1_n_0),
        .I4(n4[6]),
        .I5(n14__56_carry_0[0]),
        .O(n17__0_carry_i_9__1_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__27_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n17__27_carry_n_0,n17__27_carry_n_1,n17__27_carry_n_2,n17__27_carry_n_3,n17__27_carry_n_4,n17__27_carry_n_5,n17__27_carry_n_6,n17__27_carry_n_7}),
        .DI({n17__27_carry_i_1__1_n_0,n17__27_carry_i_2__1_n_0,n17__27_carry_i_3__1_n_0,n17__27_carry_i_4__1_n_0,n17__27_carry_i_5__1_n_0,n17__27_carry_i_6__1_n_0,n17__27_carry_i_7__1_n_0,1'b0}),
        .O({n17__27_carry_n_8,n17__27_carry_n_9,n17__27_carry_n_10,n17__27_carry_n_11,n17__27_carry_n_12,n17__27_carry_n_13,n17__27_carry_n_14,n17__27_carry_n_15}),
        .S({n17__27_carry_i_8__1_n_0,n17__27_carry_i_9__1_n_0,n17__27_carry_i_10__1_n_0,n17__27_carry_i_11__1_n_0,n17__27_carry_i_12__1_n_0,n17__27_carry_i_13__1_n_0,n17__27_carry_i_14__1_n_0,n17__27_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__27_carry__0
       (.CI(n17__27_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n17__27_carry__0_CO_UNCONNECTED[7:3],n17__27_carry__0_n_5,NLW_n17__27_carry__0_CO_UNCONNECTED[1],n17__27_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n17__27_carry__0_i_1__1_n_0,n17__27_carry__0_i_2__1_n_0}),
        .O({NLW_n17__27_carry__0_O_UNCONNECTED[7:2],n17__27_carry__0_n_14,n17__27_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n17__27_carry__0_i_3__1_n_0,n17__27_carry__0_i_4__1_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__27_carry__0_i_1__1
       (.I0(n14__56_carry_0[4]),
        .I1(n4[7]),
        .I2(n14__56_carry_0[5]),
        .I3(n4[6]),
        .O(n17__27_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n17__27_carry__0_i_2__1
       (.I0(n14__56_carry_0[5]),
        .I1(n4[5]),
        .I2(n14__56_carry_0[4]),
        .I3(n4[6]),
        .I4(n14__56_carry_0[3]),
        .I5(n4[7]),
        .O(n17__27_carry__0_i_2__1_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n17__27_carry__0_i_3__1
       (.I0(n4[6]),
        .I1(n14__56_carry_0[4]),
        .I2(n14__56_carry_0[5]),
        .I3(n4[7]),
        .O(n17__27_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n17__27_carry__0_i_4__1
       (.I0(n14__56_carry_0[3]),
        .I1(n4[5]),
        .I2(n4[6]),
        .I3(n14__56_carry_0[5]),
        .I4(n4[7]),
        .I5(n14__56_carry_0[4]),
        .O(n17__27_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__27_carry_i_10__1
       (.I0(n17__27_carry_i_3__1_n_0),
        .I1(n14__56_carry_0[4]),
        .I2(n4[4]),
        .I3(n17__27_carry_i_18__1_n_0),
        .I4(n4[5]),
        .I5(n14__56_carry_0[3]),
        .O(n17__27_carry_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__27_carry_i_11__1
       (.I0(n17__27_carry_i_4__1_n_0),
        .I1(n14__56_carry_0[4]),
        .I2(n4[3]),
        .I3(n17__27_carry_i_19__1_n_0),
        .I4(n4[4]),
        .I5(n14__56_carry_0[3]),
        .O(n17__27_carry_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n17__27_carry_i_12__1
       (.I0(n4[2]),
        .I1(n17__27_carry_i_20__1_n_0),
        .I2(n4[1]),
        .I3(n14__56_carry_0[4]),
        .I4(n4[0]),
        .I5(n14__56_carry_0[5]),
        .O(n17__27_carry_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n17__27_carry_i_13__1
       (.I0(n4[0]),
        .I1(n14__56_carry_0[5]),
        .I2(n4[1]),
        .I3(n14__56_carry_0[4]),
        .I4(n14__56_carry_0[3]),
        .I5(n4[2]),
        .O(n17__27_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__27_carry_i_14__1
       (.I0(n14__56_carry_0[3]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[4]),
        .I3(n4[0]),
        .O(n17__27_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__27_carry_i_15__1
       (.I0(n4[0]),
        .I1(n14__56_carry_0[3]),
        .O(n17__27_carry_i_15__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_16__1
       (.I0(n4[5]),
        .I1(n14__56_carry_0[5]),
        .O(n17__27_carry_i_16__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_17__1
       (.I0(n4[4]),
        .I1(n14__56_carry_0[5]),
        .O(n17__27_carry_i_17__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_18__1
       (.I0(n4[3]),
        .I1(n14__56_carry_0[5]),
        .O(n17__27_carry_i_18__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_19__1
       (.I0(n4[2]),
        .I1(n14__56_carry_0[5]),
        .O(n17__27_carry_i_19__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__27_carry_i_1__1
       (.I0(n14__56_carry_0[5]),
        .I1(n4[4]),
        .I2(n14__56_carry_0[4]),
        .I3(n4[5]),
        .I4(n14__56_carry_0[3]),
        .I5(n4[6]),
        .O(n17__27_carry_i_1__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_20__1
       (.I0(n4[3]),
        .I1(n14__56_carry_0[3]),
        .O(n17__27_carry_i_20__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__27_carry_i_2__1
       (.I0(n14__56_carry_0[5]),
        .I1(n4[3]),
        .I2(n14__56_carry_0[4]),
        .I3(n4[4]),
        .I4(n14__56_carry_0[3]),
        .I5(n4[5]),
        .O(n17__27_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__27_carry_i_3__1
       (.I0(n14__56_carry_0[5]),
        .I1(n4[2]),
        .I2(n14__56_carry_0[4]),
        .I3(n4[3]),
        .I4(n14__56_carry_0[3]),
        .I5(n4[4]),
        .O(n17__27_carry_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__27_carry_i_4__1
       (.I0(n14__56_carry_0[5]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[4]),
        .I3(n4[2]),
        .I4(n14__56_carry_0[3]),
        .I5(n4[3]),
        .O(n17__27_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n17__27_carry_i_5__1
       (.I0(n14__56_carry_0[4]),
        .I1(n4[2]),
        .I2(n14__56_carry_0[5]),
        .I3(n4[1]),
        .I4(n4[3]),
        .I5(n14__56_carry_0[3]),
        .O(n17__27_carry_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__27_carry_i_6__1
       (.I0(n14__56_carry_0[4]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[5]),
        .I3(n4[0]),
        .O(n17__27_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__27_carry_i_7__1
       (.I0(n14__56_carry_0[3]),
        .I1(n4[1]),
        .O(n17__27_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n17__27_carry_i_8__1
       (.I0(n17__27_carry_i_1__1_n_0),
        .I1(n14__56_carry_0[4]),
        .I2(n4[6]),
        .I3(n17__27_carry_i_16__1_n_0),
        .I4(n4[7]),
        .I5(n14__56_carry_0[3]),
        .O(n17__27_carry_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__27_carry_i_9__1
       (.I0(n17__27_carry_i_2__1_n_0),
        .I1(n14__56_carry_0[4]),
        .I2(n4[5]),
        .I3(n17__27_carry_i_17__1_n_0),
        .I4(n4[6]),
        .I5(n14__56_carry_0[3]),
        .O(n17__27_carry_i_9__1_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__56_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n17__56_carry_n_0,n17__56_carry_n_1,n17__56_carry_n_2,n17__56_carry_n_3,n17__56_carry_n_4,n17__56_carry_n_5,n17__56_carry_n_6,n17__56_carry_n_7}),
        .DI({n17__56_carry_i_1__1_n_0,n17__56_carry_i_2__1_n_0,n17__56_carry_i_3__1_n_0,n17__56_carry_i_4__1_n_0,n17__56_carry_i_5__1_n_0,n17__56_carry_i_6__1_n_0,n17__56_carry_i_7__1_n_0,1'b0}),
        .O({n17__56_carry_n_8,n17__56_carry_n_9,n17__56_carry_n_10,n17__56_carry_n_11,n17__56_carry_n_12,n17__56_carry_n_13,n17__56_carry_n_14,n17__56_carry_n_15}),
        .S({n17__56_carry_i_8__1_n_0,n17__56_carry_i_9__1_n_0,n17__56_carry_i_10__1_n_0,n17__56_carry_i_11__1_n_0,n17__56_carry_i_12__1_n_0,n17__56_carry_i_13__1_n_0,n17__56_carry_i_14__1_n_0,n17__56_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__56_carry__0
       (.CI(n17__56_carry_n_0),
        .CI_TOP(1'b0),
        .CO(NLW_n17__56_carry__0_CO_UNCONNECTED[7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_n17__56_carry__0_O_UNCONNECTED[7:1],n17__56_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n17__56_carry__0_i_1__1_n_0}));
  LUT4 #(
    .INIT(16'hE53F)) 
    n17__56_carry__0_i_1__1
       (.I0(n14__56_carry_0[6]),
        .I1(n4[6]),
        .I2(n14__56_carry_0[7]),
        .I3(n4[7]),
        .O(n17__56_carry__0_i_1__1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n17__56_carry_i_10__1
       (.I0(n4[3]),
        .I1(n4[4]),
        .I2(n14__56_carry_0[7]),
        .I3(n4[5]),
        .I4(n14__56_carry_0[6]),
        .O(n17__56_carry_i_10__1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n17__56_carry_i_11__1
       (.I0(n4[2]),
        .I1(n4[3]),
        .I2(n14__56_carry_0[7]),
        .I3(n4[4]),
        .I4(n14__56_carry_0[6]),
        .O(n17__56_carry_i_11__1_n_0));
  LUT5 #(
    .INIT(32'h9F606060)) 
    n17__56_carry_i_12__1
       (.I0(n4[1]),
        .I1(n4[2]),
        .I2(n14__56_carry_0[7]),
        .I3(n4[3]),
        .I4(n14__56_carry_0[6]),
        .O(n17__56_carry_i_12__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__56_carry_i_13__1
       (.I0(n14__56_carry_0[7]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[6]),
        .I3(n4[2]),
        .O(n17__56_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h8777)) 
    n17__56_carry_i_14__1
       (.I0(n14__56_carry_0[7]),
        .I1(n4[0]),
        .I2(n14__56_carry_0[6]),
        .I3(n4[1]),
        .O(n17__56_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__56_carry_i_15__1
       (.I0(n4[0]),
        .I1(n14__56_carry_0[6]),
        .O(n17__56_carry_i_15__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__56_carry_i_1__1
       (.I0(n14__56_carry_0[7]),
        .I1(n4[5]),
        .I2(n14__56_carry_0[6]),
        .I3(n4[6]),
        .O(n17__56_carry_i_1__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__56_carry_i_2__1
       (.I0(n14__56_carry_0[7]),
        .I1(n4[4]),
        .I2(n14__56_carry_0[6]),
        .I3(n4[5]),
        .O(n17__56_carry_i_2__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__56_carry_i_3__1
       (.I0(n14__56_carry_0[7]),
        .I1(n4[3]),
        .I2(n14__56_carry_0[6]),
        .I3(n4[4]),
        .O(n17__56_carry_i_3__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__56_carry_i_4__1
       (.I0(n14__56_carry_0[7]),
        .I1(n4[2]),
        .I2(n14__56_carry_0[6]),
        .I3(n4[3]),
        .O(n17__56_carry_i_4__1_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n17__56_carry_i_5__1
       (.I0(n4[1]),
        .I1(n14__56_carry_0[7]),
        .O(n17__56_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__56_carry_i_6__1
       (.I0(n14__56_carry_0[7]),
        .I1(n4[1]),
        .O(n17__56_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n17__56_carry_i_7__1
       (.I0(n4[0]),
        .I1(n14__56_carry_0[7]),
        .O(n17__56_carry_i_7__1_n_0));
  LUT5 #(
    .INIT(32'h738CC0C0)) 
    n17__56_carry_i_8__1
       (.I0(n4[5]),
        .I1(n4[6]),
        .I2(n14__56_carry_0[7]),
        .I3(n4[7]),
        .I4(n14__56_carry_0[6]),
        .O(n17__56_carry_i_8__1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n17__56_carry_i_9__1
       (.I0(n4[4]),
        .I1(n4[5]),
        .I2(n14__56_carry_0[7]),
        .I3(n4[6]),
        .I4(n14__56_carry_0[6]),
        .O(n17__56_carry_i_9__1_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__81_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n17__81_carry_n_0,n17__81_carry_n_1,n17__81_carry_n_2,n17__81_carry_n_3,n17__81_carry_n_4,n17__81_carry_n_5,n17__81_carry_n_6,n17__81_carry_n_7}),
        .DI({n17__81_carry_i_1__1_n_0,n17__81_carry_i_2__1_n_0,n17__81_carry_i_3__1_n_0,n17__81_carry_i_4__1_n_0,n17__81_carry_i_5__1_n_0,n17__81_carry_i_6__1_n_0,n17__81_carry_i_7__1_n_0,1'b0}),
        .O({n17[10:7],NLW_n17__81_carry_O_UNCONNECTED[3:0]}),
        .S({n17__81_carry_i_8__1_n_0,n17__81_carry_i_9__1_n_0,n17__81_carry_i_10__1_n_0,n17__81_carry_i_11__1_n_0,n17__81_carry_i_12__1_n_0,n17__81_carry_i_13__1_n_0,n17__81_carry_i_14__1_n_0,n17__81_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__81_carry__0
       (.CI(n17__81_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n17__81_carry__0_CO_UNCONNECTED[7:3],n17__81_carry__0_n_5,n17__81_carry__0_n_6,n17__81_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n17__81_carry__0_i_1__1_n_0,n17__81_carry__0_i_2__1_n_0,n17__81_carry__0_i_3__1_n_0}),
        .O({NLW_n17__81_carry__0_O_UNCONNECTED[7:4],n17[14:11]}),
        .S({1'b0,1'b0,1'b0,1'b0,n17__81_carry__0_i_4__1_n_0,n17__81_carry__0_i_5__1_n_0,n17__81_carry__0_i_6__1_n_0,n17__81_carry__0_i_7__1_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry__0_i_1__1
       (.I0(n17__27_carry__0_n_14),
        .I1(n17__56_carry_n_9),
        .O(n17__81_carry__0_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry__0_i_2__1
       (.I0(n17__27_carry__0_n_15),
        .I1(n17__56_carry_n_10),
        .O(n17__81_carry__0_i_2__1_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry__0_i_3__1
       (.I0(n17__56_carry_n_11),
        .I1(n17__27_carry_n_8),
        .I2(n17__0_carry__0_n_5),
        .O(n17__81_carry__0_i_3__1_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n17__81_carry__0_i_4__1
       (.I0(n17__27_carry__0_n_5),
        .I1(n17__56_carry_n_8),
        .I2(n17__56_carry__0_n_15),
        .O(n17__81_carry__0_i_4__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n17__81_carry__0_i_5__1
       (.I0(n17__27_carry__0_n_14),
        .I1(n17__56_carry_n_9),
        .I2(n17__56_carry_n_8),
        .I3(n17__27_carry__0_n_5),
        .O(n17__81_carry__0_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n17__81_carry__0_i_6__1
       (.I0(n17__27_carry__0_n_15),
        .I1(n17__56_carry_n_10),
        .I2(n17__56_carry_n_9),
        .I3(n17__27_carry__0_n_14),
        .O(n17__81_carry__0_i_6__1_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n17__81_carry__0_i_7__1
       (.I0(n17__0_carry__0_n_5),
        .I1(n17__27_carry_n_8),
        .I2(n17__56_carry_n_11),
        .I3(n17__56_carry_n_10),
        .I4(n17__27_carry__0_n_15),
        .O(n17__81_carry__0_i_7__1_n_0));
  (* HLUTNM = "lutpair26" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_10__1
       (.I0(n17__56_carry_n_13),
        .I1(n17__27_carry_n_10),
        .I2(n17__0_carry__0_n_15),
        .I3(n17__81_carry_i_3__1_n_0),
        .O(n17__81_carry_i_10__1_n_0));
  (* HLUTNM = "lutpair25" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_11__1
       (.I0(n17__56_carry_n_14),
        .I1(n17__27_carry_n_11),
        .I2(n17__0_carry_n_8),
        .I3(n17__81_carry_i_4__1_n_0),
        .O(n17__81_carry_i_11__1_n_0));
  (* HLUTNM = "lutpair24" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_12__1
       (.I0(n17__56_carry_n_15),
        .I1(n17__27_carry_n_12),
        .I2(n17__0_carry_n_9),
        .I3(n17__81_carry_i_5__1_n_0),
        .O(n17__81_carry_i_12__1_n_0));
  (* HLUTNM = "lutpair86" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n17__81_carry_i_13__1
       (.I0(n17__27_carry_n_13),
        .I1(n17__0_carry_n_10),
        .I2(n17__0_carry_n_11),
        .I3(n17__27_carry_n_14),
        .O(n17__81_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n17__81_carry_i_14__1
       (.I0(n17__0_carry_n_12),
        .I1(n17__27_carry_n_15),
        .I2(n17__27_carry_n_14),
        .I3(n17__0_carry_n_11),
        .O(n17__81_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n17__81_carry_i_15__1
       (.I0(n17__0_carry_n_12),
        .I1(n17__27_carry_n_15),
        .O(n17__81_carry_i_15__1_n_0));
  (* HLUTNM = "lutpair27" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry_i_1__1
       (.I0(n17__56_carry_n_12),
        .I1(n17__27_carry_n_9),
        .I2(n17__0_carry__0_n_14),
        .O(n17__81_carry_i_1__1_n_0));
  (* HLUTNM = "lutpair26" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry_i_2__1
       (.I0(n17__56_carry_n_13),
        .I1(n17__27_carry_n_10),
        .I2(n17__0_carry__0_n_15),
        .O(n17__81_carry_i_2__1_n_0));
  (* HLUTNM = "lutpair25" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry_i_3__1
       (.I0(n17__56_carry_n_14),
        .I1(n17__27_carry_n_11),
        .I2(n17__0_carry_n_8),
        .O(n17__81_carry_i_3__1_n_0));
  (* HLUTNM = "lutpair24" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry_i_4__1
       (.I0(n17__56_carry_n_15),
        .I1(n17__27_carry_n_12),
        .I2(n17__0_carry_n_9),
        .O(n17__81_carry_i_4__1_n_0));
  (* HLUTNM = "lutpair86" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry_i_5__1
       (.I0(n17__27_carry_n_13),
        .I1(n17__0_carry_n_10),
        .O(n17__81_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry_i_6__1
       (.I0(n17__0_carry_n_11),
        .I1(n17__27_carry_n_14),
        .O(n17__81_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry_i_7__1
       (.I0(n17__0_carry_n_12),
        .I1(n17__27_carry_n_15),
        .O(n17__81_carry_i_7__1_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_8__1
       (.I0(n17__81_carry_i_1__1_n_0),
        .I1(n17__27_carry_n_8),
        .I2(n17__56_carry_n_11),
        .I3(n17__0_carry__0_n_5),
        .O(n17__81_carry_i_8__1_n_0));
  (* HLUTNM = "lutpair27" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_9__1
       (.I0(n17__56_carry_n_12),
        .I1(n17__27_carry_n_9),
        .I2(n17__0_carry__0_n_14),
        .I3(n17__81_carry_i_2__1_n_0),
        .O(n17__81_carry_i_9__1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[14]),
        .Q(n19_reg_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__0
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[13]),
        .Q(n19_reg__0_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__1
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[12]),
        .Q(n19_reg__1_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__2
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[11]),
        .Q(n19_reg__2_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__3
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[10]),
        .Q(n19_reg__3_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__4
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[9]),
        .Q(n19_reg__4_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__5
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[8]),
        .Q(n19_reg__5_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__6
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[7]),
        .Q(n19_reg__6_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[0]),
        .Q(\n1_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[10]),
        .Q(n2[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[11]),
        .Q(n2[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[12]),
        .Q(n2[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[13]),
        .Q(n2[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[14]),
        .Q(n2[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[15]),
        .Q(n2[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[1]),
        .Q(\n1_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[2]),
        .Q(\n1_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[3]),
        .Q(\n1_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[4]),
        .Q(\n1_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[5]),
        .Q(\n1_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[6]),
        .Q(\n1_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[7]),
        .Q(\n1_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[8]),
        .Q(n2[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[9]),
        .Q(n2[1]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n20_carry
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({NLW_n20_carry_CO_UNCONNECTED[7],n20_carry_n_1,n20_carry_n_2,n20_carry_n_3,n20_carry_n_4,n20_carry_n_5,n20_carry_n_6,n20_carry_n_7}),
        .DI({1'b0,\n16_reg_n_0_[6] ,\n16_reg_n_0_[5] ,\n16_reg_n_0_[4] ,\n16_reg_n_0_[3] ,\n16_reg_n_0_[2] ,\n16_reg_n_0_[1] ,\n16_reg_n_0_[0] }),
        .O(n202_out),
        .S({n20_carry_i_1__2_n_0,n20_carry_i_2__2_n_0,n20_carry_i_3__2_n_0,n20_carry_i_4__2_n_0,n20_carry_i_5__2_n_0,n20_carry_i_6__2_n_0,n20_carry_i_7__2_n_0,n20_carry_i_8__2_n_0}));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_1__2
       (.I0(\n16_reg_n_0_[7] ),
        .I1(n19_reg_n_0),
        .O(n20_carry_i_1__2_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_2__2
       (.I0(\n16_reg_n_0_[6] ),
        .I1(n19_reg__0_n_0),
        .O(n20_carry_i_2__2_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_3__2
       (.I0(\n16_reg_n_0_[5] ),
        .I1(n19_reg__1_n_0),
        .O(n20_carry_i_3__2_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_4__2
       (.I0(\n16_reg_n_0_[4] ),
        .I1(n19_reg__2_n_0),
        .O(n20_carry_i_4__2_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_5__2
       (.I0(\n16_reg_n_0_[3] ),
        .I1(n19_reg__3_n_0),
        .O(n20_carry_i_5__2_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_6__2
       (.I0(\n16_reg_n_0_[2] ),
        .I1(n19_reg__4_n_0),
        .O(n20_carry_i_6__2_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_7__2
       (.I0(\n16_reg_n_0_[1] ),
        .I1(n19_reg__5_n_0),
        .O(n20_carry_i_7__2_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_8__2
       (.I0(\n16_reg_n_0_[0] ),
        .I1(n19_reg__6_n_0),
        .O(n20_carry_i_8__2_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[0]),
        .Q(n21[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[1]),
        .Q(n21[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[2]),
        .Q(n21[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[3]),
        .Q(n21[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[4]),
        .Q(n21[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[5]),
        .Q(n21[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[6]),
        .Q(n21[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[7]),
        .Q(n21[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[15]),
        .Q(n22_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__0
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[14]),
        .Q(n22__0_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__0_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n22__0_carry_n_0,n22__0_carry_n_1,n22__0_carry_n_2,n22__0_carry_n_3,n22__0_carry_n_4,n22__0_carry_n_5,n22__0_carry_n_6,n22__0_carry_n_7}),
        .DI({n22__0_carry_i_1__1_n_0,n22__0_carry_i_2__1_n_0,n22__0_carry_i_3__1_n_0,n22__0_carry_i_4__1_n_0,n22__0_carry_i_5__1_n_0,n22__0_carry_i_6__1_n_0,n22__0_carry_i_7__1_n_0,1'b0}),
        .O({n22__0_carry_n_8,n22__0_carry_n_9,n22__0_carry_n_10,n22__0_carry_n_11,n22__0_carry_n_12,NLW_n22__0_carry_O_UNCONNECTED[2:0]}),
        .S({n22__0_carry_i_8__1_n_0,n22__0_carry_i_9__1_n_0,n22__0_carry_i_10__1_n_0,n22__0_carry_i_11__1_n_0,n22__0_carry_i_12__1_n_0,n22__0_carry_i_13__1_n_0,n22__0_carry_i_14__1_n_0,n22__0_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__0_carry__0
       (.CI(n22__0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n22__0_carry__0_CO_UNCONNECTED[7:3],n22__0_carry__0_n_5,NLW_n22__0_carry__0_CO_UNCONNECTED[1],n22__0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n22__0_carry__0_i_1__1_n_0,n22__0_carry__0_i_2__1_n_0}),
        .O({NLW_n22__0_carry__0_O_UNCONNECTED[7:2],n22__0_carry__0_n_14,n22__0_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n22__0_carry__0_i_3__1_n_0,n22__0_carry__0_i_4__1_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__0_carry__0_i_1__1
       (.I0(n14__56_carry_0[1]),
        .I1(n22_n_0),
        .I2(n14__56_carry_0[2]),
        .I3(n22__0_n_0),
        .O(n22__0_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n22__0_carry__0_i_2__1
       (.I0(n14__56_carry_0[2]),
        .I1(n22__1_n_0),
        .I2(n14__56_carry_0[1]),
        .I3(n22__0_n_0),
        .I4(n14__56_carry_0[0]),
        .I5(n22_n_0),
        .O(n22__0_carry__0_i_2__1_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n22__0_carry__0_i_3__1
       (.I0(n22__0_n_0),
        .I1(n14__56_carry_0[1]),
        .I2(n14__56_carry_0[2]),
        .I3(n22_n_0),
        .O(n22__0_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n22__0_carry__0_i_4__1
       (.I0(n14__56_carry_0[0]),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(n14__56_carry_0[2]),
        .I4(n22_n_0),
        .I5(n14__56_carry_0[1]),
        .O(n22__0_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__0_carry_i_10__1
       (.I0(n22__0_carry_i_3__1_n_0),
        .I1(n14__56_carry_0[1]),
        .I2(n22__2_n_0),
        .I3(n22__0_carry_i_18__1_n_0),
        .I4(n22__1_n_0),
        .I5(n14__56_carry_0[0]),
        .O(n22__0_carry_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__0_carry_i_11__1
       (.I0(n22__0_carry_i_4__1_n_0),
        .I1(n14__56_carry_0[1]),
        .I2(n22__3_n_0),
        .I3(n22__0_carry_i_19__1_n_0),
        .I4(n22__2_n_0),
        .I5(n14__56_carry_0[0]),
        .O(n22__0_carry_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n22__0_carry_i_12__1
       (.I0(n22__4_n_0),
        .I1(n22__0_carry_i_20__1_n_0),
        .I2(n22__5_n_0),
        .I3(n14__56_carry_0[1]),
        .I4(n22__6_n_0),
        .I5(n14__56_carry_0[2]),
        .O(n22__0_carry_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n22__0_carry_i_13__1
       (.I0(n22__6_n_0),
        .I1(n14__56_carry_0[2]),
        .I2(n22__5_n_0),
        .I3(n14__56_carry_0[1]),
        .I4(n14__56_carry_0[0]),
        .I5(n22__4_n_0),
        .O(n22__0_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__0_carry_i_14__1
       (.I0(n14__56_carry_0[0]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[1]),
        .I3(n22__6_n_0),
        .O(n22__0_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__0_carry_i_15__1
       (.I0(n22__6_n_0),
        .I1(n14__56_carry_0[0]),
        .O(n22__0_carry_i_15__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_16__1
       (.I0(n22__1_n_0),
        .I1(n14__56_carry_0[2]),
        .O(n22__0_carry_i_16__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_17__1
       (.I0(n22__2_n_0),
        .I1(n14__56_carry_0[2]),
        .O(n22__0_carry_i_17__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_18__1
       (.I0(n22__3_n_0),
        .I1(n14__56_carry_0[2]),
        .O(n22__0_carry_i_18__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_19__1
       (.I0(n22__4_n_0),
        .I1(n14__56_carry_0[2]),
        .O(n22__0_carry_i_19__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__0_carry_i_1__1
       (.I0(n14__56_carry_0[2]),
        .I1(n22__2_n_0),
        .I2(n14__56_carry_0[1]),
        .I3(n22__1_n_0),
        .I4(n14__56_carry_0[0]),
        .I5(n22__0_n_0),
        .O(n22__0_carry_i_1__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_20__1
       (.I0(n22__3_n_0),
        .I1(n14__56_carry_0[0]),
        .O(n22__0_carry_i_20__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__0_carry_i_2__1
       (.I0(n14__56_carry_0[2]),
        .I1(n22__3_n_0),
        .I2(n14__56_carry_0[1]),
        .I3(n22__2_n_0),
        .I4(n14__56_carry_0[0]),
        .I5(n22__1_n_0),
        .O(n22__0_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__0_carry_i_3__1
       (.I0(n14__56_carry_0[2]),
        .I1(n22__4_n_0),
        .I2(n14__56_carry_0[1]),
        .I3(n22__3_n_0),
        .I4(n14__56_carry_0[0]),
        .I5(n22__2_n_0),
        .O(n22__0_carry_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__0_carry_i_4__1
       (.I0(n14__56_carry_0[2]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[1]),
        .I3(n22__4_n_0),
        .I4(n14__56_carry_0[0]),
        .I5(n22__3_n_0),
        .O(n22__0_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n22__0_carry_i_5__1
       (.I0(n14__56_carry_0[1]),
        .I1(n22__4_n_0),
        .I2(n14__56_carry_0[2]),
        .I3(n22__5_n_0),
        .I4(n22__3_n_0),
        .I5(n14__56_carry_0[0]),
        .O(n22__0_carry_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__0_carry_i_6__1
       (.I0(n14__56_carry_0[1]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[2]),
        .I3(n22__6_n_0),
        .O(n22__0_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__0_carry_i_7__1
       (.I0(n14__56_carry_0[0]),
        .I1(n22__5_n_0),
        .O(n22__0_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n22__0_carry_i_8__1
       (.I0(n22__0_carry_i_1__1_n_0),
        .I1(n14__56_carry_0[1]),
        .I2(n22__0_n_0),
        .I3(n22__0_carry_i_16__1_n_0),
        .I4(n22_n_0),
        .I5(n14__56_carry_0[0]),
        .O(n22__0_carry_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__0_carry_i_9__1
       (.I0(n22__0_carry_i_2__1_n_0),
        .I1(n14__56_carry_0[1]),
        .I2(n22__1_n_0),
        .I3(n22__0_carry_i_17__1_n_0),
        .I4(n22__0_n_0),
        .I5(n14__56_carry_0[0]),
        .O(n22__0_carry_i_9__1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    n22__1
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[13]),
        .Q(n22__1_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__2
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[12]),
        .Q(n22__2_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__27_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n22__27_carry_n_0,n22__27_carry_n_1,n22__27_carry_n_2,n22__27_carry_n_3,n22__27_carry_n_4,n22__27_carry_n_5,n22__27_carry_n_6,n22__27_carry_n_7}),
        .DI({n22__27_carry_i_1__1_n_0,n22__27_carry_i_2__1_n_0,n22__27_carry_i_3__1_n_0,n22__27_carry_i_4__1_n_0,n22__27_carry_i_5__1_n_0,n22__27_carry_i_6__1_n_0,n22__27_carry_i_7__1_n_0,1'b0}),
        .O({n22__27_carry_n_8,n22__27_carry_n_9,n22__27_carry_n_10,n22__27_carry_n_11,n22__27_carry_n_12,n22__27_carry_n_13,n22__27_carry_n_14,n22__27_carry_n_15}),
        .S({n22__27_carry_i_8__1_n_0,n22__27_carry_i_9__1_n_0,n22__27_carry_i_10__1_n_0,n22__27_carry_i_11__1_n_0,n22__27_carry_i_12__1_n_0,n22__27_carry_i_13__1_n_0,n22__27_carry_i_14__1_n_0,n22__27_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__27_carry__0
       (.CI(n22__27_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n22__27_carry__0_CO_UNCONNECTED[7:3],n22__27_carry__0_n_5,NLW_n22__27_carry__0_CO_UNCONNECTED[1],n22__27_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n22__27_carry__0_i_1__1_n_0,n22__27_carry__0_i_2__1_n_0}),
        .O({NLW_n22__27_carry__0_O_UNCONNECTED[7:2],n22__27_carry__0_n_14,n22__27_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n22__27_carry__0_i_3__1_n_0,n22__27_carry__0_i_4__1_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__27_carry__0_i_1__1
       (.I0(n14__56_carry_0[4]),
        .I1(n22_n_0),
        .I2(n14__56_carry_0[5]),
        .I3(n22__0_n_0),
        .O(n22__27_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n22__27_carry__0_i_2__1
       (.I0(n14__56_carry_0[5]),
        .I1(n22__1_n_0),
        .I2(n14__56_carry_0[4]),
        .I3(n22__0_n_0),
        .I4(n14__56_carry_0[3]),
        .I5(n22_n_0),
        .O(n22__27_carry__0_i_2__1_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n22__27_carry__0_i_3__1
       (.I0(n22__0_n_0),
        .I1(n14__56_carry_0[4]),
        .I2(n14__56_carry_0[5]),
        .I3(n22_n_0),
        .O(n22__27_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n22__27_carry__0_i_4__1
       (.I0(n14__56_carry_0[3]),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(n14__56_carry_0[5]),
        .I4(n22_n_0),
        .I5(n14__56_carry_0[4]),
        .O(n22__27_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__27_carry_i_10__1
       (.I0(n22__27_carry_i_3__1_n_0),
        .I1(n14__56_carry_0[4]),
        .I2(n22__2_n_0),
        .I3(n22__27_carry_i_18__1_n_0),
        .I4(n22__1_n_0),
        .I5(n14__56_carry_0[3]),
        .O(n22__27_carry_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__27_carry_i_11__1
       (.I0(n22__27_carry_i_4__1_n_0),
        .I1(n14__56_carry_0[4]),
        .I2(n22__3_n_0),
        .I3(n22__27_carry_i_19__1_n_0),
        .I4(n22__2_n_0),
        .I5(n14__56_carry_0[3]),
        .O(n22__27_carry_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n22__27_carry_i_12__1
       (.I0(n22__4_n_0),
        .I1(n22__27_carry_i_20__1_n_0),
        .I2(n22__5_n_0),
        .I3(n14__56_carry_0[4]),
        .I4(n22__6_n_0),
        .I5(n14__56_carry_0[5]),
        .O(n22__27_carry_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n22__27_carry_i_13__1
       (.I0(n22__6_n_0),
        .I1(n14__56_carry_0[5]),
        .I2(n22__5_n_0),
        .I3(n14__56_carry_0[4]),
        .I4(n14__56_carry_0[3]),
        .I5(n22__4_n_0),
        .O(n22__27_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__27_carry_i_14__1
       (.I0(n14__56_carry_0[3]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[4]),
        .I3(n22__6_n_0),
        .O(n22__27_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__27_carry_i_15__1
       (.I0(n22__6_n_0),
        .I1(n14__56_carry_0[3]),
        .O(n22__27_carry_i_15__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_16__1
       (.I0(n22__1_n_0),
        .I1(n14__56_carry_0[5]),
        .O(n22__27_carry_i_16__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_17__1
       (.I0(n22__2_n_0),
        .I1(n14__56_carry_0[5]),
        .O(n22__27_carry_i_17__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_18__1
       (.I0(n22__3_n_0),
        .I1(n14__56_carry_0[5]),
        .O(n22__27_carry_i_18__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_19__1
       (.I0(n22__4_n_0),
        .I1(n14__56_carry_0[5]),
        .O(n22__27_carry_i_19__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__27_carry_i_1__1
       (.I0(n14__56_carry_0[5]),
        .I1(n22__2_n_0),
        .I2(n14__56_carry_0[4]),
        .I3(n22__1_n_0),
        .I4(n14__56_carry_0[3]),
        .I5(n22__0_n_0),
        .O(n22__27_carry_i_1__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_20__1
       (.I0(n22__3_n_0),
        .I1(n14__56_carry_0[3]),
        .O(n22__27_carry_i_20__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__27_carry_i_2__1
       (.I0(n14__56_carry_0[5]),
        .I1(n22__3_n_0),
        .I2(n14__56_carry_0[4]),
        .I3(n22__2_n_0),
        .I4(n14__56_carry_0[3]),
        .I5(n22__1_n_0),
        .O(n22__27_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__27_carry_i_3__1
       (.I0(n14__56_carry_0[5]),
        .I1(n22__4_n_0),
        .I2(n14__56_carry_0[4]),
        .I3(n22__3_n_0),
        .I4(n14__56_carry_0[3]),
        .I5(n22__2_n_0),
        .O(n22__27_carry_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__27_carry_i_4__1
       (.I0(n14__56_carry_0[5]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[4]),
        .I3(n22__4_n_0),
        .I4(n14__56_carry_0[3]),
        .I5(n22__3_n_0),
        .O(n22__27_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n22__27_carry_i_5__1
       (.I0(n14__56_carry_0[4]),
        .I1(n22__4_n_0),
        .I2(n14__56_carry_0[5]),
        .I3(n22__5_n_0),
        .I4(n22__3_n_0),
        .I5(n14__56_carry_0[3]),
        .O(n22__27_carry_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__27_carry_i_6__1
       (.I0(n14__56_carry_0[4]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[5]),
        .I3(n22__6_n_0),
        .O(n22__27_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__27_carry_i_7__1
       (.I0(n14__56_carry_0[3]),
        .I1(n22__5_n_0),
        .O(n22__27_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n22__27_carry_i_8__1
       (.I0(n22__27_carry_i_1__1_n_0),
        .I1(n14__56_carry_0[4]),
        .I2(n22__0_n_0),
        .I3(n22__27_carry_i_16__1_n_0),
        .I4(n22_n_0),
        .I5(n14__56_carry_0[3]),
        .O(n22__27_carry_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__27_carry_i_9__1
       (.I0(n22__27_carry_i_2__1_n_0),
        .I1(n14__56_carry_0[4]),
        .I2(n22__1_n_0),
        .I3(n22__27_carry_i_17__1_n_0),
        .I4(n22__0_n_0),
        .I5(n14__56_carry_0[3]),
        .O(n22__27_carry_i_9__1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    n22__3
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[11]),
        .Q(n22__3_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__4
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[10]),
        .Q(n22__4_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__5
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[9]),
        .Q(n22__5_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__56_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n22__56_carry_n_0,n22__56_carry_n_1,n22__56_carry_n_2,n22__56_carry_n_3,n22__56_carry_n_4,n22__56_carry_n_5,n22__56_carry_n_6,n22__56_carry_n_7}),
        .DI({n22__56_carry_i_1__1_n_0,n22__56_carry_i_2__1_n_0,n22__56_carry_i_3__1_n_0,n22__56_carry_i_4__1_n_0,n22__56_carry_i_5__1_n_0,n22__56_carry_i_6__1_n_0,n22__56_carry_i_7__1_n_0,1'b0}),
        .O({n22__56_carry_n_8,n22__56_carry_n_9,n22__56_carry_n_10,n22__56_carry_n_11,n22__56_carry_n_12,n22__56_carry_n_13,n22__56_carry_n_14,n22__56_carry_n_15}),
        .S({n22__56_carry_i_8__1_n_0,n22__56_carry_i_9__1_n_0,n22__56_carry_i_10__1_n_0,n22__56_carry_i_11__1_n_0,n22__56_carry_i_12__1_n_0,n22__56_carry_i_13__1_n_0,n22__56_carry_i_14__1_n_0,n22__56_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__56_carry__0
       (.CI(n22__56_carry_n_0),
        .CI_TOP(1'b0),
        .CO(NLW_n22__56_carry__0_CO_UNCONNECTED[7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_n22__56_carry__0_O_UNCONNECTED[7:1],n22__56_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n22__56_carry__0_i_1__1_n_0}));
  LUT4 #(
    .INIT(16'hE53F)) 
    n22__56_carry__0_i_1__1
       (.I0(n14__56_carry_0[6]),
        .I1(n22__0_n_0),
        .I2(n14__56_carry_0[7]),
        .I3(n22_n_0),
        .O(n22__56_carry__0_i_1__1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n22__56_carry_i_10__1
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(n14__56_carry_0[7]),
        .I3(n22__1_n_0),
        .I4(n14__56_carry_0[6]),
        .O(n22__56_carry_i_10__1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n22__56_carry_i_11__1
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n14__56_carry_0[7]),
        .I3(n22__2_n_0),
        .I4(n14__56_carry_0[6]),
        .O(n22__56_carry_i_11__1_n_0));
  LUT5 #(
    .INIT(32'h9F606060)) 
    n22__56_carry_i_12__1
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(n14__56_carry_0[7]),
        .I3(n22__3_n_0),
        .I4(n14__56_carry_0[6]),
        .O(n22__56_carry_i_12__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__56_carry_i_13__1
       (.I0(n14__56_carry_0[7]),
        .I1(n22__5_n_0),
        .I2(n14__56_carry_0[6]),
        .I3(n22__4_n_0),
        .O(n22__56_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h8777)) 
    n22__56_carry_i_14__1
       (.I0(n14__56_carry_0[7]),
        .I1(n22__6_n_0),
        .I2(n14__56_carry_0[6]),
        .I3(n22__5_n_0),
        .O(n22__56_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__56_carry_i_15__1
       (.I0(n22__6_n_0),
        .I1(n14__56_carry_0[6]),
        .O(n22__56_carry_i_15__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__56_carry_i_1__1
       (.I0(n14__56_carry_0[7]),
        .I1(n22__1_n_0),
        .I2(n14__56_carry_0[6]),
        .I3(n22__0_n_0),
        .O(n22__56_carry_i_1__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__56_carry_i_2__1
       (.I0(n14__56_carry_0[7]),
        .I1(n22__2_n_0),
        .I2(n14__56_carry_0[6]),
        .I3(n22__1_n_0),
        .O(n22__56_carry_i_2__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__56_carry_i_3__1
       (.I0(n14__56_carry_0[7]),
        .I1(n22__3_n_0),
        .I2(n14__56_carry_0[6]),
        .I3(n22__2_n_0),
        .O(n22__56_carry_i_3__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__56_carry_i_4__1
       (.I0(n14__56_carry_0[7]),
        .I1(n22__4_n_0),
        .I2(n14__56_carry_0[6]),
        .I3(n22__3_n_0),
        .O(n22__56_carry_i_4__1_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n22__56_carry_i_5__1
       (.I0(n22__5_n_0),
        .I1(n14__56_carry_0[7]),
        .O(n22__56_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__56_carry_i_6__1
       (.I0(n14__56_carry_0[7]),
        .I1(n22__5_n_0),
        .O(n22__56_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n22__56_carry_i_7__1
       (.I0(n22__6_n_0),
        .I1(n14__56_carry_0[7]),
        .O(n22__56_carry_i_7__1_n_0));
  LUT5 #(
    .INIT(32'h738CC0C0)) 
    n22__56_carry_i_8__1
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n14__56_carry_0[7]),
        .I3(n22_n_0),
        .I4(n14__56_carry_0[6]),
        .O(n22__56_carry_i_8__1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n22__56_carry_i_9__1
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(n14__56_carry_0[7]),
        .I3(n22__0_n_0),
        .I4(n14__56_carry_0[6]),
        .O(n22__56_carry_i_9__1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    n22__6
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[8]),
        .Q(n22__6_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__81_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n22__81_carry_n_0,n22__81_carry_n_1,n22__81_carry_n_2,n22__81_carry_n_3,n22__81_carry_n_4,n22__81_carry_n_5,n22__81_carry_n_6,n22__81_carry_n_7}),
        .DI({n22__81_carry_i_1__1_n_0,n22__81_carry_i_2__1_n_0,n22__81_carry_i_3__1_n_0,n22__81_carry_i_4__1_n_0,n22__81_carry_i_5__1_n_0,n22__81_carry_i_6__1_n_0,n22__81_carry_i_7__1_n_0,1'b0}),
        .O({n23[3:0],NLW_n22__81_carry_O_UNCONNECTED[3:0]}),
        .S({n22__81_carry_i_8__1_n_0,n22__81_carry_i_9__1_n_0,n22__81_carry_i_10__1_n_0,n22__81_carry_i_11__1_n_0,n22__81_carry_i_12__1_n_0,n22__81_carry_i_13__1_n_0,n22__81_carry_i_14__1_n_0,n22__81_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__81_carry__0
       (.CI(n22__81_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n22__81_carry__0_CO_UNCONNECTED[7:3],n22__81_carry__0_n_5,n22__81_carry__0_n_6,n22__81_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n22__81_carry__0_i_1__1_n_0,n22__81_carry__0_i_2__1_n_0,n22__81_carry__0_i_3__1_n_0}),
        .O({NLW_n22__81_carry__0_O_UNCONNECTED[7:4],n23[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n22__81_carry__0_i_4__1_n_0,n22__81_carry__0_i_5__1_n_0,n22__81_carry__0_i_6__1_n_0,n22__81_carry__0_i_7__1_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry__0_i_1__1
       (.I0(n22__27_carry__0_n_14),
        .I1(n22__56_carry_n_9),
        .O(n22__81_carry__0_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry__0_i_2__1
       (.I0(n22__27_carry__0_n_15),
        .I1(n22__56_carry_n_10),
        .O(n22__81_carry__0_i_2__1_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry__0_i_3__1
       (.I0(n22__56_carry_n_11),
        .I1(n22__27_carry_n_8),
        .I2(n22__0_carry__0_n_5),
        .O(n22__81_carry__0_i_3__1_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n22__81_carry__0_i_4__1
       (.I0(n22__27_carry__0_n_5),
        .I1(n22__56_carry_n_8),
        .I2(n22__56_carry__0_n_15),
        .O(n22__81_carry__0_i_4__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n22__81_carry__0_i_5__1
       (.I0(n22__27_carry__0_n_14),
        .I1(n22__56_carry_n_9),
        .I2(n22__56_carry_n_8),
        .I3(n22__27_carry__0_n_5),
        .O(n22__81_carry__0_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n22__81_carry__0_i_6__1
       (.I0(n22__27_carry__0_n_15),
        .I1(n22__56_carry_n_10),
        .I2(n22__56_carry_n_9),
        .I3(n22__27_carry__0_n_14),
        .O(n22__81_carry__0_i_6__1_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n22__81_carry__0_i_7__1
       (.I0(n22__0_carry__0_n_5),
        .I1(n22__27_carry_n_8),
        .I2(n22__56_carry_n_11),
        .I3(n22__56_carry_n_10),
        .I4(n22__27_carry__0_n_15),
        .O(n22__81_carry__0_i_7__1_n_0));
  (* HLUTNM = "lutpair22" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_10__1
       (.I0(n22__56_carry_n_13),
        .I1(n22__27_carry_n_10),
        .I2(n22__0_carry__0_n_15),
        .I3(n22__81_carry_i_3__1_n_0),
        .O(n22__81_carry_i_10__1_n_0));
  (* HLUTNM = "lutpair21" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_11__1
       (.I0(n22__56_carry_n_14),
        .I1(n22__27_carry_n_11),
        .I2(n22__0_carry_n_8),
        .I3(n22__81_carry_i_4__1_n_0),
        .O(n22__81_carry_i_11__1_n_0));
  (* HLUTNM = "lutpair20" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_12__1
       (.I0(n22__56_carry_n_15),
        .I1(n22__27_carry_n_12),
        .I2(n22__0_carry_n_9),
        .I3(n22__81_carry_i_5__1_n_0),
        .O(n22__81_carry_i_12__1_n_0));
  (* HLUTNM = "lutpair85" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n22__81_carry_i_13__1
       (.I0(n22__27_carry_n_13),
        .I1(n22__0_carry_n_10),
        .I2(n22__0_carry_n_11),
        .I3(n22__27_carry_n_14),
        .O(n22__81_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n22__81_carry_i_14__1
       (.I0(n22__0_carry_n_12),
        .I1(n22__27_carry_n_15),
        .I2(n22__27_carry_n_14),
        .I3(n22__0_carry_n_11),
        .O(n22__81_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n22__81_carry_i_15__1
       (.I0(n22__0_carry_n_12),
        .I1(n22__27_carry_n_15),
        .O(n22__81_carry_i_15__1_n_0));
  (* HLUTNM = "lutpair23" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry_i_1__1
       (.I0(n22__56_carry_n_12),
        .I1(n22__27_carry_n_9),
        .I2(n22__0_carry__0_n_14),
        .O(n22__81_carry_i_1__1_n_0));
  (* HLUTNM = "lutpair22" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry_i_2__1
       (.I0(n22__56_carry_n_13),
        .I1(n22__27_carry_n_10),
        .I2(n22__0_carry__0_n_15),
        .O(n22__81_carry_i_2__1_n_0));
  (* HLUTNM = "lutpair21" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry_i_3__1
       (.I0(n22__56_carry_n_14),
        .I1(n22__27_carry_n_11),
        .I2(n22__0_carry_n_8),
        .O(n22__81_carry_i_3__1_n_0));
  (* HLUTNM = "lutpair20" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry_i_4__1
       (.I0(n22__56_carry_n_15),
        .I1(n22__27_carry_n_12),
        .I2(n22__0_carry_n_9),
        .O(n22__81_carry_i_4__1_n_0));
  (* HLUTNM = "lutpair85" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry_i_5__1
       (.I0(n22__27_carry_n_13),
        .I1(n22__0_carry_n_10),
        .O(n22__81_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry_i_6__1
       (.I0(n22__0_carry_n_11),
        .I1(n22__27_carry_n_14),
        .O(n22__81_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry_i_7__1
       (.I0(n22__0_carry_n_12),
        .I1(n22__27_carry_n_15),
        .O(n22__81_carry_i_7__1_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_8__1
       (.I0(n22__81_carry_i_1__1_n_0),
        .I1(n22__27_carry_n_8),
        .I2(n22__56_carry_n_11),
        .I3(n22__0_carry__0_n_5),
        .O(n22__81_carry_i_8__1_n_0));
  (* HLUTNM = "lutpair23" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_9__1
       (.I0(n22__56_carry_n_12),
        .I1(n22__27_carry_n_9),
        .I2(n22__0_carry__0_n_14),
        .I3(n22__81_carry_i_2__1_n_0),
        .O(n22__81_carry_i_9__1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[0]),
        .Q(n24[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[1]),
        .Q(n24[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[2]),
        .Q(n24[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[3]),
        .Q(n24[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[4]),
        .Q(n24[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[5]),
        .Q(n24[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[6]),
        .Q(n24[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[7]),
        .Q(n24[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__0_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__0_carry_n_0,n25__0_carry_n_1,n25__0_carry_n_2,n25__0_carry_n_3,n25__0_carry_n_4,n25__0_carry_n_5,n25__0_carry_n_6,n25__0_carry_n_7}),
        .DI({n25__0_carry_i_1__1_n_0,n25__0_carry_i_2__1_n_0,n25__0_carry_i_3__1_n_0,n25__0_carry_i_4__1_n_0,n25__0_carry_i_5__1_n_0,n25__0_carry_i_6__1_n_0,n25__0_carry_i_7__1_n_0,1'b0}),
        .O({n25__0_carry_n_8,n25__0_carry_n_9,n25__0_carry_n_10,n25__0_carry_n_11,n25__0_carry_n_12,NLW_n25__0_carry_O_UNCONNECTED[2:0]}),
        .S({n25__0_carry_i_8__1_n_0,n25__0_carry_i_9__1_n_0,n25__0_carry_i_10__1_n_0,n25__0_carry_i_11__1_n_0,n25__0_carry_i_12__1_n_0,n25__0_carry_i_13__1_n_0,n25__0_carry_i_14__1_n_0,n25__0_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__0_carry__0
       (.CI(n25__0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__0_carry__0_CO_UNCONNECTED[7:3],n25__0_carry__0_n_5,NLW_n25__0_carry__0_CO_UNCONNECTED[1],n25__0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25__0_carry__0_i_1__1_n_0,n25__0_carry__0_i_2__1_n_0}),
        .O({NLW_n25__0_carry__0_O_UNCONNECTED[7:2],n25__0_carry__0_n_14,n25__0_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n25__0_carry__0_i_3__1_n_0,n25__0_carry__0_i_4__1_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__0_carry__0_i_1__1
       (.I0(n14__56_carry_0[9]),
        .I1(n4[7]),
        .I2(n14__56_carry_0[10]),
        .I3(n4[6]),
        .O(n25__0_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n25__0_carry__0_i_2__1
       (.I0(n14__56_carry_0[10]),
        .I1(n4[5]),
        .I2(n14__56_carry_0[9]),
        .I3(n4[6]),
        .I4(n14__56_carry_0[8]),
        .I5(n4[7]),
        .O(n25__0_carry__0_i_2__1_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n25__0_carry__0_i_3__1
       (.I0(n4[6]),
        .I1(n14__56_carry_0[9]),
        .I2(n14__56_carry_0[10]),
        .I3(n4[7]),
        .O(n25__0_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n25__0_carry__0_i_4__1
       (.I0(n14__56_carry_0[8]),
        .I1(n4[5]),
        .I2(n4[6]),
        .I3(n14__56_carry_0[10]),
        .I4(n4[7]),
        .I5(n14__56_carry_0[9]),
        .O(n25__0_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__0_carry_i_10__1
       (.I0(n25__0_carry_i_3__1_n_0),
        .I1(n14__56_carry_0[9]),
        .I2(n4[4]),
        .I3(n25__0_carry_i_19__1_n_0),
        .I4(n4[5]),
        .I5(n14__56_carry_0[8]),
        .O(n25__0_carry_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__0_carry_i_11__1
       (.I0(n25__0_carry_i_4__1_n_0),
        .I1(n14__56_carry_0[9]),
        .I2(n4[3]),
        .I3(n25__0_carry_i_20__1_n_0),
        .I4(n4[4]),
        .I5(n14__56_carry_0[8]),
        .O(n25__0_carry_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n25__0_carry_i_12__1
       (.I0(n4[2]),
        .I1(n25__0_carry_i_21__0_n_0),
        .I2(n4[1]),
        .I3(n14__56_carry_0[9]),
        .I4(n4[0]),
        .I5(n14__56_carry_0[10]),
        .O(n25__0_carry_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n25__0_carry_i_13__1
       (.I0(n4[0]),
        .I1(n14__56_carry_0[10]),
        .I2(n4[1]),
        .I3(n14__56_carry_0[9]),
        .I4(n14__56_carry_0[8]),
        .I5(n4[2]),
        .O(n25__0_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__0_carry_i_14__1
       (.I0(n14__56_carry_0[8]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[9]),
        .I3(n4[0]),
        .O(n25__0_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__0_carry_i_15__1
       (.I0(n4[0]),
        .I1(n14__56_carry_0[8]),
        .O(n25__0_carry_i_15__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_17__1
       (.I0(n4[5]),
        .I1(n14__56_carry_0[10]),
        .O(n25__0_carry_i_17__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_18__1
       (.I0(n4[4]),
        .I1(n14__56_carry_0[10]),
        .O(n25__0_carry_i_18__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_19__1
       (.I0(n4[3]),
        .I1(n14__56_carry_0[10]),
        .O(n25__0_carry_i_19__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__0_carry_i_1__1
       (.I0(n14__56_carry_0[10]),
        .I1(n4[4]),
        .I2(n14__56_carry_0[9]),
        .I3(n4[5]),
        .I4(n14__56_carry_0[8]),
        .I5(n4[6]),
        .O(n25__0_carry_i_1__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_20__1
       (.I0(n4[2]),
        .I1(n14__56_carry_0[10]),
        .O(n25__0_carry_i_20__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_21__0
       (.I0(n4[3]),
        .I1(n14__56_carry_0[8]),
        .O(n25__0_carry_i_21__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__0_carry_i_2__1
       (.I0(n14__56_carry_0[10]),
        .I1(n4[3]),
        .I2(n14__56_carry_0[9]),
        .I3(n4[4]),
        .I4(n14__56_carry_0[8]),
        .I5(n4[5]),
        .O(n25__0_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__0_carry_i_3__1
       (.I0(n14__56_carry_0[10]),
        .I1(n4[2]),
        .I2(n14__56_carry_0[9]),
        .I3(n4[3]),
        .I4(n14__56_carry_0[8]),
        .I5(n4[4]),
        .O(n25__0_carry_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__0_carry_i_4__1
       (.I0(n14__56_carry_0[10]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[9]),
        .I3(n4[2]),
        .I4(n14__56_carry_0[8]),
        .I5(n4[3]),
        .O(n25__0_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n25__0_carry_i_5__1
       (.I0(n14__56_carry_0[9]),
        .I1(n4[2]),
        .I2(n14__56_carry_0[10]),
        .I3(n4[1]),
        .I4(n4[3]),
        .I5(n14__56_carry_0[8]),
        .O(n25__0_carry_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__0_carry_i_6__1
       (.I0(n14__56_carry_0[9]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[10]),
        .I3(n4[0]),
        .O(n25__0_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__0_carry_i_7__1
       (.I0(n14__56_carry_0[8]),
        .I1(n4[1]),
        .O(n25__0_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n25__0_carry_i_8__1
       (.I0(n25__0_carry_i_1__1_n_0),
        .I1(n14__56_carry_0[9]),
        .I2(n4[6]),
        .I3(n25__0_carry_i_17__1_n_0),
        .I4(n4[7]),
        .I5(n14__56_carry_0[8]),
        .O(n25__0_carry_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__0_carry_i_9__1
       (.I0(n25__0_carry_i_2__1_n_0),
        .I1(n14__56_carry_0[9]),
        .I2(n4[5]),
        .I3(n25__0_carry_i_18__1_n_0),
        .I4(n4[6]),
        .I5(n14__56_carry_0[8]),
        .O(n25__0_carry_i_9__1_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__27_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__27_carry_n_0,n25__27_carry_n_1,n25__27_carry_n_2,n25__27_carry_n_3,n25__27_carry_n_4,n25__27_carry_n_5,n25__27_carry_n_6,n25__27_carry_n_7}),
        .DI({n25__27_carry_i_1__1_n_0,n25__27_carry_i_2__1_n_0,n25__27_carry_i_3__1_n_0,n25__27_carry_i_4__1_n_0,n25__27_carry_i_5__1_n_0,n25__27_carry_i_6__1_n_0,n25__27_carry_i_7__1_n_0,1'b0}),
        .O({n25__27_carry_n_8,n25__27_carry_n_9,n25__27_carry_n_10,n25__27_carry_n_11,n25__27_carry_n_12,n25__27_carry_n_13,n25__27_carry_n_14,n25__27_carry_n_15}),
        .S({n25__27_carry_i_8__1_n_0,n25__27_carry_i_9__1_n_0,n25__27_carry_i_10__1_n_0,n25__27_carry_i_11__1_n_0,n25__27_carry_i_12__1_n_0,n25__27_carry_i_13__1_n_0,n25__27_carry_i_14__1_n_0,n25__27_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__27_carry__0
       (.CI(n25__27_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__27_carry__0_CO_UNCONNECTED[7:3],n25__27_carry__0_n_5,NLW_n25__27_carry__0_CO_UNCONNECTED[1],n25__27_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25__27_carry__0_i_1__1_n_0,n25__27_carry__0_i_2__1_n_0}),
        .O({NLW_n25__27_carry__0_O_UNCONNECTED[7:2],n25__27_carry__0_n_14,n25__27_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n25__27_carry__0_i_3__1_n_0,n25__27_carry__0_i_4__1_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__27_carry__0_i_1__1
       (.I0(n14__56_carry_0[12]),
        .I1(n4[7]),
        .I2(n14__56_carry_0[13]),
        .I3(n4[6]),
        .O(n25__27_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n25__27_carry__0_i_2__1
       (.I0(n14__56_carry_0[13]),
        .I1(n4[5]),
        .I2(n14__56_carry_0[12]),
        .I3(n4[6]),
        .I4(n14__56_carry_0[11]),
        .I5(n4[7]),
        .O(n25__27_carry__0_i_2__1_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n25__27_carry__0_i_3__1
       (.I0(n4[6]),
        .I1(n14__56_carry_0[12]),
        .I2(n14__56_carry_0[13]),
        .I3(n4[7]),
        .O(n25__27_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n25__27_carry__0_i_4__1
       (.I0(n14__56_carry_0[11]),
        .I1(n4[5]),
        .I2(n4[6]),
        .I3(n14__56_carry_0[13]),
        .I4(n4[7]),
        .I5(n14__56_carry_0[12]),
        .O(n25__27_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__27_carry_i_10__1
       (.I0(n25__27_carry_i_3__1_n_0),
        .I1(n14__56_carry_0[12]),
        .I2(n4[4]),
        .I3(n25__27_carry_i_18__1_n_0),
        .I4(n4[5]),
        .I5(n14__56_carry_0[11]),
        .O(n25__27_carry_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__27_carry_i_11__1
       (.I0(n25__27_carry_i_4__1_n_0),
        .I1(n14__56_carry_0[12]),
        .I2(n4[3]),
        .I3(n25__27_carry_i_19__1_n_0),
        .I4(n4[4]),
        .I5(n14__56_carry_0[11]),
        .O(n25__27_carry_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n25__27_carry_i_12__1
       (.I0(n4[2]),
        .I1(n25__27_carry_i_20__1_n_0),
        .I2(n4[1]),
        .I3(n14__56_carry_0[12]),
        .I4(n4[0]),
        .I5(n14__56_carry_0[13]),
        .O(n25__27_carry_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n25__27_carry_i_13__1
       (.I0(n4[0]),
        .I1(n14__56_carry_0[13]),
        .I2(n4[1]),
        .I3(n14__56_carry_0[12]),
        .I4(n14__56_carry_0[11]),
        .I5(n4[2]),
        .O(n25__27_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__27_carry_i_14__1
       (.I0(n14__56_carry_0[11]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[12]),
        .I3(n4[0]),
        .O(n25__27_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__27_carry_i_15__1
       (.I0(n4[0]),
        .I1(n14__56_carry_0[11]),
        .O(n25__27_carry_i_15__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_16__1
       (.I0(n4[5]),
        .I1(n14__56_carry_0[13]),
        .O(n25__27_carry_i_16__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_17__1
       (.I0(n4[4]),
        .I1(n14__56_carry_0[13]),
        .O(n25__27_carry_i_17__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_18__1
       (.I0(n4[3]),
        .I1(n14__56_carry_0[13]),
        .O(n25__27_carry_i_18__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_19__1
       (.I0(n4[2]),
        .I1(n14__56_carry_0[13]),
        .O(n25__27_carry_i_19__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__27_carry_i_1__1
       (.I0(n14__56_carry_0[13]),
        .I1(n4[4]),
        .I2(n14__56_carry_0[12]),
        .I3(n4[5]),
        .I4(n14__56_carry_0[11]),
        .I5(n4[6]),
        .O(n25__27_carry_i_1__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_20__1
       (.I0(n4[3]),
        .I1(n14__56_carry_0[11]),
        .O(n25__27_carry_i_20__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__27_carry_i_2__1
       (.I0(n14__56_carry_0[13]),
        .I1(n4[3]),
        .I2(n14__56_carry_0[12]),
        .I3(n4[4]),
        .I4(n14__56_carry_0[11]),
        .I5(n4[5]),
        .O(n25__27_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__27_carry_i_3__1
       (.I0(n14__56_carry_0[13]),
        .I1(n4[2]),
        .I2(n14__56_carry_0[12]),
        .I3(n4[3]),
        .I4(n14__56_carry_0[11]),
        .I5(n4[4]),
        .O(n25__27_carry_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__27_carry_i_4__1
       (.I0(n14__56_carry_0[13]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[12]),
        .I3(n4[2]),
        .I4(n14__56_carry_0[11]),
        .I5(n4[3]),
        .O(n25__27_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n25__27_carry_i_5__1
       (.I0(n14__56_carry_0[12]),
        .I1(n4[2]),
        .I2(n14__56_carry_0[13]),
        .I3(n4[1]),
        .I4(n4[3]),
        .I5(n14__56_carry_0[11]),
        .O(n25__27_carry_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__27_carry_i_6__1
       (.I0(n14__56_carry_0[12]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[13]),
        .I3(n4[0]),
        .O(n25__27_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__27_carry_i_7__1
       (.I0(n14__56_carry_0[11]),
        .I1(n4[1]),
        .O(n25__27_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n25__27_carry_i_8__1
       (.I0(n25__27_carry_i_1__1_n_0),
        .I1(n14__56_carry_0[12]),
        .I2(n4[6]),
        .I3(n25__27_carry_i_16__1_n_0),
        .I4(n4[7]),
        .I5(n14__56_carry_0[11]),
        .O(n25__27_carry_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__27_carry_i_9__1
       (.I0(n25__27_carry_i_2__1_n_0),
        .I1(n14__56_carry_0[12]),
        .I2(n4[5]),
        .I3(n25__27_carry_i_17__1_n_0),
        .I4(n4[6]),
        .I5(n14__56_carry_0[11]),
        .O(n25__27_carry_i_9__1_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__56_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__56_carry_n_0,n25__56_carry_n_1,n25__56_carry_n_2,n25__56_carry_n_3,n25__56_carry_n_4,n25__56_carry_n_5,n25__56_carry_n_6,n25__56_carry_n_7}),
        .DI({n25__56_carry_i_1__1_n_0,n25__56_carry_i_2__1_n_0,n25__56_carry_i_3__1_n_0,n25__56_carry_i_4__1_n_0,n25__56_carry_i_5__1_n_0,n25__56_carry_i_6__1_n_0,n25__56_carry_i_7__1_n_0,1'b0}),
        .O({n25__56_carry_n_8,n25__56_carry_n_9,n25__56_carry_n_10,n25__56_carry_n_11,n25__56_carry_n_12,n25__56_carry_n_13,n25__56_carry_n_14,n25__56_carry_n_15}),
        .S({n25__56_carry_i_8__1_n_0,n25__56_carry_i_9__1_n_0,n25__56_carry_i_10__1_n_0,n25__56_carry_i_11__1_n_0,n25__56_carry_i_12__1_n_0,n25__56_carry_i_13__1_n_0,n25__56_carry_i_14__1_n_0,n25__56_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__56_carry__0
       (.CI(n25__56_carry_n_0),
        .CI_TOP(1'b0),
        .CO(NLW_n25__56_carry__0_CO_UNCONNECTED[7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_n25__56_carry__0_O_UNCONNECTED[7:1],n25__56_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25__56_carry__0_i_1__1_n_0}));
  LUT4 #(
    .INIT(16'hE53F)) 
    n25__56_carry__0_i_1__1
       (.I0(n14__56_carry_0[14]),
        .I1(n4[6]),
        .I2(n14__56_carry_0[15]),
        .I3(n4[7]),
        .O(n25__56_carry__0_i_1__1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n25__56_carry_i_10__1
       (.I0(n4[3]),
        .I1(n4[4]),
        .I2(n14__56_carry_0[15]),
        .I3(n4[5]),
        .I4(n14__56_carry_0[14]),
        .O(n25__56_carry_i_10__1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n25__56_carry_i_11__1
       (.I0(n4[2]),
        .I1(n4[3]),
        .I2(n14__56_carry_0[15]),
        .I3(n4[4]),
        .I4(n14__56_carry_0[14]),
        .O(n25__56_carry_i_11__1_n_0));
  LUT5 #(
    .INIT(32'h9F606060)) 
    n25__56_carry_i_12__1
       (.I0(n4[1]),
        .I1(n4[2]),
        .I2(n14__56_carry_0[15]),
        .I3(n4[3]),
        .I4(n14__56_carry_0[14]),
        .O(n25__56_carry_i_12__1_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__56_carry_i_13__1
       (.I0(n14__56_carry_0[15]),
        .I1(n4[1]),
        .I2(n14__56_carry_0[14]),
        .I3(n4[2]),
        .O(n25__56_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h8777)) 
    n25__56_carry_i_14__1
       (.I0(n14__56_carry_0[15]),
        .I1(n4[0]),
        .I2(n14__56_carry_0[14]),
        .I3(n4[1]),
        .O(n25__56_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__56_carry_i_15__1
       (.I0(n4[0]),
        .I1(n14__56_carry_0[14]),
        .O(n25__56_carry_i_15__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__56_carry_i_1__1
       (.I0(n14__56_carry_0[15]),
        .I1(n4[5]),
        .I2(n14__56_carry_0[14]),
        .I3(n4[6]),
        .O(n25__56_carry_i_1__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__56_carry_i_2__1
       (.I0(n14__56_carry_0[15]),
        .I1(n4[4]),
        .I2(n14__56_carry_0[14]),
        .I3(n4[5]),
        .O(n25__56_carry_i_2__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__56_carry_i_3__1
       (.I0(n14__56_carry_0[15]),
        .I1(n4[3]),
        .I2(n14__56_carry_0[14]),
        .I3(n4[4]),
        .O(n25__56_carry_i_3__1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__56_carry_i_4__1
       (.I0(n14__56_carry_0[15]),
        .I1(n4[2]),
        .I2(n14__56_carry_0[14]),
        .I3(n4[3]),
        .O(n25__56_carry_i_4__1_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n25__56_carry_i_5__1
       (.I0(n4[1]),
        .I1(n14__56_carry_0[15]),
        .O(n25__56_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__56_carry_i_6__1
       (.I0(n14__56_carry_0[15]),
        .I1(n4[1]),
        .O(n25__56_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n25__56_carry_i_7__1
       (.I0(n4[0]),
        .I1(n14__56_carry_0[15]),
        .O(n25__56_carry_i_7__1_n_0));
  LUT5 #(
    .INIT(32'h738CC0C0)) 
    n25__56_carry_i_8__1
       (.I0(n4[5]),
        .I1(n4[6]),
        .I2(n14__56_carry_0[15]),
        .I3(n4[7]),
        .I4(n14__56_carry_0[14]),
        .O(n25__56_carry_i_8__1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n25__56_carry_i_9__1
       (.I0(n4[4]),
        .I1(n4[5]),
        .I2(n14__56_carry_0[15]),
        .I3(n4[6]),
        .I4(n14__56_carry_0[14]),
        .O(n25__56_carry_i_9__1_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__81_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__81_carry_n_0,n25__81_carry_n_1,n25__81_carry_n_2,n25__81_carry_n_3,n25__81_carry_n_4,n25__81_carry_n_5,n25__81_carry_n_6,n25__81_carry_n_7}),
        .DI({n25__81_carry_i_1__1_n_0,n25__81_carry_i_2__1_n_0,n25__81_carry_i_3__1_n_0,n25__81_carry_i_4__1_n_0,n25__81_carry_i_5__1_n_0,n25__81_carry_i_6__1_n_0,n25__81_carry_i_7__1_n_0,1'b0}),
        .O({n26[3:0],NLW_n25__81_carry_O_UNCONNECTED[3:0]}),
        .S({n25__81_carry_i_8__1_n_0,n25__81_carry_i_9__1_n_0,n25__81_carry_i_10__1_n_0,n25__81_carry_i_11__1_n_0,n25__81_carry_i_12__1_n_0,n25__81_carry_i_13__1_n_0,n25__81_carry_i_14__1_n_0,n25__81_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__81_carry__0
       (.CI(n25__81_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__81_carry__0_CO_UNCONNECTED[7:3],n25__81_carry__0_n_5,n25__81_carry__0_n_6,n25__81_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n25__81_carry__0_i_1__1_n_0,n25__81_carry__0_i_2__1_n_0,n25__81_carry__0_i_3__1_n_0}),
        .O({NLW_n25__81_carry__0_O_UNCONNECTED[7:4],n26[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n25__81_carry__0_i_4__1_n_0,n25__81_carry__0_i_5__1_n_0,n25__81_carry__0_i_6__1_n_0,n25__81_carry__0_i_7__1_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry__0_i_1__1
       (.I0(n25__27_carry__0_n_14),
        .I1(n25__56_carry_n_9),
        .O(n25__81_carry__0_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry__0_i_2__1
       (.I0(n25__27_carry__0_n_15),
        .I1(n25__56_carry_n_10),
        .O(n25__81_carry__0_i_2__1_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry__0_i_3__1
       (.I0(n25__56_carry_n_11),
        .I1(n25__27_carry_n_8),
        .I2(n25__0_carry__0_n_5),
        .O(n25__81_carry__0_i_3__1_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n25__81_carry__0_i_4__1
       (.I0(n25__27_carry__0_n_5),
        .I1(n25__56_carry_n_8),
        .I2(n25__56_carry__0_n_15),
        .O(n25__81_carry__0_i_4__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__81_carry__0_i_5__1
       (.I0(n25__27_carry__0_n_14),
        .I1(n25__56_carry_n_9),
        .I2(n25__56_carry_n_8),
        .I3(n25__27_carry__0_n_5),
        .O(n25__81_carry__0_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__81_carry__0_i_6__1
       (.I0(n25__27_carry__0_n_15),
        .I1(n25__56_carry_n_10),
        .I2(n25__56_carry_n_9),
        .I3(n25__27_carry__0_n_14),
        .O(n25__81_carry__0_i_6__1_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n25__81_carry__0_i_7__1
       (.I0(n25__0_carry__0_n_5),
        .I1(n25__27_carry_n_8),
        .I2(n25__56_carry_n_11),
        .I3(n25__56_carry_n_10),
        .I4(n25__27_carry__0_n_15),
        .O(n25__81_carry__0_i_7__1_n_0));
  (* HLUTNM = "lutpair18" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_10__1
       (.I0(n25__56_carry_n_13),
        .I1(n25__27_carry_n_10),
        .I2(n25__0_carry__0_n_15),
        .I3(n25__81_carry_i_3__1_n_0),
        .O(n25__81_carry_i_10__1_n_0));
  (* HLUTNM = "lutpair17" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_11__1
       (.I0(n25__56_carry_n_14),
        .I1(n25__27_carry_n_11),
        .I2(n25__0_carry_n_8),
        .I3(n25__81_carry_i_4__1_n_0),
        .O(n25__81_carry_i_11__1_n_0));
  (* HLUTNM = "lutpair16" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_12__1
       (.I0(n25__56_carry_n_15),
        .I1(n25__27_carry_n_12),
        .I2(n25__0_carry_n_9),
        .I3(n25__81_carry_i_5__1_n_0),
        .O(n25__81_carry_i_12__1_n_0));
  (* HLUTNM = "lutpair84" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n25__81_carry_i_13__1
       (.I0(n25__27_carry_n_13),
        .I1(n25__0_carry_n_10),
        .I2(n25__0_carry_n_11),
        .I3(n25__27_carry_n_14),
        .O(n25__81_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__81_carry_i_14__1
       (.I0(n25__0_carry_n_12),
        .I1(n25__27_carry_n_15),
        .I2(n25__27_carry_n_14),
        .I3(n25__0_carry_n_11),
        .O(n25__81_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n25__81_carry_i_15__1
       (.I0(n25__0_carry_n_12),
        .I1(n25__27_carry_n_15),
        .O(n25__81_carry_i_15__1_n_0));
  (* HLUTNM = "lutpair19" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry_i_1__1
       (.I0(n25__56_carry_n_12),
        .I1(n25__27_carry_n_9),
        .I2(n25__0_carry__0_n_14),
        .O(n25__81_carry_i_1__1_n_0));
  (* HLUTNM = "lutpair18" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry_i_2__1
       (.I0(n25__56_carry_n_13),
        .I1(n25__27_carry_n_10),
        .I2(n25__0_carry__0_n_15),
        .O(n25__81_carry_i_2__1_n_0));
  (* HLUTNM = "lutpair17" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry_i_3__1
       (.I0(n25__56_carry_n_14),
        .I1(n25__27_carry_n_11),
        .I2(n25__0_carry_n_8),
        .O(n25__81_carry_i_3__1_n_0));
  (* HLUTNM = "lutpair16" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry_i_4__1
       (.I0(n25__56_carry_n_15),
        .I1(n25__27_carry_n_12),
        .I2(n25__0_carry_n_9),
        .O(n25__81_carry_i_4__1_n_0));
  (* HLUTNM = "lutpair84" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry_i_5__1
       (.I0(n25__27_carry_n_13),
        .I1(n25__0_carry_n_10),
        .O(n25__81_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry_i_6__1
       (.I0(n25__0_carry_n_11),
        .I1(n25__27_carry_n_14),
        .O(n25__81_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry_i_7__1
       (.I0(n25__0_carry_n_12),
        .I1(n25__27_carry_n_15),
        .O(n25__81_carry_i_7__1_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_8__1
       (.I0(n25__81_carry_i_1__1_n_0),
        .I1(n25__27_carry_n_8),
        .I2(n25__56_carry_n_11),
        .I3(n25__0_carry__0_n_5),
        .O(n25__81_carry_i_8__1_n_0));
  (* HLUTNM = "lutpair19" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_9__1
       (.I0(n25__56_carry_n_12),
        .I1(n25__27_carry_n_9),
        .I2(n25__0_carry__0_n_14),
        .I3(n25__81_carry_i_2__1_n_0),
        .O(n25__81_carry_i_9__1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[0]),
        .Q(n27[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[1]),
        .Q(n27[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[2]),
        .Q(n27[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[3]),
        .Q(n27[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[4]),
        .Q(n27[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[5]),
        .Q(n27[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[6]),
        .Q(n27[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[7]),
        .Q(n27[7]),
        .R(rst_i));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_2 
       (.I0(n24[7]),
        .I1(n27[7]),
        .O(\n29[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_3 
       (.I0(n24[6]),
        .I1(n27[6]),
        .O(\n29[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_4 
       (.I0(n24[5]),
        .I1(n27[5]),
        .O(\n29[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_5 
       (.I0(n24[4]),
        .I1(n27[4]),
        .O(\n29[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_6 
       (.I0(n24[3]),
        .I1(n27[3]),
        .O(\n29[7]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_7 
       (.I0(n24[2]),
        .I1(n27[2]),
        .O(\n29[7]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_8 
       (.I0(n24[1]),
        .I1(n27[1]),
        .O(\n29[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_9 
       (.I0(n24[0]),
        .I1(n27[0]),
        .O(\n29[7]_i_9_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[0]),
        .Q(n29[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[1]),
        .Q(n29[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[2]),
        .Q(n29[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[3]),
        .Q(n29[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[4]),
        .Q(n29[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[5]),
        .Q(n29[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[6]),
        .Q(n29[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[7]),
        .Q(n29[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n29_reg[7]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\NLW_n29_reg[7]_i_1_CO_UNCONNECTED [7],\n29_reg[7]_i_1_n_1 ,\n29_reg[7]_i_1_n_2 ,\n29_reg[7]_i_1_n_3 ,\n29_reg[7]_i_1_n_4 ,\n29_reg[7]_i_1_n_5 ,\n29_reg[7]_i_1_n_6 ,\n29_reg[7]_i_1_n_7 }),
        .DI({1'b0,n24[6:0]}),
        .O(n28),
        .S({\n29[7]_i_2_n_0 ,\n29[7]_i_3_n_0 ,\n29[7]_i_4_n_0 ,\n29[7]_i_5_n_0 ,\n29[7]_i_6_n_0 ,\n29[7]_i_7_n_0 ,\n29[7]_i_8_n_0 ,\n29[7]_i_9_n_0 }));
  LUT2 #(
    .INIT(4'h6)) 
    \n33[0]_i_1__1 
       (.I0(n29[0]),
        .I1(n10[0]),
        .O(n31[0]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[10]_i_1__1 
       (.I0(n21[2]),
        .I1(\n8_reg_n_0_[2] ),
        .I2(\n8_reg_n_0_[1] ),
        .I3(n21[1]),
        .I4(\n8_reg_n_0_[0] ),
        .I5(n21[0]),
        .O(\n33[10]_i_1__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[11]_i_1__1 
       (.I0(n21[3]),
        .I1(\n8_reg_n_0_[3] ),
        .I2(\n33[12]_i_2__1_n_0 ),
        .O(\n33[11]_i_1__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[12]_i_1__1 
       (.I0(n21[4]),
        .I1(\n8_reg_n_0_[4] ),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[3]),
        .I4(\n33[12]_i_2__1_n_0 ),
        .O(\n33[12]_i_1__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[12]_i_2__1 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n33[12]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[13]_i_1__1 
       (.I0(n21[5]),
        .I1(\n8_reg_n_0_[5] ),
        .I2(\n33[14]_i_2__1_n_0 ),
        .O(\n33[13]_i_1__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[14]_i_1__1 
       (.I0(n21[6]),
        .I1(\n8_reg_n_0_[6] ),
        .I2(\n8_reg_n_0_[5] ),
        .I3(n21[5]),
        .I4(\n33[14]_i_2__1_n_0 ),
        .O(\n33[14]_i_1__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[14]_i_2__1 
       (.I0(\n33[12]_i_2__1_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n33[14]_i_2__1_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[15]_i_1__1 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n33[15]_i_2__1_n_0 ),
        .O(n30[7]));
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[15]_i_2__1 
       (.I0(\n33[14]_i_2__1_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n33[15]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[1]_i_1__1 
       (.I0(n29[1]),
        .I1(n10[1]),
        .I2(n10[0]),
        .I3(n29[0]),
        .O(n31[1]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[2]_i_1__1 
       (.I0(n29[2]),
        .I1(n10[2]),
        .I2(n10[1]),
        .I3(n29[1]),
        .I4(n10[0]),
        .I5(n29[0]),
        .O(\n33[2]_i_1__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[3]_i_1__1 
       (.I0(n29[3]),
        .I1(n10[3]),
        .I2(\n33[4]_i_2__1_n_0 ),
        .O(\n33[3]_i_1__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[4]_i_1__1 
       (.I0(n29[4]),
        .I1(n10[4]),
        .I2(n10[3]),
        .I3(n29[3]),
        .I4(\n33[4]_i_2__1_n_0 ),
        .O(\n33[4]_i_1__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[4]_i_2__1 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n33[4]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[5]_i_1__1 
       (.I0(n29[5]),
        .I1(n10[5]),
        .I2(\n33[6]_i_2__1_n_0 ),
        .O(\n33[5]_i_1__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[6]_i_1__1 
       (.I0(n29[6]),
        .I1(n10[6]),
        .I2(n10[5]),
        .I3(n29[5]),
        .I4(\n33[6]_i_2__1_n_0 ),
        .O(\n33[6]_i_1__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[6]_i_2__1 
       (.I0(\n33[4]_i_2__1_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n33[6]_i_2__1_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[7]_i_1__1 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n33[7]_i_2__1_n_0 ),
        .O(n31[7]));
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[7]_i_2__1 
       (.I0(\n33[6]_i_2__1_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n33[7]_i_2__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n33[8]_i_1__0 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .O(n30[0]));
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[9]_i_1__1 
       (.I0(n21[1]),
        .I1(\n8_reg_n_0_[1] ),
        .I2(\n8_reg_n_0_[0] ),
        .I3(n21[0]),
        .O(\n33[9]_i_1__1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[0]),
        .Q(i1[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[10]_i_1__1_n_0 ),
        .Q(i1[24]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[11]_i_1__1_n_0 ),
        .Q(i1[25]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[12]_i_1__1_n_0 ),
        .Q(i1[26]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[13]_i_1__1_n_0 ),
        .Q(i1[27]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[14]_i_1__1_n_0 ),
        .Q(i1[28]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n30[7]),
        .Q(i1[29]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[1]),
        .Q(i1[15]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[2]_i_1__1_n_0 ),
        .Q(i1[16]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[3]_i_1__1_n_0 ),
        .Q(i1[17]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[4]_i_1__1_n_0 ),
        .Q(i1[18]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[5]_i_1__1_n_0 ),
        .Q(i1[19]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[6]_i_1__1_n_0 ),
        .Q(i1[20]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[7]),
        .Q(i1[21]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n30[0]),
        .Q(i1[22]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[9]_i_1__1_n_0 ),
        .Q(i1[23]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[10]_i_1__1 
       (.I0(\n8_reg_n_0_[1] ),
        .I1(n21[1]),
        .I2(n21[0]),
        .I3(\n8_reg_n_0_[0] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(n341_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[11]_i_1__1 
       (.I0(\n37[12]_i_2__1_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .O(n341_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[12]_i_1__1 
       (.I0(\n8_reg_n_0_[3] ),
        .I1(n21[3]),
        .I2(\n37[12]_i_2__1_n_0 ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(n341_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[12]_i_2__1 
       (.I0(\n8_reg_n_0_[0] ),
        .I1(n21[0]),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n37[12]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[13]_i_1__1 
       (.I0(\n37[14]_i_2__1_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(n341_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[14]_i_1__1 
       (.I0(\n8_reg_n_0_[5] ),
        .I1(n21[5]),
        .I2(\n37[14]_i_2__1_n_0 ),
        .I3(n21[6]),
        .I4(\n8_reg_n_0_[6] ),
        .O(n341_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[14]_i_2__1 
       (.I0(\n37[12]_i_2__1_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n37[14]_i_2__1_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[15]_i_1__1 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n37[15]_i_2__1_n_0 ),
        .O(n341_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[15]_i_2__1 
       (.I0(\n37[14]_i_2__1_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n37[15]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[1]_i_1__1 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .O(n350_out[1]));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[2]_i_1__1 
       (.I0(n10[1]),
        .I1(n29[1]),
        .I2(n29[0]),
        .I3(n10[0]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(n350_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[3]_i_1__1 
       (.I0(\n37[4]_i_2__1_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .O(n350_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[4]_i_1__1 
       (.I0(n10[3]),
        .I1(n29[3]),
        .I2(\n37[4]_i_2__1_n_0 ),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(n350_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[4]_i_2__1 
       (.I0(n10[0]),
        .I1(n29[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n37[4]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[5]_i_1__1 
       (.I0(\n37[6]_i_2__1_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(n350_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[6]_i_1__1 
       (.I0(n10[5]),
        .I1(n29[5]),
        .I2(\n37[6]_i_2__1_n_0 ),
        .I3(n29[6]),
        .I4(n10[6]),
        .O(n350_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[6]_i_2__1 
       (.I0(\n37[4]_i_2__1_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n37[6]_i_2__1_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[7]_i_1__1 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n37[7]_i_2__1_n_0 ),
        .O(n350_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[7]_i_2__1 
       (.I0(\n37[6]_i_2__1_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n37[7]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[9]_i_1__1 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .O(n341_out[1]));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[2]),
        .Q(i1[9]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[3]),
        .Q(i1[10]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[4]),
        .Q(i1[11]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[5]),
        .Q(i1[12]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[6]),
        .Q(i1[13]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[7]),
        .Q(i1[14]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[1]),
        .Q(i1[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[2]),
        .Q(i1[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[3]),
        .Q(i1[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[4]),
        .Q(i1[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[5]),
        .Q(i1[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[6]),
        .Q(i1[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[7]),
        .Q(i1[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[1]),
        .Q(i1[8]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[0]),
        .Q(n4[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[1]),
        .Q(n4[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[2]),
        .Q(n4[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[3]),
        .Q(n4[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[4]),
        .Q(n4[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[5]),
        .Q(n4[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[6]),
        .Q(n4[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s4_3[7]),
        .Q(n4[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[0]),
        .Q(\n7_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[1]),
        .Q(\n7_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[2]),
        .Q(\n7_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[3]),
        .Q(\n7_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[4]),
        .Q(\n7_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[5]),
        .Q(\n7_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[6]),
        .Q(\n7_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[7]),
        .Q(\n7_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[0] ),
        .Q(\n8_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[1] ),
        .Q(\n8_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[2] ),
        .Q(\n8_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[3] ),
        .Q(\n8_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[4] ),
        .Q(\n8_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[5] ),
        .Q(\n8_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[6] ),
        .Q(\n8_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[7] ),
        .Q(\n8_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[0] ),
        .Q(\n9_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[1] ),
        .Q(\n9_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[2] ),
        .Q(\n9_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[3] ),
        .Q(\n9_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[4] ),
        .Q(\n9_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[5] ),
        .Q(\n9_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[6] ),
        .Q(\n9_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[7] ),
        .Q(\n9_reg_n_0_[7] ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_17" *) 
module switch_elements_cf_fft_512_8_17
   (\n9_reg[0] ,
    s2_3,
    rst_i,
    enable_i,
    clk_i,
    DOUTADOUT,
    s3_3,
    D);
  output [15:0]\n9_reg[0] ;
  output [15:0]s2_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]DOUTADOUT;
  input [15:0]s3_3;
  input [15:0]D;

  wire [15:0]D;
  wire [15:0]DOUTADOUT;
  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire [15:0]n33;
  wire [15:1]n37;
  wire n4;
  wire [15:0]\n9_reg[0] ;
  wire rst_i;
  wire s28_n_0;
  wire [15:0]s2_3;
  wire [15:0]s3_3;

  switch_elements_cf_fft_512_8_18 s25
       (.D(D),
        .DOUTADOUT(DOUTADOUT),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:1],n37[15:9],n37[7:1],n33[0]}),
        .rst_i(rst_i),
        .s3_3(s3_3));
  switch_elements_cf_fft_512_8_31_16 s26
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i8(i8),
        .n4(n4),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_27_17 s28
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:1],n37[15:9],n37[7:1],n33[0]}),
        .i8(i8),
        .\n9_reg[0]_0 (s28_n_0),
        .rst_i(rst_i),
        .s2_3(s2_3));
  switch_elements_cf_fft_512_8_26_18 s29
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33,n37[15:9],n37[7:1]}),
        .i8(i8),
        .\n1_reg[0] (s28_n_0),
        .n4(n4),
        .\n9_reg[0] (\n9_reg[0] ),
        .rst_i(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_18" *) 
module switch_elements_cf_fft_512_8_18
   (i1,
    rst_i,
    enable_i,
    clk_i,
    DOUTADOUT,
    s3_3,
    D);
  output [29:0]i1;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]DOUTADOUT;
  input [15:0]s3_3;
  input [15:0]D;

  wire [15:0]D;
  wire [15:0]DOUTADOUT;
  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [7:0]n10;
  wire n14__0_carry__0_i_1__0_n_0;
  wire n14__0_carry__0_i_2__0_n_0;
  wire n14__0_carry__0_i_3__0_n_0;
  wire n14__0_carry__0_i_4__0_n_0;
  wire n14__0_carry__0_n_14;
  wire n14__0_carry__0_n_15;
  wire n14__0_carry__0_n_5;
  wire n14__0_carry__0_n_7;
  wire n14__0_carry_i_10__0_n_0;
  wire n14__0_carry_i_11__0_n_0;
  wire n14__0_carry_i_12__0_n_0;
  wire n14__0_carry_i_13__0_n_0;
  wire n14__0_carry_i_14__0_n_0;
  wire n14__0_carry_i_15__0_n_0;
  wire n14__0_carry_i_16__0_n_0;
  wire n14__0_carry_i_17__0_n_0;
  wire n14__0_carry_i_18__0_n_0;
  wire n14__0_carry_i_19__0_n_0;
  wire n14__0_carry_i_1__0_n_0;
  wire n14__0_carry_i_20__0_n_0;
  wire n14__0_carry_i_2__0_n_0;
  wire n14__0_carry_i_3__0_n_0;
  wire n14__0_carry_i_4__0_n_0;
  wire n14__0_carry_i_5__0_n_0;
  wire n14__0_carry_i_6__0_n_0;
  wire n14__0_carry_i_7__0_n_0;
  wire n14__0_carry_i_8__0_n_0;
  wire n14__0_carry_i_9__0_n_0;
  wire n14__0_carry_n_0;
  wire n14__0_carry_n_1;
  wire n14__0_carry_n_10;
  wire n14__0_carry_n_11;
  wire n14__0_carry_n_12;
  wire n14__0_carry_n_2;
  wire n14__0_carry_n_3;
  wire n14__0_carry_n_4;
  wire n14__0_carry_n_5;
  wire n14__0_carry_n_6;
  wire n14__0_carry_n_7;
  wire n14__0_carry_n_8;
  wire n14__0_carry_n_9;
  wire n14__27_carry__0_i_1__0_n_0;
  wire n14__27_carry__0_i_2__0_n_0;
  wire n14__27_carry__0_i_3__0_n_0;
  wire n14__27_carry__0_i_4__0_n_0;
  wire n14__27_carry__0_n_14;
  wire n14__27_carry__0_n_15;
  wire n14__27_carry__0_n_5;
  wire n14__27_carry__0_n_7;
  wire n14__27_carry_i_10__0_n_0;
  wire n14__27_carry_i_11__0_n_0;
  wire n14__27_carry_i_12__0_n_0;
  wire n14__27_carry_i_13__0_n_0;
  wire n14__27_carry_i_14__0_n_0;
  wire n14__27_carry_i_15__0_n_0;
  wire n14__27_carry_i_16__0_n_0;
  wire n14__27_carry_i_17__0_n_0;
  wire n14__27_carry_i_18__0_n_0;
  wire n14__27_carry_i_19__0_n_0;
  wire n14__27_carry_i_1__0_n_0;
  wire n14__27_carry_i_20__0_n_0;
  wire n14__27_carry_i_2__0_n_0;
  wire n14__27_carry_i_3__0_n_0;
  wire n14__27_carry_i_4__0_n_0;
  wire n14__27_carry_i_5__0_n_0;
  wire n14__27_carry_i_6__0_n_0;
  wire n14__27_carry_i_7__0_n_0;
  wire n14__27_carry_i_8__0_n_0;
  wire n14__27_carry_i_9__0_n_0;
  wire n14__27_carry_n_0;
  wire n14__27_carry_n_1;
  wire n14__27_carry_n_10;
  wire n14__27_carry_n_11;
  wire n14__27_carry_n_12;
  wire n14__27_carry_n_13;
  wire n14__27_carry_n_14;
  wire n14__27_carry_n_15;
  wire n14__27_carry_n_2;
  wire n14__27_carry_n_3;
  wire n14__27_carry_n_4;
  wire n14__27_carry_n_5;
  wire n14__27_carry_n_6;
  wire n14__27_carry_n_7;
  wire n14__27_carry_n_8;
  wire n14__27_carry_n_9;
  wire n14__56_carry__0_i_1__0_n_0;
  wire n14__56_carry__0_n_15;
  wire n14__56_carry_i_10__0_n_0;
  wire n14__56_carry_i_11__0_n_0;
  wire n14__56_carry_i_12__0_n_0;
  wire n14__56_carry_i_13__0_n_0;
  wire n14__56_carry_i_14__0_n_0;
  wire n14__56_carry_i_15__0_n_0;
  wire n14__56_carry_i_1__0_n_0;
  wire n14__56_carry_i_2__0_n_0;
  wire n14__56_carry_i_3__0_n_0;
  wire n14__56_carry_i_4__0_n_0;
  wire n14__56_carry_i_5__0_n_0;
  wire n14__56_carry_i_6__0_n_0;
  wire n14__56_carry_i_7__0_n_0;
  wire n14__56_carry_i_8__0_n_0;
  wire n14__56_carry_i_9__0_n_0;
  wire n14__56_carry_n_0;
  wire n14__56_carry_n_1;
  wire n14__56_carry_n_10;
  wire n14__56_carry_n_11;
  wire n14__56_carry_n_12;
  wire n14__56_carry_n_13;
  wire n14__56_carry_n_14;
  wire n14__56_carry_n_15;
  wire n14__56_carry_n_2;
  wire n14__56_carry_n_3;
  wire n14__56_carry_n_4;
  wire n14__56_carry_n_5;
  wire n14__56_carry_n_6;
  wire n14__56_carry_n_7;
  wire n14__56_carry_n_8;
  wire n14__56_carry_n_9;
  wire n14__81_carry__0_i_1__0_n_0;
  wire n14__81_carry__0_i_2__0_n_0;
  wire n14__81_carry__0_i_3__0_n_0;
  wire n14__81_carry__0_i_4__0_n_0;
  wire n14__81_carry__0_i_5__0_n_0;
  wire n14__81_carry__0_i_6__0_n_0;
  wire n14__81_carry__0_i_7__0_n_0;
  wire n14__81_carry__0_n_5;
  wire n14__81_carry__0_n_6;
  wire n14__81_carry__0_n_7;
  wire n14__81_carry_i_10__0_n_0;
  wire n14__81_carry_i_11__0_n_0;
  wire n14__81_carry_i_12__0_n_0;
  wire n14__81_carry_i_13__0_n_0;
  wire n14__81_carry_i_14__0_n_0;
  wire n14__81_carry_i_15__0_n_0;
  wire n14__81_carry_i_1__0_n_0;
  wire n14__81_carry_i_2__0_n_0;
  wire n14__81_carry_i_3__0_n_0;
  wire n14__81_carry_i_4__0_n_0;
  wire n14__81_carry_i_5__0_n_0;
  wire n14__81_carry_i_6__0_n_0;
  wire n14__81_carry_i_7__0_n_0;
  wire n14__81_carry_i_8__0_n_0;
  wire n14__81_carry_i_9__0_n_0;
  wire n14__81_carry_n_0;
  wire n14__81_carry_n_1;
  wire n14__81_carry_n_2;
  wire n14__81_carry_n_3;
  wire n14__81_carry_n_4;
  wire n14__81_carry_n_5;
  wire n14__81_carry_n_6;
  wire n14__81_carry_n_7;
  wire [7:0]n15;
  wire \n16_reg_n_0_[0] ;
  wire \n16_reg_n_0_[1] ;
  wire \n16_reg_n_0_[2] ;
  wire \n16_reg_n_0_[3] ;
  wire \n16_reg_n_0_[4] ;
  wire \n16_reg_n_0_[5] ;
  wire \n16_reg_n_0_[6] ;
  wire \n16_reg_n_0_[7] ;
  wire [14:7]n17;
  wire n17__0_carry__0_i_1__0_n_0;
  wire n17__0_carry__0_i_2__0_n_0;
  wire n17__0_carry__0_i_3__0_n_0;
  wire n17__0_carry__0_i_4__0_n_0;
  wire n17__0_carry__0_n_14;
  wire n17__0_carry__0_n_15;
  wire n17__0_carry__0_n_5;
  wire n17__0_carry__0_n_7;
  wire n17__0_carry_i_10__0_n_0;
  wire n17__0_carry_i_11__0_n_0;
  wire n17__0_carry_i_12__0_n_0;
  wire n17__0_carry_i_13__0_n_0;
  wire n17__0_carry_i_14__0_n_0;
  wire n17__0_carry_i_15__0_n_0;
  wire n17__0_carry_i_16__0_n_0;
  wire n17__0_carry_i_17__0_n_0;
  wire n17__0_carry_i_18__0_n_0;
  wire n17__0_carry_i_19__0_n_0;
  wire n17__0_carry_i_1__0_n_0;
  wire n17__0_carry_i_20__0_n_0;
  wire n17__0_carry_i_2__0_n_0;
  wire n17__0_carry_i_3__0_n_0;
  wire n17__0_carry_i_4__0_n_0;
  wire n17__0_carry_i_5__0_n_0;
  wire n17__0_carry_i_6__0_n_0;
  wire n17__0_carry_i_7__0_n_0;
  wire n17__0_carry_i_8__0_n_0;
  wire n17__0_carry_i_9__0_n_0;
  wire n17__0_carry_n_0;
  wire n17__0_carry_n_1;
  wire n17__0_carry_n_10;
  wire n17__0_carry_n_11;
  wire n17__0_carry_n_12;
  wire n17__0_carry_n_2;
  wire n17__0_carry_n_3;
  wire n17__0_carry_n_4;
  wire n17__0_carry_n_5;
  wire n17__0_carry_n_6;
  wire n17__0_carry_n_7;
  wire n17__0_carry_n_8;
  wire n17__0_carry_n_9;
  wire n17__27_carry__0_i_1__0_n_0;
  wire n17__27_carry__0_i_2__0_n_0;
  wire n17__27_carry__0_i_3__0_n_0;
  wire n17__27_carry__0_i_4__0_n_0;
  wire n17__27_carry__0_n_14;
  wire n17__27_carry__0_n_15;
  wire n17__27_carry__0_n_5;
  wire n17__27_carry__0_n_7;
  wire n17__27_carry_i_10__0_n_0;
  wire n17__27_carry_i_11__0_n_0;
  wire n17__27_carry_i_12__0_n_0;
  wire n17__27_carry_i_13__0_n_0;
  wire n17__27_carry_i_14__0_n_0;
  wire n17__27_carry_i_15__0_n_0;
  wire n17__27_carry_i_16__0_n_0;
  wire n17__27_carry_i_17__0_n_0;
  wire n17__27_carry_i_18__0_n_0;
  wire n17__27_carry_i_19__0_n_0;
  wire n17__27_carry_i_1__0_n_0;
  wire n17__27_carry_i_20__0_n_0;
  wire n17__27_carry_i_2__0_n_0;
  wire n17__27_carry_i_3__0_n_0;
  wire n17__27_carry_i_4__0_n_0;
  wire n17__27_carry_i_5__0_n_0;
  wire n17__27_carry_i_6__0_n_0;
  wire n17__27_carry_i_7__0_n_0;
  wire n17__27_carry_i_8__0_n_0;
  wire n17__27_carry_i_9__0_n_0;
  wire n17__27_carry_n_0;
  wire n17__27_carry_n_1;
  wire n17__27_carry_n_10;
  wire n17__27_carry_n_11;
  wire n17__27_carry_n_12;
  wire n17__27_carry_n_13;
  wire n17__27_carry_n_14;
  wire n17__27_carry_n_15;
  wire n17__27_carry_n_2;
  wire n17__27_carry_n_3;
  wire n17__27_carry_n_4;
  wire n17__27_carry_n_5;
  wire n17__27_carry_n_6;
  wire n17__27_carry_n_7;
  wire n17__27_carry_n_8;
  wire n17__27_carry_n_9;
  wire n17__56_carry__0_i_1__0_n_0;
  wire n17__56_carry__0_n_15;
  wire n17__56_carry_i_10__0_n_0;
  wire n17__56_carry_i_11__0_n_0;
  wire n17__56_carry_i_12__0_n_0;
  wire n17__56_carry_i_13__0_n_0;
  wire n17__56_carry_i_14__0_n_0;
  wire n17__56_carry_i_15__0_n_0;
  wire n17__56_carry_i_1__0_n_0;
  wire n17__56_carry_i_2__0_n_0;
  wire n17__56_carry_i_3__0_n_0;
  wire n17__56_carry_i_4__0_n_0;
  wire n17__56_carry_i_5__0_n_0;
  wire n17__56_carry_i_6__0_n_0;
  wire n17__56_carry_i_7__0_n_0;
  wire n17__56_carry_i_8__0_n_0;
  wire n17__56_carry_i_9__0_n_0;
  wire n17__56_carry_n_0;
  wire n17__56_carry_n_1;
  wire n17__56_carry_n_10;
  wire n17__56_carry_n_11;
  wire n17__56_carry_n_12;
  wire n17__56_carry_n_13;
  wire n17__56_carry_n_14;
  wire n17__56_carry_n_15;
  wire n17__56_carry_n_2;
  wire n17__56_carry_n_3;
  wire n17__56_carry_n_4;
  wire n17__56_carry_n_5;
  wire n17__56_carry_n_6;
  wire n17__56_carry_n_7;
  wire n17__56_carry_n_8;
  wire n17__56_carry_n_9;
  wire n17__81_carry__0_i_1__0_n_0;
  wire n17__81_carry__0_i_2__0_n_0;
  wire n17__81_carry__0_i_3__0_n_0;
  wire n17__81_carry__0_i_4__0_n_0;
  wire n17__81_carry__0_i_5__0_n_0;
  wire n17__81_carry__0_i_6__0_n_0;
  wire n17__81_carry__0_i_7__0_n_0;
  wire n17__81_carry__0_n_5;
  wire n17__81_carry__0_n_6;
  wire n17__81_carry__0_n_7;
  wire n17__81_carry_i_10__0_n_0;
  wire n17__81_carry_i_11__0_n_0;
  wire n17__81_carry_i_12__0_n_0;
  wire n17__81_carry_i_13__0_n_0;
  wire n17__81_carry_i_14__0_n_0;
  wire n17__81_carry_i_15__0_n_0;
  wire n17__81_carry_i_1__0_n_0;
  wire n17__81_carry_i_2__0_n_0;
  wire n17__81_carry_i_3__0_n_0;
  wire n17__81_carry_i_4__0_n_0;
  wire n17__81_carry_i_5__0_n_0;
  wire n17__81_carry_i_6__0_n_0;
  wire n17__81_carry_i_7__0_n_0;
  wire n17__81_carry_i_8__0_n_0;
  wire n17__81_carry_i_9__0_n_0;
  wire n17__81_carry_n_0;
  wire n17__81_carry_n_1;
  wire n17__81_carry_n_2;
  wire n17__81_carry_n_3;
  wire n17__81_carry_n_4;
  wire n17__81_carry_n_5;
  wire n17__81_carry_n_6;
  wire n17__81_carry_n_7;
  wire n19_reg__0_n_0;
  wire n19_reg__1_n_0;
  wire n19_reg__2_n_0;
  wire n19_reg__3_n_0;
  wire n19_reg__4_n_0;
  wire n19_reg__5_n_0;
  wire n19_reg__6_n_0;
  wire n19_reg_n_0;
  wire \n1_reg_n_0_[0] ;
  wire \n1_reg_n_0_[1] ;
  wire \n1_reg_n_0_[2] ;
  wire \n1_reg_n_0_[3] ;
  wire \n1_reg_n_0_[4] ;
  wire \n1_reg_n_0_[5] ;
  wire \n1_reg_n_0_[6] ;
  wire \n1_reg_n_0_[7] ;
  wire [7:0]n2;
  wire [7:0]n202_out;
  wire n20_carry_i_1__1_n_0;
  wire n20_carry_i_2__1_n_0;
  wire n20_carry_i_3__1_n_0;
  wire n20_carry_i_4__1_n_0;
  wire n20_carry_i_5__1_n_0;
  wire n20_carry_i_6__1_n_0;
  wire n20_carry_i_7__1_n_0;
  wire n20_carry_i_8__1_n_0;
  wire n20_carry_n_1;
  wire n20_carry_n_2;
  wire n20_carry_n_3;
  wire n20_carry_n_4;
  wire n20_carry_n_5;
  wire n20_carry_n_6;
  wire n20_carry_n_7;
  wire [7:0]n21;
  wire n22__0_carry__0_i_1__0_n_0;
  wire n22__0_carry__0_i_2__0_n_0;
  wire n22__0_carry__0_i_3__0_n_0;
  wire n22__0_carry__0_i_4__0_n_0;
  wire n22__0_carry__0_n_14;
  wire n22__0_carry__0_n_15;
  wire n22__0_carry__0_n_5;
  wire n22__0_carry__0_n_7;
  wire n22__0_carry_i_10__0_n_0;
  wire n22__0_carry_i_11__0_n_0;
  wire n22__0_carry_i_12__0_n_0;
  wire n22__0_carry_i_13__0_n_0;
  wire n22__0_carry_i_14__0_n_0;
  wire n22__0_carry_i_15__0_n_0;
  wire n22__0_carry_i_16__0_n_0;
  wire n22__0_carry_i_17__0_n_0;
  wire n22__0_carry_i_18__0_n_0;
  wire n22__0_carry_i_19__0_n_0;
  wire n22__0_carry_i_1__0_n_0;
  wire n22__0_carry_i_20__0_n_0;
  wire n22__0_carry_i_2__0_n_0;
  wire n22__0_carry_i_3__0_n_0;
  wire n22__0_carry_i_4__0_n_0;
  wire n22__0_carry_i_5__0_n_0;
  wire n22__0_carry_i_6__0_n_0;
  wire n22__0_carry_i_7__0_n_0;
  wire n22__0_carry_i_8__0_n_0;
  wire n22__0_carry_i_9__0_n_0;
  wire n22__0_carry_n_0;
  wire n22__0_carry_n_1;
  wire n22__0_carry_n_10;
  wire n22__0_carry_n_11;
  wire n22__0_carry_n_12;
  wire n22__0_carry_n_2;
  wire n22__0_carry_n_3;
  wire n22__0_carry_n_4;
  wire n22__0_carry_n_5;
  wire n22__0_carry_n_6;
  wire n22__0_carry_n_7;
  wire n22__0_carry_n_8;
  wire n22__0_carry_n_9;
  wire n22__0_n_0;
  wire n22__1_n_0;
  wire n22__27_carry__0_i_1__0_n_0;
  wire n22__27_carry__0_i_2__0_n_0;
  wire n22__27_carry__0_i_3__0_n_0;
  wire n22__27_carry__0_i_4__0_n_0;
  wire n22__27_carry__0_n_14;
  wire n22__27_carry__0_n_15;
  wire n22__27_carry__0_n_5;
  wire n22__27_carry__0_n_7;
  wire n22__27_carry_i_10__0_n_0;
  wire n22__27_carry_i_11__0_n_0;
  wire n22__27_carry_i_12__0_n_0;
  wire n22__27_carry_i_13__0_n_0;
  wire n22__27_carry_i_14__0_n_0;
  wire n22__27_carry_i_15__0_n_0;
  wire n22__27_carry_i_16__0_n_0;
  wire n22__27_carry_i_17__0_n_0;
  wire n22__27_carry_i_18__0_n_0;
  wire n22__27_carry_i_19__0_n_0;
  wire n22__27_carry_i_1__0_n_0;
  wire n22__27_carry_i_20__0_n_0;
  wire n22__27_carry_i_2__0_n_0;
  wire n22__27_carry_i_3__0_n_0;
  wire n22__27_carry_i_4__0_n_0;
  wire n22__27_carry_i_5__0_n_0;
  wire n22__27_carry_i_6__0_n_0;
  wire n22__27_carry_i_7__0_n_0;
  wire n22__27_carry_i_8__0_n_0;
  wire n22__27_carry_i_9__0_n_0;
  wire n22__27_carry_n_0;
  wire n22__27_carry_n_1;
  wire n22__27_carry_n_10;
  wire n22__27_carry_n_11;
  wire n22__27_carry_n_12;
  wire n22__27_carry_n_13;
  wire n22__27_carry_n_14;
  wire n22__27_carry_n_15;
  wire n22__27_carry_n_2;
  wire n22__27_carry_n_3;
  wire n22__27_carry_n_4;
  wire n22__27_carry_n_5;
  wire n22__27_carry_n_6;
  wire n22__27_carry_n_7;
  wire n22__27_carry_n_8;
  wire n22__27_carry_n_9;
  wire n22__2_n_0;
  wire n22__3_n_0;
  wire n22__4_n_0;
  wire n22__56_carry__0_i_1__0_n_0;
  wire n22__56_carry__0_n_15;
  wire n22__56_carry_i_10__0_n_0;
  wire n22__56_carry_i_11__0_n_0;
  wire n22__56_carry_i_12__0_n_0;
  wire n22__56_carry_i_13__0_n_0;
  wire n22__56_carry_i_14__0_n_0;
  wire n22__56_carry_i_15__0_n_0;
  wire n22__56_carry_i_1__0_n_0;
  wire n22__56_carry_i_2__0_n_0;
  wire n22__56_carry_i_3__0_n_0;
  wire n22__56_carry_i_4__0_n_0;
  wire n22__56_carry_i_5__0_n_0;
  wire n22__56_carry_i_6__0_n_0;
  wire n22__56_carry_i_7__0_n_0;
  wire n22__56_carry_i_8__0_n_0;
  wire n22__56_carry_i_9__0_n_0;
  wire n22__56_carry_n_0;
  wire n22__56_carry_n_1;
  wire n22__56_carry_n_10;
  wire n22__56_carry_n_11;
  wire n22__56_carry_n_12;
  wire n22__56_carry_n_13;
  wire n22__56_carry_n_14;
  wire n22__56_carry_n_15;
  wire n22__56_carry_n_2;
  wire n22__56_carry_n_3;
  wire n22__56_carry_n_4;
  wire n22__56_carry_n_5;
  wire n22__56_carry_n_6;
  wire n22__56_carry_n_7;
  wire n22__56_carry_n_8;
  wire n22__56_carry_n_9;
  wire n22__5_n_0;
  wire n22__6_n_0;
  wire n22__81_carry__0_i_1__0_n_0;
  wire n22__81_carry__0_i_2__0_n_0;
  wire n22__81_carry__0_i_3__0_n_0;
  wire n22__81_carry__0_i_4__0_n_0;
  wire n22__81_carry__0_i_5__0_n_0;
  wire n22__81_carry__0_i_6__0_n_0;
  wire n22__81_carry__0_i_7__0_n_0;
  wire n22__81_carry__0_n_5;
  wire n22__81_carry__0_n_6;
  wire n22__81_carry__0_n_7;
  wire n22__81_carry_i_10__0_n_0;
  wire n22__81_carry_i_11__0_n_0;
  wire n22__81_carry_i_12__0_n_0;
  wire n22__81_carry_i_13__0_n_0;
  wire n22__81_carry_i_14__0_n_0;
  wire n22__81_carry_i_15__0_n_0;
  wire n22__81_carry_i_1__0_n_0;
  wire n22__81_carry_i_2__0_n_0;
  wire n22__81_carry_i_3__0_n_0;
  wire n22__81_carry_i_4__0_n_0;
  wire n22__81_carry_i_5__0_n_0;
  wire n22__81_carry_i_6__0_n_0;
  wire n22__81_carry_i_7__0_n_0;
  wire n22__81_carry_i_8__0_n_0;
  wire n22__81_carry_i_9__0_n_0;
  wire n22__81_carry_n_0;
  wire n22__81_carry_n_1;
  wire n22__81_carry_n_2;
  wire n22__81_carry_n_3;
  wire n22__81_carry_n_4;
  wire n22__81_carry_n_5;
  wire n22__81_carry_n_6;
  wire n22__81_carry_n_7;
  wire n22_n_0;
  wire [7:0]n23;
  wire [7:0]n24;
  wire n25__0_carry__0_i_1__0_n_0;
  wire n25__0_carry__0_i_2__0_n_0;
  wire n25__0_carry__0_i_3__0_n_0;
  wire n25__0_carry__0_i_4__0_n_0;
  wire n25__0_carry__0_n_14;
  wire n25__0_carry__0_n_15;
  wire n25__0_carry__0_n_5;
  wire n25__0_carry__0_n_7;
  wire n25__0_carry_i_10__0_n_0;
  wire n25__0_carry_i_11__0_n_0;
  wire n25__0_carry_i_12__0_n_0;
  wire n25__0_carry_i_13__0_n_0;
  wire n25__0_carry_i_14__0_n_0;
  wire n25__0_carry_i_15__0_n_0;
  wire n25__0_carry_i_17__0_n_0;
  wire n25__0_carry_i_18__0_n_0;
  wire n25__0_carry_i_19__0_n_0;
  wire n25__0_carry_i_1__0_n_0;
  wire n25__0_carry_i_20__0_n_0;
  wire n25__0_carry_i_21_n_0;
  wire n25__0_carry_i_2__0_n_0;
  wire n25__0_carry_i_3__0_n_0;
  wire n25__0_carry_i_4__0_n_0;
  wire n25__0_carry_i_5__0_n_0;
  wire n25__0_carry_i_6__0_n_0;
  wire n25__0_carry_i_7__0_n_0;
  wire n25__0_carry_i_8__0_n_0;
  wire n25__0_carry_i_9__0_n_0;
  wire n25__0_carry_n_0;
  wire n25__0_carry_n_1;
  wire n25__0_carry_n_10;
  wire n25__0_carry_n_11;
  wire n25__0_carry_n_12;
  wire n25__0_carry_n_2;
  wire n25__0_carry_n_3;
  wire n25__0_carry_n_4;
  wire n25__0_carry_n_5;
  wire n25__0_carry_n_6;
  wire n25__0_carry_n_7;
  wire n25__0_carry_n_8;
  wire n25__0_carry_n_9;
  wire n25__27_carry__0_i_1__0_n_0;
  wire n25__27_carry__0_i_2__0_n_0;
  wire n25__27_carry__0_i_3__0_n_0;
  wire n25__27_carry__0_i_4__0_n_0;
  wire n25__27_carry__0_n_14;
  wire n25__27_carry__0_n_15;
  wire n25__27_carry__0_n_5;
  wire n25__27_carry__0_n_7;
  wire n25__27_carry_i_10__0_n_0;
  wire n25__27_carry_i_11__0_n_0;
  wire n25__27_carry_i_12__0_n_0;
  wire n25__27_carry_i_13__0_n_0;
  wire n25__27_carry_i_14__0_n_0;
  wire n25__27_carry_i_15__0_n_0;
  wire n25__27_carry_i_16__0_n_0;
  wire n25__27_carry_i_17__0_n_0;
  wire n25__27_carry_i_18__0_n_0;
  wire n25__27_carry_i_19__0_n_0;
  wire n25__27_carry_i_1__0_n_0;
  wire n25__27_carry_i_20__0_n_0;
  wire n25__27_carry_i_2__0_n_0;
  wire n25__27_carry_i_3__0_n_0;
  wire n25__27_carry_i_4__0_n_0;
  wire n25__27_carry_i_5__0_n_0;
  wire n25__27_carry_i_6__0_n_0;
  wire n25__27_carry_i_7__0_n_0;
  wire n25__27_carry_i_8__0_n_0;
  wire n25__27_carry_i_9__0_n_0;
  wire n25__27_carry_n_0;
  wire n25__27_carry_n_1;
  wire n25__27_carry_n_10;
  wire n25__27_carry_n_11;
  wire n25__27_carry_n_12;
  wire n25__27_carry_n_13;
  wire n25__27_carry_n_14;
  wire n25__27_carry_n_15;
  wire n25__27_carry_n_2;
  wire n25__27_carry_n_3;
  wire n25__27_carry_n_4;
  wire n25__27_carry_n_5;
  wire n25__27_carry_n_6;
  wire n25__27_carry_n_7;
  wire n25__27_carry_n_8;
  wire n25__27_carry_n_9;
  wire n25__56_carry__0_i_1__0_n_0;
  wire n25__56_carry__0_n_15;
  wire n25__56_carry_i_10__0_n_0;
  wire n25__56_carry_i_11__0_n_0;
  wire n25__56_carry_i_12__0_n_0;
  wire n25__56_carry_i_13__0_n_0;
  wire n25__56_carry_i_14__0_n_0;
  wire n25__56_carry_i_15__0_n_0;
  wire n25__56_carry_i_1__0_n_0;
  wire n25__56_carry_i_2__0_n_0;
  wire n25__56_carry_i_3__0_n_0;
  wire n25__56_carry_i_4__0_n_0;
  wire n25__56_carry_i_5__0_n_0;
  wire n25__56_carry_i_6__0_n_0;
  wire n25__56_carry_i_7__0_n_0;
  wire n25__56_carry_i_8__0_n_0;
  wire n25__56_carry_i_9__0_n_0;
  wire n25__56_carry_n_0;
  wire n25__56_carry_n_1;
  wire n25__56_carry_n_10;
  wire n25__56_carry_n_11;
  wire n25__56_carry_n_12;
  wire n25__56_carry_n_13;
  wire n25__56_carry_n_14;
  wire n25__56_carry_n_15;
  wire n25__56_carry_n_2;
  wire n25__56_carry_n_3;
  wire n25__56_carry_n_4;
  wire n25__56_carry_n_5;
  wire n25__56_carry_n_6;
  wire n25__56_carry_n_7;
  wire n25__56_carry_n_8;
  wire n25__56_carry_n_9;
  wire n25__81_carry__0_i_1__0_n_0;
  wire n25__81_carry__0_i_2__0_n_0;
  wire n25__81_carry__0_i_3__0_n_0;
  wire n25__81_carry__0_i_4__0_n_0;
  wire n25__81_carry__0_i_5__0_n_0;
  wire n25__81_carry__0_i_6__0_n_0;
  wire n25__81_carry__0_i_7__0_n_0;
  wire n25__81_carry__0_n_5;
  wire n25__81_carry__0_n_6;
  wire n25__81_carry__0_n_7;
  wire n25__81_carry_i_10__0_n_0;
  wire n25__81_carry_i_11__0_n_0;
  wire n25__81_carry_i_12__0_n_0;
  wire n25__81_carry_i_13__0_n_0;
  wire n25__81_carry_i_14__0_n_0;
  wire n25__81_carry_i_15__0_n_0;
  wire n25__81_carry_i_1__0_n_0;
  wire n25__81_carry_i_2__0_n_0;
  wire n25__81_carry_i_3__0_n_0;
  wire n25__81_carry_i_4__0_n_0;
  wire n25__81_carry_i_5__0_n_0;
  wire n25__81_carry_i_6__0_n_0;
  wire n25__81_carry_i_7__0_n_0;
  wire n25__81_carry_i_8__0_n_0;
  wire n25__81_carry_i_9__0_n_0;
  wire n25__81_carry_n_0;
  wire n25__81_carry_n_1;
  wire n25__81_carry_n_2;
  wire n25__81_carry_n_3;
  wire n25__81_carry_n_4;
  wire n25__81_carry_n_5;
  wire n25__81_carry_n_6;
  wire n25__81_carry_n_7;
  wire [7:0]n26;
  wire [7:0]n27;
  wire [7:0]n28;
  wire [7:0]n29;
  wire \n29[7]_i_2_n_0 ;
  wire \n29[7]_i_3_n_0 ;
  wire \n29[7]_i_4_n_0 ;
  wire \n29[7]_i_5_n_0 ;
  wire \n29[7]_i_6_n_0 ;
  wire \n29[7]_i_7_n_0 ;
  wire \n29[7]_i_8_n_0 ;
  wire \n29[7]_i_9_n_0 ;
  wire \n29_reg[7]_i_1_n_1 ;
  wire \n29_reg[7]_i_1_n_2 ;
  wire \n29_reg[7]_i_1_n_3 ;
  wire \n29_reg[7]_i_1_n_4 ;
  wire \n29_reg[7]_i_1_n_5 ;
  wire \n29_reg[7]_i_1_n_6 ;
  wire \n29_reg[7]_i_1_n_7 ;
  wire [7:0]n30;
  wire [7:0]n31;
  wire \n33[10]_i_1__0_n_0 ;
  wire \n33[11]_i_1__0_n_0 ;
  wire \n33[12]_i_1__0_n_0 ;
  wire \n33[12]_i_2__0_n_0 ;
  wire \n33[13]_i_1__0_n_0 ;
  wire \n33[14]_i_1__0_n_0 ;
  wire \n33[14]_i_2__0_n_0 ;
  wire \n33[15]_i_2__0_n_0 ;
  wire \n33[2]_i_1__0_n_0 ;
  wire \n33[3]_i_1__0_n_0 ;
  wire \n33[4]_i_1__0_n_0 ;
  wire \n33[4]_i_2__0_n_0 ;
  wire \n33[5]_i_1__0_n_0 ;
  wire \n33[6]_i_1__0_n_0 ;
  wire \n33[6]_i_2__0_n_0 ;
  wire \n33[7]_i_2__0_n_0 ;
  wire \n33[9]_i_1__0_n_0 ;
  wire [7:1]n341_out;
  wire [7:1]n350_out;
  wire \n37[12]_i_2__0_n_0 ;
  wire \n37[14]_i_2__0_n_0 ;
  wire \n37[15]_i_2__0_n_0 ;
  wire \n37[4]_i_2__0_n_0 ;
  wire \n37[6]_i_2__0_n_0 ;
  wire \n37[7]_i_2__0_n_0 ;
  wire [7:0]n4;
  wire \n7_reg_n_0_[0] ;
  wire \n7_reg_n_0_[1] ;
  wire \n7_reg_n_0_[2] ;
  wire \n7_reg_n_0_[3] ;
  wire \n7_reg_n_0_[4] ;
  wire \n7_reg_n_0_[5] ;
  wire \n7_reg_n_0_[6] ;
  wire \n7_reg_n_0_[7] ;
  wire \n8_reg_n_0_[0] ;
  wire \n8_reg_n_0_[1] ;
  wire \n8_reg_n_0_[2] ;
  wire \n8_reg_n_0_[3] ;
  wire \n8_reg_n_0_[4] ;
  wire \n8_reg_n_0_[5] ;
  wire \n8_reg_n_0_[6] ;
  wire \n8_reg_n_0_[7] ;
  wire \n9_reg_n_0_[0] ;
  wire \n9_reg_n_0_[1] ;
  wire \n9_reg_n_0_[2] ;
  wire \n9_reg_n_0_[3] ;
  wire \n9_reg_n_0_[4] ;
  wire \n9_reg_n_0_[5] ;
  wire \n9_reg_n_0_[6] ;
  wire \n9_reg_n_0_[7] ;
  wire rst_i;
  wire [15:0]s3_3;
  wire [2:0]NLW_n14__0_carry_O_UNCONNECTED;
  wire [7:1]NLW_n14__0_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n14__0_carry__0_O_UNCONNECTED;
  wire [7:1]NLW_n14__27_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n14__27_carry__0_O_UNCONNECTED;
  wire [7:0]NLW_n14__56_carry__0_CO_UNCONNECTED;
  wire [7:1]NLW_n14__56_carry__0_O_UNCONNECTED;
  wire [3:0]NLW_n14__81_carry_O_UNCONNECTED;
  wire [7:3]NLW_n14__81_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n14__81_carry__0_O_UNCONNECTED;
  wire [2:0]NLW_n17__0_carry_O_UNCONNECTED;
  wire [7:1]NLW_n17__0_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n17__0_carry__0_O_UNCONNECTED;
  wire [7:1]NLW_n17__27_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n17__27_carry__0_O_UNCONNECTED;
  wire [7:0]NLW_n17__56_carry__0_CO_UNCONNECTED;
  wire [7:1]NLW_n17__56_carry__0_O_UNCONNECTED;
  wire [3:0]NLW_n17__81_carry_O_UNCONNECTED;
  wire [7:3]NLW_n17__81_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n17__81_carry__0_O_UNCONNECTED;
  wire [7:7]NLW_n20_carry_CO_UNCONNECTED;
  wire [2:0]NLW_n22__0_carry_O_UNCONNECTED;
  wire [7:1]NLW_n22__0_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n22__0_carry__0_O_UNCONNECTED;
  wire [7:1]NLW_n22__27_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n22__27_carry__0_O_UNCONNECTED;
  wire [7:0]NLW_n22__56_carry__0_CO_UNCONNECTED;
  wire [7:1]NLW_n22__56_carry__0_O_UNCONNECTED;
  wire [3:0]NLW_n22__81_carry_O_UNCONNECTED;
  wire [7:3]NLW_n22__81_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n22__81_carry__0_O_UNCONNECTED;
  wire [2:0]NLW_n25__0_carry_O_UNCONNECTED;
  wire [7:1]NLW_n25__0_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n25__0_carry__0_O_UNCONNECTED;
  wire [7:1]NLW_n25__27_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n25__27_carry__0_O_UNCONNECTED;
  wire [7:0]NLW_n25__56_carry__0_CO_UNCONNECTED;
  wire [7:1]NLW_n25__56_carry__0_O_UNCONNECTED;
  wire [3:0]NLW_n25__81_carry_O_UNCONNECTED;
  wire [7:3]NLW_n25__81_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n25__81_carry__0_O_UNCONNECTED;
  wire [7:7]\NLW_n29_reg[7]_i_1_CO_UNCONNECTED ;

  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[0] ),
        .Q(n10[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[1] ),
        .Q(n10[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[2] ),
        .Q(n10[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[3] ),
        .Q(n10[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[4] ),
        .Q(n10[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[5] ),
        .Q(n10[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[6] ),
        .Q(n10[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[7] ),
        .Q(n10[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__0_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__0_carry_n_0,n14__0_carry_n_1,n14__0_carry_n_2,n14__0_carry_n_3,n14__0_carry_n_4,n14__0_carry_n_5,n14__0_carry_n_6,n14__0_carry_n_7}),
        .DI({n14__0_carry_i_1__0_n_0,n14__0_carry_i_2__0_n_0,n14__0_carry_i_3__0_n_0,n14__0_carry_i_4__0_n_0,n14__0_carry_i_5__0_n_0,n14__0_carry_i_6__0_n_0,n14__0_carry_i_7__0_n_0,1'b0}),
        .O({n14__0_carry_n_8,n14__0_carry_n_9,n14__0_carry_n_10,n14__0_carry_n_11,n14__0_carry_n_12,NLW_n14__0_carry_O_UNCONNECTED[2:0]}),
        .S({n14__0_carry_i_8__0_n_0,n14__0_carry_i_9__0_n_0,n14__0_carry_i_10__0_n_0,n14__0_carry_i_11__0_n_0,n14__0_carry_i_12__0_n_0,n14__0_carry_i_13__0_n_0,n14__0_carry_i_14__0_n_0,n14__0_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__0_carry__0
       (.CI(n14__0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__0_carry__0_CO_UNCONNECTED[7:3],n14__0_carry__0_n_5,NLW_n14__0_carry__0_CO_UNCONNECTED[1],n14__0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14__0_carry__0_i_1__0_n_0,n14__0_carry__0_i_2__0_n_0}),
        .O({NLW_n14__0_carry__0_O_UNCONNECTED[7:2],n14__0_carry__0_n_14,n14__0_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n14__0_carry__0_i_3__0_n_0,n14__0_carry__0_i_4__0_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__0_carry__0_i_1__0
       (.I0(DOUTADOUT[9]),
        .I1(n22_n_0),
        .I2(DOUTADOUT[10]),
        .I3(n22__0_n_0),
        .O(n14__0_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n14__0_carry__0_i_2__0
       (.I0(DOUTADOUT[10]),
        .I1(n22__1_n_0),
        .I2(DOUTADOUT[9]),
        .I3(n22__0_n_0),
        .I4(DOUTADOUT[8]),
        .I5(n22_n_0),
        .O(n14__0_carry__0_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n14__0_carry__0_i_3__0
       (.I0(n22__0_n_0),
        .I1(DOUTADOUT[9]),
        .I2(DOUTADOUT[10]),
        .I3(n22_n_0),
        .O(n14__0_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n14__0_carry__0_i_4__0
       (.I0(DOUTADOUT[8]),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(DOUTADOUT[10]),
        .I4(n22_n_0),
        .I5(DOUTADOUT[9]),
        .O(n14__0_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__0_carry_i_10__0
       (.I0(n14__0_carry_i_3__0_n_0),
        .I1(DOUTADOUT[9]),
        .I2(n22__2_n_0),
        .I3(n14__0_carry_i_18__0_n_0),
        .I4(n22__1_n_0),
        .I5(DOUTADOUT[8]),
        .O(n14__0_carry_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__0_carry_i_11__0
       (.I0(n14__0_carry_i_4__0_n_0),
        .I1(DOUTADOUT[9]),
        .I2(n22__3_n_0),
        .I3(n14__0_carry_i_19__0_n_0),
        .I4(n22__2_n_0),
        .I5(DOUTADOUT[8]),
        .O(n14__0_carry_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n14__0_carry_i_12__0
       (.I0(n22__4_n_0),
        .I1(n14__0_carry_i_20__0_n_0),
        .I2(n22__5_n_0),
        .I3(DOUTADOUT[9]),
        .I4(n22__6_n_0),
        .I5(DOUTADOUT[10]),
        .O(n14__0_carry_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n14__0_carry_i_13__0
       (.I0(n22__6_n_0),
        .I1(DOUTADOUT[10]),
        .I2(n22__5_n_0),
        .I3(DOUTADOUT[9]),
        .I4(DOUTADOUT[8]),
        .I5(n22__4_n_0),
        .O(n14__0_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__0_carry_i_14__0
       (.I0(DOUTADOUT[8]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[9]),
        .I3(n22__6_n_0),
        .O(n14__0_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__0_carry_i_15__0
       (.I0(n22__6_n_0),
        .I1(DOUTADOUT[8]),
        .O(n14__0_carry_i_15__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_16__0
       (.I0(n22__1_n_0),
        .I1(DOUTADOUT[10]),
        .O(n14__0_carry_i_16__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_17__0
       (.I0(n22__2_n_0),
        .I1(DOUTADOUT[10]),
        .O(n14__0_carry_i_17__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_18__0
       (.I0(n22__3_n_0),
        .I1(DOUTADOUT[10]),
        .O(n14__0_carry_i_18__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_19__0
       (.I0(n22__4_n_0),
        .I1(DOUTADOUT[10]),
        .O(n14__0_carry_i_19__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__0_carry_i_1__0
       (.I0(DOUTADOUT[10]),
        .I1(n22__2_n_0),
        .I2(DOUTADOUT[9]),
        .I3(n22__1_n_0),
        .I4(DOUTADOUT[8]),
        .I5(n22__0_n_0),
        .O(n14__0_carry_i_1__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_20__0
       (.I0(n22__3_n_0),
        .I1(DOUTADOUT[8]),
        .O(n14__0_carry_i_20__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__0_carry_i_2__0
       (.I0(DOUTADOUT[10]),
        .I1(n22__3_n_0),
        .I2(DOUTADOUT[9]),
        .I3(n22__2_n_0),
        .I4(DOUTADOUT[8]),
        .I5(n22__1_n_0),
        .O(n14__0_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__0_carry_i_3__0
       (.I0(DOUTADOUT[10]),
        .I1(n22__4_n_0),
        .I2(DOUTADOUT[9]),
        .I3(n22__3_n_0),
        .I4(DOUTADOUT[8]),
        .I5(n22__2_n_0),
        .O(n14__0_carry_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__0_carry_i_4__0
       (.I0(DOUTADOUT[10]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[9]),
        .I3(n22__4_n_0),
        .I4(DOUTADOUT[8]),
        .I5(n22__3_n_0),
        .O(n14__0_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n14__0_carry_i_5__0
       (.I0(DOUTADOUT[9]),
        .I1(n22__4_n_0),
        .I2(DOUTADOUT[10]),
        .I3(n22__5_n_0),
        .I4(n22__3_n_0),
        .I5(DOUTADOUT[8]),
        .O(n14__0_carry_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__0_carry_i_6__0
       (.I0(DOUTADOUT[9]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[10]),
        .I3(n22__6_n_0),
        .O(n14__0_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__0_carry_i_7__0
       (.I0(DOUTADOUT[8]),
        .I1(n22__5_n_0),
        .O(n14__0_carry_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n14__0_carry_i_8__0
       (.I0(n14__0_carry_i_1__0_n_0),
        .I1(DOUTADOUT[9]),
        .I2(n22__0_n_0),
        .I3(n14__0_carry_i_16__0_n_0),
        .I4(n22_n_0),
        .I5(DOUTADOUT[8]),
        .O(n14__0_carry_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__0_carry_i_9__0
       (.I0(n14__0_carry_i_2__0_n_0),
        .I1(DOUTADOUT[9]),
        .I2(n22__1_n_0),
        .I3(n14__0_carry_i_17__0_n_0),
        .I4(n22__0_n_0),
        .I5(DOUTADOUT[8]),
        .O(n14__0_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__27_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__27_carry_n_0,n14__27_carry_n_1,n14__27_carry_n_2,n14__27_carry_n_3,n14__27_carry_n_4,n14__27_carry_n_5,n14__27_carry_n_6,n14__27_carry_n_7}),
        .DI({n14__27_carry_i_1__0_n_0,n14__27_carry_i_2__0_n_0,n14__27_carry_i_3__0_n_0,n14__27_carry_i_4__0_n_0,n14__27_carry_i_5__0_n_0,n14__27_carry_i_6__0_n_0,n14__27_carry_i_7__0_n_0,1'b0}),
        .O({n14__27_carry_n_8,n14__27_carry_n_9,n14__27_carry_n_10,n14__27_carry_n_11,n14__27_carry_n_12,n14__27_carry_n_13,n14__27_carry_n_14,n14__27_carry_n_15}),
        .S({n14__27_carry_i_8__0_n_0,n14__27_carry_i_9__0_n_0,n14__27_carry_i_10__0_n_0,n14__27_carry_i_11__0_n_0,n14__27_carry_i_12__0_n_0,n14__27_carry_i_13__0_n_0,n14__27_carry_i_14__0_n_0,n14__27_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__27_carry__0
       (.CI(n14__27_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__27_carry__0_CO_UNCONNECTED[7:3],n14__27_carry__0_n_5,NLW_n14__27_carry__0_CO_UNCONNECTED[1],n14__27_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14__27_carry__0_i_1__0_n_0,n14__27_carry__0_i_2__0_n_0}),
        .O({NLW_n14__27_carry__0_O_UNCONNECTED[7:2],n14__27_carry__0_n_14,n14__27_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n14__27_carry__0_i_3__0_n_0,n14__27_carry__0_i_4__0_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__27_carry__0_i_1__0
       (.I0(DOUTADOUT[12]),
        .I1(n22_n_0),
        .I2(DOUTADOUT[13]),
        .I3(n22__0_n_0),
        .O(n14__27_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n14__27_carry__0_i_2__0
       (.I0(DOUTADOUT[13]),
        .I1(n22__1_n_0),
        .I2(DOUTADOUT[12]),
        .I3(n22__0_n_0),
        .I4(DOUTADOUT[11]),
        .I5(n22_n_0),
        .O(n14__27_carry__0_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n14__27_carry__0_i_3__0
       (.I0(n22__0_n_0),
        .I1(DOUTADOUT[12]),
        .I2(DOUTADOUT[13]),
        .I3(n22_n_0),
        .O(n14__27_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n14__27_carry__0_i_4__0
       (.I0(DOUTADOUT[11]),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(DOUTADOUT[13]),
        .I4(n22_n_0),
        .I5(DOUTADOUT[12]),
        .O(n14__27_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__27_carry_i_10__0
       (.I0(n14__27_carry_i_3__0_n_0),
        .I1(DOUTADOUT[12]),
        .I2(n22__2_n_0),
        .I3(n14__27_carry_i_18__0_n_0),
        .I4(n22__1_n_0),
        .I5(DOUTADOUT[11]),
        .O(n14__27_carry_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__27_carry_i_11__0
       (.I0(n14__27_carry_i_4__0_n_0),
        .I1(DOUTADOUT[12]),
        .I2(n22__3_n_0),
        .I3(n14__27_carry_i_19__0_n_0),
        .I4(n22__2_n_0),
        .I5(DOUTADOUT[11]),
        .O(n14__27_carry_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n14__27_carry_i_12__0
       (.I0(n22__4_n_0),
        .I1(n14__27_carry_i_20__0_n_0),
        .I2(n22__5_n_0),
        .I3(DOUTADOUT[12]),
        .I4(n22__6_n_0),
        .I5(DOUTADOUT[13]),
        .O(n14__27_carry_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n14__27_carry_i_13__0
       (.I0(n22__6_n_0),
        .I1(DOUTADOUT[13]),
        .I2(n22__5_n_0),
        .I3(DOUTADOUT[12]),
        .I4(DOUTADOUT[11]),
        .I5(n22__4_n_0),
        .O(n14__27_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__27_carry_i_14__0
       (.I0(DOUTADOUT[11]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[12]),
        .I3(n22__6_n_0),
        .O(n14__27_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__27_carry_i_15__0
       (.I0(n22__6_n_0),
        .I1(DOUTADOUT[11]),
        .O(n14__27_carry_i_15__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_16__0
       (.I0(n22__1_n_0),
        .I1(DOUTADOUT[13]),
        .O(n14__27_carry_i_16__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_17__0
       (.I0(n22__2_n_0),
        .I1(DOUTADOUT[13]),
        .O(n14__27_carry_i_17__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_18__0
       (.I0(n22__3_n_0),
        .I1(DOUTADOUT[13]),
        .O(n14__27_carry_i_18__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_19__0
       (.I0(n22__4_n_0),
        .I1(DOUTADOUT[13]),
        .O(n14__27_carry_i_19__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__27_carry_i_1__0
       (.I0(DOUTADOUT[13]),
        .I1(n22__2_n_0),
        .I2(DOUTADOUT[12]),
        .I3(n22__1_n_0),
        .I4(DOUTADOUT[11]),
        .I5(n22__0_n_0),
        .O(n14__27_carry_i_1__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_20__0
       (.I0(n22__3_n_0),
        .I1(DOUTADOUT[11]),
        .O(n14__27_carry_i_20__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__27_carry_i_2__0
       (.I0(DOUTADOUT[13]),
        .I1(n22__3_n_0),
        .I2(DOUTADOUT[12]),
        .I3(n22__2_n_0),
        .I4(DOUTADOUT[11]),
        .I5(n22__1_n_0),
        .O(n14__27_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__27_carry_i_3__0
       (.I0(DOUTADOUT[13]),
        .I1(n22__4_n_0),
        .I2(DOUTADOUT[12]),
        .I3(n22__3_n_0),
        .I4(DOUTADOUT[11]),
        .I5(n22__2_n_0),
        .O(n14__27_carry_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__27_carry_i_4__0
       (.I0(DOUTADOUT[13]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[12]),
        .I3(n22__4_n_0),
        .I4(DOUTADOUT[11]),
        .I5(n22__3_n_0),
        .O(n14__27_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n14__27_carry_i_5__0
       (.I0(DOUTADOUT[12]),
        .I1(n22__4_n_0),
        .I2(DOUTADOUT[13]),
        .I3(n22__5_n_0),
        .I4(n22__3_n_0),
        .I5(DOUTADOUT[11]),
        .O(n14__27_carry_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__27_carry_i_6__0
       (.I0(DOUTADOUT[12]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[13]),
        .I3(n22__6_n_0),
        .O(n14__27_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__27_carry_i_7__0
       (.I0(DOUTADOUT[11]),
        .I1(n22__5_n_0),
        .O(n14__27_carry_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n14__27_carry_i_8__0
       (.I0(n14__27_carry_i_1__0_n_0),
        .I1(DOUTADOUT[12]),
        .I2(n22__0_n_0),
        .I3(n14__27_carry_i_16__0_n_0),
        .I4(n22_n_0),
        .I5(DOUTADOUT[11]),
        .O(n14__27_carry_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__27_carry_i_9__0
       (.I0(n14__27_carry_i_2__0_n_0),
        .I1(DOUTADOUT[12]),
        .I2(n22__1_n_0),
        .I3(n14__27_carry_i_17__0_n_0),
        .I4(n22__0_n_0),
        .I5(DOUTADOUT[11]),
        .O(n14__27_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__56_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__56_carry_n_0,n14__56_carry_n_1,n14__56_carry_n_2,n14__56_carry_n_3,n14__56_carry_n_4,n14__56_carry_n_5,n14__56_carry_n_6,n14__56_carry_n_7}),
        .DI({n14__56_carry_i_1__0_n_0,n14__56_carry_i_2__0_n_0,n14__56_carry_i_3__0_n_0,n14__56_carry_i_4__0_n_0,n14__56_carry_i_5__0_n_0,n14__56_carry_i_6__0_n_0,n14__56_carry_i_7__0_n_0,1'b0}),
        .O({n14__56_carry_n_8,n14__56_carry_n_9,n14__56_carry_n_10,n14__56_carry_n_11,n14__56_carry_n_12,n14__56_carry_n_13,n14__56_carry_n_14,n14__56_carry_n_15}),
        .S({n14__56_carry_i_8__0_n_0,n14__56_carry_i_9__0_n_0,n14__56_carry_i_10__0_n_0,n14__56_carry_i_11__0_n_0,n14__56_carry_i_12__0_n_0,n14__56_carry_i_13__0_n_0,n14__56_carry_i_14__0_n_0,n14__56_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__56_carry__0
       (.CI(n14__56_carry_n_0),
        .CI_TOP(1'b0),
        .CO(NLW_n14__56_carry__0_CO_UNCONNECTED[7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_n14__56_carry__0_O_UNCONNECTED[7:1],n14__56_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14__56_carry__0_i_1__0_n_0}));
  LUT4 #(
    .INIT(16'hE53F)) 
    n14__56_carry__0_i_1__0
       (.I0(DOUTADOUT[14]),
        .I1(n22__0_n_0),
        .I2(DOUTADOUT[15]),
        .I3(n22_n_0),
        .O(n14__56_carry__0_i_1__0_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n14__56_carry_i_10__0
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(DOUTADOUT[15]),
        .I3(n22__1_n_0),
        .I4(DOUTADOUT[14]),
        .O(n14__56_carry_i_10__0_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n14__56_carry_i_11__0
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(DOUTADOUT[15]),
        .I3(n22__2_n_0),
        .I4(DOUTADOUT[14]),
        .O(n14__56_carry_i_11__0_n_0));
  LUT5 #(
    .INIT(32'h9F606060)) 
    n14__56_carry_i_12__0
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(DOUTADOUT[15]),
        .I3(n22__3_n_0),
        .I4(DOUTADOUT[14]),
        .O(n14__56_carry_i_12__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__56_carry_i_13__0
       (.I0(DOUTADOUT[15]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[14]),
        .I3(n22__4_n_0),
        .O(n14__56_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h8777)) 
    n14__56_carry_i_14__0
       (.I0(DOUTADOUT[15]),
        .I1(n22__6_n_0),
        .I2(DOUTADOUT[14]),
        .I3(n22__5_n_0),
        .O(n14__56_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__56_carry_i_15__0
       (.I0(n22__6_n_0),
        .I1(DOUTADOUT[14]),
        .O(n14__56_carry_i_15__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__56_carry_i_1__0
       (.I0(DOUTADOUT[15]),
        .I1(n22__1_n_0),
        .I2(DOUTADOUT[14]),
        .I3(n22__0_n_0),
        .O(n14__56_carry_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__56_carry_i_2__0
       (.I0(DOUTADOUT[15]),
        .I1(n22__2_n_0),
        .I2(DOUTADOUT[14]),
        .I3(n22__1_n_0),
        .O(n14__56_carry_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__56_carry_i_3__0
       (.I0(DOUTADOUT[15]),
        .I1(n22__3_n_0),
        .I2(DOUTADOUT[14]),
        .I3(n22__2_n_0),
        .O(n14__56_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__56_carry_i_4__0
       (.I0(DOUTADOUT[15]),
        .I1(n22__4_n_0),
        .I2(DOUTADOUT[14]),
        .I3(n22__3_n_0),
        .O(n14__56_carry_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n14__56_carry_i_5__0
       (.I0(n22__5_n_0),
        .I1(DOUTADOUT[15]),
        .O(n14__56_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__56_carry_i_6__0
       (.I0(DOUTADOUT[15]),
        .I1(n22__5_n_0),
        .O(n14__56_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n14__56_carry_i_7__0
       (.I0(n22__6_n_0),
        .I1(DOUTADOUT[15]),
        .O(n14__56_carry_i_7__0_n_0));
  LUT5 #(
    .INIT(32'h738CC0C0)) 
    n14__56_carry_i_8__0
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(DOUTADOUT[15]),
        .I3(n22_n_0),
        .I4(DOUTADOUT[14]),
        .O(n14__56_carry_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n14__56_carry_i_9__0
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(DOUTADOUT[15]),
        .I3(n22__0_n_0),
        .I4(DOUTADOUT[14]),
        .O(n14__56_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__81_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__81_carry_n_0,n14__81_carry_n_1,n14__81_carry_n_2,n14__81_carry_n_3,n14__81_carry_n_4,n14__81_carry_n_5,n14__81_carry_n_6,n14__81_carry_n_7}),
        .DI({n14__81_carry_i_1__0_n_0,n14__81_carry_i_2__0_n_0,n14__81_carry_i_3__0_n_0,n14__81_carry_i_4__0_n_0,n14__81_carry_i_5__0_n_0,n14__81_carry_i_6__0_n_0,n14__81_carry_i_7__0_n_0,1'b0}),
        .O({n15[3:0],NLW_n14__81_carry_O_UNCONNECTED[3:0]}),
        .S({n14__81_carry_i_8__0_n_0,n14__81_carry_i_9__0_n_0,n14__81_carry_i_10__0_n_0,n14__81_carry_i_11__0_n_0,n14__81_carry_i_12__0_n_0,n14__81_carry_i_13__0_n_0,n14__81_carry_i_14__0_n_0,n14__81_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__81_carry__0
       (.CI(n14__81_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__81_carry__0_CO_UNCONNECTED[7:3],n14__81_carry__0_n_5,n14__81_carry__0_n_6,n14__81_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n14__81_carry__0_i_1__0_n_0,n14__81_carry__0_i_2__0_n_0,n14__81_carry__0_i_3__0_n_0}),
        .O({NLW_n14__81_carry__0_O_UNCONNECTED[7:4],n15[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n14__81_carry__0_i_4__0_n_0,n14__81_carry__0_i_5__0_n_0,n14__81_carry__0_i_6__0_n_0,n14__81_carry__0_i_7__0_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry__0_i_1__0
       (.I0(n14__27_carry__0_n_14),
        .I1(n14__56_carry_n_9),
        .O(n14__81_carry__0_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry__0_i_2__0
       (.I0(n14__27_carry__0_n_15),
        .I1(n14__56_carry_n_10),
        .O(n14__81_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry__0_i_3__0
       (.I0(n14__56_carry_n_11),
        .I1(n14__27_carry_n_8),
        .I2(n14__0_carry__0_n_5),
        .O(n14__81_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n14__81_carry__0_i_4__0
       (.I0(n14__27_carry__0_n_5),
        .I1(n14__56_carry_n_8),
        .I2(n14__56_carry__0_n_15),
        .O(n14__81_carry__0_i_4__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__81_carry__0_i_5__0
       (.I0(n14__27_carry__0_n_14),
        .I1(n14__56_carry_n_9),
        .I2(n14__56_carry_n_8),
        .I3(n14__27_carry__0_n_5),
        .O(n14__81_carry__0_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__81_carry__0_i_6__0
       (.I0(n14__27_carry__0_n_15),
        .I1(n14__56_carry_n_10),
        .I2(n14__56_carry_n_9),
        .I3(n14__27_carry__0_n_14),
        .O(n14__81_carry__0_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n14__81_carry__0_i_7__0
       (.I0(n14__0_carry__0_n_5),
        .I1(n14__27_carry_n_8),
        .I2(n14__56_carry_n_11),
        .I3(n14__56_carry_n_10),
        .I4(n14__27_carry__0_n_15),
        .O(n14__81_carry__0_i_7__0_n_0));
  (* HLUTNM = "lutpair14" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_10__0
       (.I0(n14__56_carry_n_13),
        .I1(n14__27_carry_n_10),
        .I2(n14__0_carry__0_n_15),
        .I3(n14__81_carry_i_3__0_n_0),
        .O(n14__81_carry_i_10__0_n_0));
  (* HLUTNM = "lutpair13" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_11__0
       (.I0(n14__56_carry_n_14),
        .I1(n14__27_carry_n_11),
        .I2(n14__0_carry_n_8),
        .I3(n14__81_carry_i_4__0_n_0),
        .O(n14__81_carry_i_11__0_n_0));
  (* HLUTNM = "lutpair12" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_12__0
       (.I0(n14__56_carry_n_15),
        .I1(n14__27_carry_n_12),
        .I2(n14__0_carry_n_9),
        .I3(n14__81_carry_i_5__0_n_0),
        .O(n14__81_carry_i_12__0_n_0));
  (* HLUTNM = "lutpair83" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n14__81_carry_i_13__0
       (.I0(n14__27_carry_n_13),
        .I1(n14__0_carry_n_10),
        .I2(n14__0_carry_n_11),
        .I3(n14__27_carry_n_14),
        .O(n14__81_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__81_carry_i_14__0
       (.I0(n14__0_carry_n_12),
        .I1(n14__27_carry_n_15),
        .I2(n14__27_carry_n_14),
        .I3(n14__0_carry_n_11),
        .O(n14__81_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n14__81_carry_i_15__0
       (.I0(n14__0_carry_n_12),
        .I1(n14__27_carry_n_15),
        .O(n14__81_carry_i_15__0_n_0));
  (* HLUTNM = "lutpair15" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry_i_1__0
       (.I0(n14__56_carry_n_12),
        .I1(n14__27_carry_n_9),
        .I2(n14__0_carry__0_n_14),
        .O(n14__81_carry_i_1__0_n_0));
  (* HLUTNM = "lutpair14" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry_i_2__0
       (.I0(n14__56_carry_n_13),
        .I1(n14__27_carry_n_10),
        .I2(n14__0_carry__0_n_15),
        .O(n14__81_carry_i_2__0_n_0));
  (* HLUTNM = "lutpair13" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry_i_3__0
       (.I0(n14__56_carry_n_14),
        .I1(n14__27_carry_n_11),
        .I2(n14__0_carry_n_8),
        .O(n14__81_carry_i_3__0_n_0));
  (* HLUTNM = "lutpair12" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry_i_4__0
       (.I0(n14__56_carry_n_15),
        .I1(n14__27_carry_n_12),
        .I2(n14__0_carry_n_9),
        .O(n14__81_carry_i_4__0_n_0));
  (* HLUTNM = "lutpair83" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry_i_5__0
       (.I0(n14__27_carry_n_13),
        .I1(n14__0_carry_n_10),
        .O(n14__81_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry_i_6__0
       (.I0(n14__0_carry_n_11),
        .I1(n14__27_carry_n_14),
        .O(n14__81_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry_i_7__0
       (.I0(n14__0_carry_n_12),
        .I1(n14__27_carry_n_15),
        .O(n14__81_carry_i_7__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_8__0
       (.I0(n14__81_carry_i_1__0_n_0),
        .I1(n14__27_carry_n_8),
        .I2(n14__56_carry_n_11),
        .I3(n14__0_carry__0_n_5),
        .O(n14__81_carry_i_8__0_n_0));
  (* HLUTNM = "lutpair15" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_9__0
       (.I0(n14__56_carry_n_12),
        .I1(n14__27_carry_n_9),
        .I2(n14__0_carry__0_n_14),
        .I3(n14__81_carry_i_2__0_n_0),
        .O(n14__81_carry_i_9__0_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[0]),
        .Q(\n16_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[1]),
        .Q(\n16_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[2]),
        .Q(\n16_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[3]),
        .Q(\n16_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[4]),
        .Q(\n16_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[5]),
        .Q(\n16_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[6]),
        .Q(\n16_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[7]),
        .Q(\n16_reg_n_0_[7] ),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__0_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n17__0_carry_n_0,n17__0_carry_n_1,n17__0_carry_n_2,n17__0_carry_n_3,n17__0_carry_n_4,n17__0_carry_n_5,n17__0_carry_n_6,n17__0_carry_n_7}),
        .DI({n17__0_carry_i_1__0_n_0,n17__0_carry_i_2__0_n_0,n17__0_carry_i_3__0_n_0,n17__0_carry_i_4__0_n_0,n17__0_carry_i_5__0_n_0,n17__0_carry_i_6__0_n_0,n17__0_carry_i_7__0_n_0,1'b0}),
        .O({n17__0_carry_n_8,n17__0_carry_n_9,n17__0_carry_n_10,n17__0_carry_n_11,n17__0_carry_n_12,NLW_n17__0_carry_O_UNCONNECTED[2:0]}),
        .S({n17__0_carry_i_8__0_n_0,n17__0_carry_i_9__0_n_0,n17__0_carry_i_10__0_n_0,n17__0_carry_i_11__0_n_0,n17__0_carry_i_12__0_n_0,n17__0_carry_i_13__0_n_0,n17__0_carry_i_14__0_n_0,n17__0_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__0_carry__0
       (.CI(n17__0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n17__0_carry__0_CO_UNCONNECTED[7:3],n17__0_carry__0_n_5,NLW_n17__0_carry__0_CO_UNCONNECTED[1],n17__0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n17__0_carry__0_i_1__0_n_0,n17__0_carry__0_i_2__0_n_0}),
        .O({NLW_n17__0_carry__0_O_UNCONNECTED[7:2],n17__0_carry__0_n_14,n17__0_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n17__0_carry__0_i_3__0_n_0,n17__0_carry__0_i_4__0_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__0_carry__0_i_1__0
       (.I0(DOUTADOUT[1]),
        .I1(n4[7]),
        .I2(DOUTADOUT[2]),
        .I3(n4[6]),
        .O(n17__0_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n17__0_carry__0_i_2__0
       (.I0(DOUTADOUT[2]),
        .I1(n4[5]),
        .I2(DOUTADOUT[1]),
        .I3(n4[6]),
        .I4(DOUTADOUT[0]),
        .I5(n4[7]),
        .O(n17__0_carry__0_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n17__0_carry__0_i_3__0
       (.I0(n4[6]),
        .I1(DOUTADOUT[1]),
        .I2(DOUTADOUT[2]),
        .I3(n4[7]),
        .O(n17__0_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n17__0_carry__0_i_4__0
       (.I0(DOUTADOUT[0]),
        .I1(n4[5]),
        .I2(n4[6]),
        .I3(DOUTADOUT[2]),
        .I4(n4[7]),
        .I5(DOUTADOUT[1]),
        .O(n17__0_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__0_carry_i_10__0
       (.I0(n17__0_carry_i_3__0_n_0),
        .I1(DOUTADOUT[1]),
        .I2(n4[4]),
        .I3(n17__0_carry_i_18__0_n_0),
        .I4(n4[5]),
        .I5(DOUTADOUT[0]),
        .O(n17__0_carry_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__0_carry_i_11__0
       (.I0(n17__0_carry_i_4__0_n_0),
        .I1(DOUTADOUT[1]),
        .I2(n4[3]),
        .I3(n17__0_carry_i_19__0_n_0),
        .I4(n4[4]),
        .I5(DOUTADOUT[0]),
        .O(n17__0_carry_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n17__0_carry_i_12__0
       (.I0(n4[2]),
        .I1(n17__0_carry_i_20__0_n_0),
        .I2(n4[1]),
        .I3(DOUTADOUT[1]),
        .I4(n4[0]),
        .I5(DOUTADOUT[2]),
        .O(n17__0_carry_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n17__0_carry_i_13__0
       (.I0(n4[0]),
        .I1(DOUTADOUT[2]),
        .I2(n4[1]),
        .I3(DOUTADOUT[1]),
        .I4(DOUTADOUT[0]),
        .I5(n4[2]),
        .O(n17__0_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__0_carry_i_14__0
       (.I0(DOUTADOUT[0]),
        .I1(n4[1]),
        .I2(DOUTADOUT[1]),
        .I3(n4[0]),
        .O(n17__0_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__0_carry_i_15__0
       (.I0(n4[0]),
        .I1(DOUTADOUT[0]),
        .O(n17__0_carry_i_15__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_16__0
       (.I0(n4[5]),
        .I1(DOUTADOUT[2]),
        .O(n17__0_carry_i_16__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_17__0
       (.I0(n4[4]),
        .I1(DOUTADOUT[2]),
        .O(n17__0_carry_i_17__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_18__0
       (.I0(n4[3]),
        .I1(DOUTADOUT[2]),
        .O(n17__0_carry_i_18__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_19__0
       (.I0(n4[2]),
        .I1(DOUTADOUT[2]),
        .O(n17__0_carry_i_19__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__0_carry_i_1__0
       (.I0(DOUTADOUT[2]),
        .I1(n4[4]),
        .I2(DOUTADOUT[1]),
        .I3(n4[5]),
        .I4(DOUTADOUT[0]),
        .I5(n4[6]),
        .O(n17__0_carry_i_1__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_20__0
       (.I0(n4[3]),
        .I1(DOUTADOUT[0]),
        .O(n17__0_carry_i_20__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__0_carry_i_2__0
       (.I0(DOUTADOUT[2]),
        .I1(n4[3]),
        .I2(DOUTADOUT[1]),
        .I3(n4[4]),
        .I4(DOUTADOUT[0]),
        .I5(n4[5]),
        .O(n17__0_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__0_carry_i_3__0
       (.I0(DOUTADOUT[2]),
        .I1(n4[2]),
        .I2(DOUTADOUT[1]),
        .I3(n4[3]),
        .I4(DOUTADOUT[0]),
        .I5(n4[4]),
        .O(n17__0_carry_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__0_carry_i_4__0
       (.I0(DOUTADOUT[2]),
        .I1(n4[1]),
        .I2(DOUTADOUT[1]),
        .I3(n4[2]),
        .I4(DOUTADOUT[0]),
        .I5(n4[3]),
        .O(n17__0_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n17__0_carry_i_5__0
       (.I0(DOUTADOUT[1]),
        .I1(n4[2]),
        .I2(DOUTADOUT[2]),
        .I3(n4[1]),
        .I4(n4[3]),
        .I5(DOUTADOUT[0]),
        .O(n17__0_carry_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__0_carry_i_6__0
       (.I0(DOUTADOUT[1]),
        .I1(n4[1]),
        .I2(DOUTADOUT[2]),
        .I3(n4[0]),
        .O(n17__0_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__0_carry_i_7__0
       (.I0(DOUTADOUT[0]),
        .I1(n4[1]),
        .O(n17__0_carry_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n17__0_carry_i_8__0
       (.I0(n17__0_carry_i_1__0_n_0),
        .I1(DOUTADOUT[1]),
        .I2(n4[6]),
        .I3(n17__0_carry_i_16__0_n_0),
        .I4(n4[7]),
        .I5(DOUTADOUT[0]),
        .O(n17__0_carry_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__0_carry_i_9__0
       (.I0(n17__0_carry_i_2__0_n_0),
        .I1(DOUTADOUT[1]),
        .I2(n4[5]),
        .I3(n17__0_carry_i_17__0_n_0),
        .I4(n4[6]),
        .I5(DOUTADOUT[0]),
        .O(n17__0_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__27_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n17__27_carry_n_0,n17__27_carry_n_1,n17__27_carry_n_2,n17__27_carry_n_3,n17__27_carry_n_4,n17__27_carry_n_5,n17__27_carry_n_6,n17__27_carry_n_7}),
        .DI({n17__27_carry_i_1__0_n_0,n17__27_carry_i_2__0_n_0,n17__27_carry_i_3__0_n_0,n17__27_carry_i_4__0_n_0,n17__27_carry_i_5__0_n_0,n17__27_carry_i_6__0_n_0,n17__27_carry_i_7__0_n_0,1'b0}),
        .O({n17__27_carry_n_8,n17__27_carry_n_9,n17__27_carry_n_10,n17__27_carry_n_11,n17__27_carry_n_12,n17__27_carry_n_13,n17__27_carry_n_14,n17__27_carry_n_15}),
        .S({n17__27_carry_i_8__0_n_0,n17__27_carry_i_9__0_n_0,n17__27_carry_i_10__0_n_0,n17__27_carry_i_11__0_n_0,n17__27_carry_i_12__0_n_0,n17__27_carry_i_13__0_n_0,n17__27_carry_i_14__0_n_0,n17__27_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__27_carry__0
       (.CI(n17__27_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n17__27_carry__0_CO_UNCONNECTED[7:3],n17__27_carry__0_n_5,NLW_n17__27_carry__0_CO_UNCONNECTED[1],n17__27_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n17__27_carry__0_i_1__0_n_0,n17__27_carry__0_i_2__0_n_0}),
        .O({NLW_n17__27_carry__0_O_UNCONNECTED[7:2],n17__27_carry__0_n_14,n17__27_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n17__27_carry__0_i_3__0_n_0,n17__27_carry__0_i_4__0_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__27_carry__0_i_1__0
       (.I0(DOUTADOUT[4]),
        .I1(n4[7]),
        .I2(DOUTADOUT[5]),
        .I3(n4[6]),
        .O(n17__27_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n17__27_carry__0_i_2__0
       (.I0(DOUTADOUT[5]),
        .I1(n4[5]),
        .I2(DOUTADOUT[4]),
        .I3(n4[6]),
        .I4(DOUTADOUT[3]),
        .I5(n4[7]),
        .O(n17__27_carry__0_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n17__27_carry__0_i_3__0
       (.I0(n4[6]),
        .I1(DOUTADOUT[4]),
        .I2(DOUTADOUT[5]),
        .I3(n4[7]),
        .O(n17__27_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n17__27_carry__0_i_4__0
       (.I0(DOUTADOUT[3]),
        .I1(n4[5]),
        .I2(n4[6]),
        .I3(DOUTADOUT[5]),
        .I4(n4[7]),
        .I5(DOUTADOUT[4]),
        .O(n17__27_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__27_carry_i_10__0
       (.I0(n17__27_carry_i_3__0_n_0),
        .I1(DOUTADOUT[4]),
        .I2(n4[4]),
        .I3(n17__27_carry_i_18__0_n_0),
        .I4(n4[5]),
        .I5(DOUTADOUT[3]),
        .O(n17__27_carry_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__27_carry_i_11__0
       (.I0(n17__27_carry_i_4__0_n_0),
        .I1(DOUTADOUT[4]),
        .I2(n4[3]),
        .I3(n17__27_carry_i_19__0_n_0),
        .I4(n4[4]),
        .I5(DOUTADOUT[3]),
        .O(n17__27_carry_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n17__27_carry_i_12__0
       (.I0(n4[2]),
        .I1(n17__27_carry_i_20__0_n_0),
        .I2(n4[1]),
        .I3(DOUTADOUT[4]),
        .I4(n4[0]),
        .I5(DOUTADOUT[5]),
        .O(n17__27_carry_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n17__27_carry_i_13__0
       (.I0(n4[0]),
        .I1(DOUTADOUT[5]),
        .I2(n4[1]),
        .I3(DOUTADOUT[4]),
        .I4(DOUTADOUT[3]),
        .I5(n4[2]),
        .O(n17__27_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__27_carry_i_14__0
       (.I0(DOUTADOUT[3]),
        .I1(n4[1]),
        .I2(DOUTADOUT[4]),
        .I3(n4[0]),
        .O(n17__27_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__27_carry_i_15__0
       (.I0(n4[0]),
        .I1(DOUTADOUT[3]),
        .O(n17__27_carry_i_15__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_16__0
       (.I0(n4[5]),
        .I1(DOUTADOUT[5]),
        .O(n17__27_carry_i_16__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_17__0
       (.I0(n4[4]),
        .I1(DOUTADOUT[5]),
        .O(n17__27_carry_i_17__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_18__0
       (.I0(n4[3]),
        .I1(DOUTADOUT[5]),
        .O(n17__27_carry_i_18__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_19__0
       (.I0(n4[2]),
        .I1(DOUTADOUT[5]),
        .O(n17__27_carry_i_19__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__27_carry_i_1__0
       (.I0(DOUTADOUT[5]),
        .I1(n4[4]),
        .I2(DOUTADOUT[4]),
        .I3(n4[5]),
        .I4(DOUTADOUT[3]),
        .I5(n4[6]),
        .O(n17__27_carry_i_1__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_20__0
       (.I0(n4[3]),
        .I1(DOUTADOUT[3]),
        .O(n17__27_carry_i_20__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__27_carry_i_2__0
       (.I0(DOUTADOUT[5]),
        .I1(n4[3]),
        .I2(DOUTADOUT[4]),
        .I3(n4[4]),
        .I4(DOUTADOUT[3]),
        .I5(n4[5]),
        .O(n17__27_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__27_carry_i_3__0
       (.I0(DOUTADOUT[5]),
        .I1(n4[2]),
        .I2(DOUTADOUT[4]),
        .I3(n4[3]),
        .I4(DOUTADOUT[3]),
        .I5(n4[4]),
        .O(n17__27_carry_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__27_carry_i_4__0
       (.I0(DOUTADOUT[5]),
        .I1(n4[1]),
        .I2(DOUTADOUT[4]),
        .I3(n4[2]),
        .I4(DOUTADOUT[3]),
        .I5(n4[3]),
        .O(n17__27_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n17__27_carry_i_5__0
       (.I0(DOUTADOUT[4]),
        .I1(n4[2]),
        .I2(DOUTADOUT[5]),
        .I3(n4[1]),
        .I4(n4[3]),
        .I5(DOUTADOUT[3]),
        .O(n17__27_carry_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__27_carry_i_6__0
       (.I0(DOUTADOUT[4]),
        .I1(n4[1]),
        .I2(DOUTADOUT[5]),
        .I3(n4[0]),
        .O(n17__27_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__27_carry_i_7__0
       (.I0(DOUTADOUT[3]),
        .I1(n4[1]),
        .O(n17__27_carry_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n17__27_carry_i_8__0
       (.I0(n17__27_carry_i_1__0_n_0),
        .I1(DOUTADOUT[4]),
        .I2(n4[6]),
        .I3(n17__27_carry_i_16__0_n_0),
        .I4(n4[7]),
        .I5(DOUTADOUT[3]),
        .O(n17__27_carry_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__27_carry_i_9__0
       (.I0(n17__27_carry_i_2__0_n_0),
        .I1(DOUTADOUT[4]),
        .I2(n4[5]),
        .I3(n17__27_carry_i_17__0_n_0),
        .I4(n4[6]),
        .I5(DOUTADOUT[3]),
        .O(n17__27_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__56_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n17__56_carry_n_0,n17__56_carry_n_1,n17__56_carry_n_2,n17__56_carry_n_3,n17__56_carry_n_4,n17__56_carry_n_5,n17__56_carry_n_6,n17__56_carry_n_7}),
        .DI({n17__56_carry_i_1__0_n_0,n17__56_carry_i_2__0_n_0,n17__56_carry_i_3__0_n_0,n17__56_carry_i_4__0_n_0,n17__56_carry_i_5__0_n_0,n17__56_carry_i_6__0_n_0,n17__56_carry_i_7__0_n_0,1'b0}),
        .O({n17__56_carry_n_8,n17__56_carry_n_9,n17__56_carry_n_10,n17__56_carry_n_11,n17__56_carry_n_12,n17__56_carry_n_13,n17__56_carry_n_14,n17__56_carry_n_15}),
        .S({n17__56_carry_i_8__0_n_0,n17__56_carry_i_9__0_n_0,n17__56_carry_i_10__0_n_0,n17__56_carry_i_11__0_n_0,n17__56_carry_i_12__0_n_0,n17__56_carry_i_13__0_n_0,n17__56_carry_i_14__0_n_0,n17__56_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__56_carry__0
       (.CI(n17__56_carry_n_0),
        .CI_TOP(1'b0),
        .CO(NLW_n17__56_carry__0_CO_UNCONNECTED[7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_n17__56_carry__0_O_UNCONNECTED[7:1],n17__56_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n17__56_carry__0_i_1__0_n_0}));
  LUT4 #(
    .INIT(16'hE53F)) 
    n17__56_carry__0_i_1__0
       (.I0(DOUTADOUT[6]),
        .I1(n4[6]),
        .I2(DOUTADOUT[7]),
        .I3(n4[7]),
        .O(n17__56_carry__0_i_1__0_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n17__56_carry_i_10__0
       (.I0(n4[3]),
        .I1(n4[4]),
        .I2(DOUTADOUT[7]),
        .I3(n4[5]),
        .I4(DOUTADOUT[6]),
        .O(n17__56_carry_i_10__0_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n17__56_carry_i_11__0
       (.I0(n4[2]),
        .I1(n4[3]),
        .I2(DOUTADOUT[7]),
        .I3(n4[4]),
        .I4(DOUTADOUT[6]),
        .O(n17__56_carry_i_11__0_n_0));
  LUT5 #(
    .INIT(32'h9F606060)) 
    n17__56_carry_i_12__0
       (.I0(n4[1]),
        .I1(n4[2]),
        .I2(DOUTADOUT[7]),
        .I3(n4[3]),
        .I4(DOUTADOUT[6]),
        .O(n17__56_carry_i_12__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__56_carry_i_13__0
       (.I0(DOUTADOUT[7]),
        .I1(n4[1]),
        .I2(DOUTADOUT[6]),
        .I3(n4[2]),
        .O(n17__56_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h8777)) 
    n17__56_carry_i_14__0
       (.I0(DOUTADOUT[7]),
        .I1(n4[0]),
        .I2(DOUTADOUT[6]),
        .I3(n4[1]),
        .O(n17__56_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__56_carry_i_15__0
       (.I0(n4[0]),
        .I1(DOUTADOUT[6]),
        .O(n17__56_carry_i_15__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__56_carry_i_1__0
       (.I0(DOUTADOUT[7]),
        .I1(n4[5]),
        .I2(DOUTADOUT[6]),
        .I3(n4[6]),
        .O(n17__56_carry_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__56_carry_i_2__0
       (.I0(DOUTADOUT[7]),
        .I1(n4[4]),
        .I2(DOUTADOUT[6]),
        .I3(n4[5]),
        .O(n17__56_carry_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__56_carry_i_3__0
       (.I0(DOUTADOUT[7]),
        .I1(n4[3]),
        .I2(DOUTADOUT[6]),
        .I3(n4[4]),
        .O(n17__56_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__56_carry_i_4__0
       (.I0(DOUTADOUT[7]),
        .I1(n4[2]),
        .I2(DOUTADOUT[6]),
        .I3(n4[3]),
        .O(n17__56_carry_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n17__56_carry_i_5__0
       (.I0(n4[1]),
        .I1(DOUTADOUT[7]),
        .O(n17__56_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__56_carry_i_6__0
       (.I0(DOUTADOUT[7]),
        .I1(n4[1]),
        .O(n17__56_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n17__56_carry_i_7__0
       (.I0(n4[0]),
        .I1(DOUTADOUT[7]),
        .O(n17__56_carry_i_7__0_n_0));
  LUT5 #(
    .INIT(32'h738CC0C0)) 
    n17__56_carry_i_8__0
       (.I0(n4[5]),
        .I1(n4[6]),
        .I2(DOUTADOUT[7]),
        .I3(n4[7]),
        .I4(DOUTADOUT[6]),
        .O(n17__56_carry_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n17__56_carry_i_9__0
       (.I0(n4[4]),
        .I1(n4[5]),
        .I2(DOUTADOUT[7]),
        .I3(n4[6]),
        .I4(DOUTADOUT[6]),
        .O(n17__56_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__81_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n17__81_carry_n_0,n17__81_carry_n_1,n17__81_carry_n_2,n17__81_carry_n_3,n17__81_carry_n_4,n17__81_carry_n_5,n17__81_carry_n_6,n17__81_carry_n_7}),
        .DI({n17__81_carry_i_1__0_n_0,n17__81_carry_i_2__0_n_0,n17__81_carry_i_3__0_n_0,n17__81_carry_i_4__0_n_0,n17__81_carry_i_5__0_n_0,n17__81_carry_i_6__0_n_0,n17__81_carry_i_7__0_n_0,1'b0}),
        .O({n17[10:7],NLW_n17__81_carry_O_UNCONNECTED[3:0]}),
        .S({n17__81_carry_i_8__0_n_0,n17__81_carry_i_9__0_n_0,n17__81_carry_i_10__0_n_0,n17__81_carry_i_11__0_n_0,n17__81_carry_i_12__0_n_0,n17__81_carry_i_13__0_n_0,n17__81_carry_i_14__0_n_0,n17__81_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__81_carry__0
       (.CI(n17__81_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n17__81_carry__0_CO_UNCONNECTED[7:3],n17__81_carry__0_n_5,n17__81_carry__0_n_6,n17__81_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n17__81_carry__0_i_1__0_n_0,n17__81_carry__0_i_2__0_n_0,n17__81_carry__0_i_3__0_n_0}),
        .O({NLW_n17__81_carry__0_O_UNCONNECTED[7:4],n17[14:11]}),
        .S({1'b0,1'b0,1'b0,1'b0,n17__81_carry__0_i_4__0_n_0,n17__81_carry__0_i_5__0_n_0,n17__81_carry__0_i_6__0_n_0,n17__81_carry__0_i_7__0_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry__0_i_1__0
       (.I0(n17__27_carry__0_n_14),
        .I1(n17__56_carry_n_9),
        .O(n17__81_carry__0_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry__0_i_2__0
       (.I0(n17__27_carry__0_n_15),
        .I1(n17__56_carry_n_10),
        .O(n17__81_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry__0_i_3__0
       (.I0(n17__56_carry_n_11),
        .I1(n17__27_carry_n_8),
        .I2(n17__0_carry__0_n_5),
        .O(n17__81_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n17__81_carry__0_i_4__0
       (.I0(n17__27_carry__0_n_5),
        .I1(n17__56_carry_n_8),
        .I2(n17__56_carry__0_n_15),
        .O(n17__81_carry__0_i_4__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n17__81_carry__0_i_5__0
       (.I0(n17__27_carry__0_n_14),
        .I1(n17__56_carry_n_9),
        .I2(n17__56_carry_n_8),
        .I3(n17__27_carry__0_n_5),
        .O(n17__81_carry__0_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n17__81_carry__0_i_6__0
       (.I0(n17__27_carry__0_n_15),
        .I1(n17__56_carry_n_10),
        .I2(n17__56_carry_n_9),
        .I3(n17__27_carry__0_n_14),
        .O(n17__81_carry__0_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n17__81_carry__0_i_7__0
       (.I0(n17__0_carry__0_n_5),
        .I1(n17__27_carry_n_8),
        .I2(n17__56_carry_n_11),
        .I3(n17__56_carry_n_10),
        .I4(n17__27_carry__0_n_15),
        .O(n17__81_carry__0_i_7__0_n_0));
  (* HLUTNM = "lutpair10" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_10__0
       (.I0(n17__56_carry_n_13),
        .I1(n17__27_carry_n_10),
        .I2(n17__0_carry__0_n_15),
        .I3(n17__81_carry_i_3__0_n_0),
        .O(n17__81_carry_i_10__0_n_0));
  (* HLUTNM = "lutpair9" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_11__0
       (.I0(n17__56_carry_n_14),
        .I1(n17__27_carry_n_11),
        .I2(n17__0_carry_n_8),
        .I3(n17__81_carry_i_4__0_n_0),
        .O(n17__81_carry_i_11__0_n_0));
  (* HLUTNM = "lutpair8" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_12__0
       (.I0(n17__56_carry_n_15),
        .I1(n17__27_carry_n_12),
        .I2(n17__0_carry_n_9),
        .I3(n17__81_carry_i_5__0_n_0),
        .O(n17__81_carry_i_12__0_n_0));
  (* HLUTNM = "lutpair82" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n17__81_carry_i_13__0
       (.I0(n17__27_carry_n_13),
        .I1(n17__0_carry_n_10),
        .I2(n17__0_carry_n_11),
        .I3(n17__27_carry_n_14),
        .O(n17__81_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n17__81_carry_i_14__0
       (.I0(n17__0_carry_n_12),
        .I1(n17__27_carry_n_15),
        .I2(n17__27_carry_n_14),
        .I3(n17__0_carry_n_11),
        .O(n17__81_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n17__81_carry_i_15__0
       (.I0(n17__0_carry_n_12),
        .I1(n17__27_carry_n_15),
        .O(n17__81_carry_i_15__0_n_0));
  (* HLUTNM = "lutpair11" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry_i_1__0
       (.I0(n17__56_carry_n_12),
        .I1(n17__27_carry_n_9),
        .I2(n17__0_carry__0_n_14),
        .O(n17__81_carry_i_1__0_n_0));
  (* HLUTNM = "lutpair10" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry_i_2__0
       (.I0(n17__56_carry_n_13),
        .I1(n17__27_carry_n_10),
        .I2(n17__0_carry__0_n_15),
        .O(n17__81_carry_i_2__0_n_0));
  (* HLUTNM = "lutpair9" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry_i_3__0
       (.I0(n17__56_carry_n_14),
        .I1(n17__27_carry_n_11),
        .I2(n17__0_carry_n_8),
        .O(n17__81_carry_i_3__0_n_0));
  (* HLUTNM = "lutpair8" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry_i_4__0
       (.I0(n17__56_carry_n_15),
        .I1(n17__27_carry_n_12),
        .I2(n17__0_carry_n_9),
        .O(n17__81_carry_i_4__0_n_0));
  (* HLUTNM = "lutpair82" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry_i_5__0
       (.I0(n17__27_carry_n_13),
        .I1(n17__0_carry_n_10),
        .O(n17__81_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry_i_6__0
       (.I0(n17__0_carry_n_11),
        .I1(n17__27_carry_n_14),
        .O(n17__81_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry_i_7__0
       (.I0(n17__0_carry_n_12),
        .I1(n17__27_carry_n_15),
        .O(n17__81_carry_i_7__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_8__0
       (.I0(n17__81_carry_i_1__0_n_0),
        .I1(n17__27_carry_n_8),
        .I2(n17__56_carry_n_11),
        .I3(n17__0_carry__0_n_5),
        .O(n17__81_carry_i_8__0_n_0));
  (* HLUTNM = "lutpair11" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_9__0
       (.I0(n17__56_carry_n_12),
        .I1(n17__27_carry_n_9),
        .I2(n17__0_carry__0_n_14),
        .I3(n17__81_carry_i_2__0_n_0),
        .O(n17__81_carry_i_9__0_n_0));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[14]),
        .Q(n19_reg_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__0
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[13]),
        .Q(n19_reg__0_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__1
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[12]),
        .Q(n19_reg__1_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__2
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[11]),
        .Q(n19_reg__2_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__3
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[10]),
        .Q(n19_reg__3_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__4
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[9]),
        .Q(n19_reg__4_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__5
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[8]),
        .Q(n19_reg__5_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__6
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[7]),
        .Q(n19_reg__6_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[0]),
        .Q(\n1_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[10]),
        .Q(n2[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[11]),
        .Q(n2[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[12]),
        .Q(n2[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[13]),
        .Q(n2[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[14]),
        .Q(n2[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[15]),
        .Q(n2[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[1]),
        .Q(\n1_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[2]),
        .Q(\n1_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[3]),
        .Q(\n1_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[4]),
        .Q(\n1_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[5]),
        .Q(\n1_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[6]),
        .Q(\n1_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[7]),
        .Q(\n1_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[8]),
        .Q(n2[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[9]),
        .Q(n2[1]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n20_carry
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({NLW_n20_carry_CO_UNCONNECTED[7],n20_carry_n_1,n20_carry_n_2,n20_carry_n_3,n20_carry_n_4,n20_carry_n_5,n20_carry_n_6,n20_carry_n_7}),
        .DI({1'b0,\n16_reg_n_0_[6] ,\n16_reg_n_0_[5] ,\n16_reg_n_0_[4] ,\n16_reg_n_0_[3] ,\n16_reg_n_0_[2] ,\n16_reg_n_0_[1] ,\n16_reg_n_0_[0] }),
        .O(n202_out),
        .S({n20_carry_i_1__1_n_0,n20_carry_i_2__1_n_0,n20_carry_i_3__1_n_0,n20_carry_i_4__1_n_0,n20_carry_i_5__1_n_0,n20_carry_i_6__1_n_0,n20_carry_i_7__1_n_0,n20_carry_i_8__1_n_0}));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_1__1
       (.I0(\n16_reg_n_0_[7] ),
        .I1(n19_reg_n_0),
        .O(n20_carry_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_2__1
       (.I0(\n16_reg_n_0_[6] ),
        .I1(n19_reg__0_n_0),
        .O(n20_carry_i_2__1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_3__1
       (.I0(\n16_reg_n_0_[5] ),
        .I1(n19_reg__1_n_0),
        .O(n20_carry_i_3__1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_4__1
       (.I0(\n16_reg_n_0_[4] ),
        .I1(n19_reg__2_n_0),
        .O(n20_carry_i_4__1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_5__1
       (.I0(\n16_reg_n_0_[3] ),
        .I1(n19_reg__3_n_0),
        .O(n20_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_6__1
       (.I0(\n16_reg_n_0_[2] ),
        .I1(n19_reg__4_n_0),
        .O(n20_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_7__1
       (.I0(\n16_reg_n_0_[1] ),
        .I1(n19_reg__5_n_0),
        .O(n20_carry_i_7__1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_8__1
       (.I0(\n16_reg_n_0_[0] ),
        .I1(n19_reg__6_n_0),
        .O(n20_carry_i_8__1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[0]),
        .Q(n21[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[1]),
        .Q(n21[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[2]),
        .Q(n21[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[3]),
        .Q(n21[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[4]),
        .Q(n21[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[5]),
        .Q(n21[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[6]),
        .Q(n21[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[7]),
        .Q(n21[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[15]),
        .Q(n22_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__0
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[14]),
        .Q(n22__0_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__0_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n22__0_carry_n_0,n22__0_carry_n_1,n22__0_carry_n_2,n22__0_carry_n_3,n22__0_carry_n_4,n22__0_carry_n_5,n22__0_carry_n_6,n22__0_carry_n_7}),
        .DI({n22__0_carry_i_1__0_n_0,n22__0_carry_i_2__0_n_0,n22__0_carry_i_3__0_n_0,n22__0_carry_i_4__0_n_0,n22__0_carry_i_5__0_n_0,n22__0_carry_i_6__0_n_0,n22__0_carry_i_7__0_n_0,1'b0}),
        .O({n22__0_carry_n_8,n22__0_carry_n_9,n22__0_carry_n_10,n22__0_carry_n_11,n22__0_carry_n_12,NLW_n22__0_carry_O_UNCONNECTED[2:0]}),
        .S({n22__0_carry_i_8__0_n_0,n22__0_carry_i_9__0_n_0,n22__0_carry_i_10__0_n_0,n22__0_carry_i_11__0_n_0,n22__0_carry_i_12__0_n_0,n22__0_carry_i_13__0_n_0,n22__0_carry_i_14__0_n_0,n22__0_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__0_carry__0
       (.CI(n22__0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n22__0_carry__0_CO_UNCONNECTED[7:3],n22__0_carry__0_n_5,NLW_n22__0_carry__0_CO_UNCONNECTED[1],n22__0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n22__0_carry__0_i_1__0_n_0,n22__0_carry__0_i_2__0_n_0}),
        .O({NLW_n22__0_carry__0_O_UNCONNECTED[7:2],n22__0_carry__0_n_14,n22__0_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n22__0_carry__0_i_3__0_n_0,n22__0_carry__0_i_4__0_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__0_carry__0_i_1__0
       (.I0(DOUTADOUT[1]),
        .I1(n22_n_0),
        .I2(DOUTADOUT[2]),
        .I3(n22__0_n_0),
        .O(n22__0_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n22__0_carry__0_i_2__0
       (.I0(DOUTADOUT[2]),
        .I1(n22__1_n_0),
        .I2(DOUTADOUT[1]),
        .I3(n22__0_n_0),
        .I4(DOUTADOUT[0]),
        .I5(n22_n_0),
        .O(n22__0_carry__0_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n22__0_carry__0_i_3__0
       (.I0(n22__0_n_0),
        .I1(DOUTADOUT[1]),
        .I2(DOUTADOUT[2]),
        .I3(n22_n_0),
        .O(n22__0_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n22__0_carry__0_i_4__0
       (.I0(DOUTADOUT[0]),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(DOUTADOUT[2]),
        .I4(n22_n_0),
        .I5(DOUTADOUT[1]),
        .O(n22__0_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__0_carry_i_10__0
       (.I0(n22__0_carry_i_3__0_n_0),
        .I1(DOUTADOUT[1]),
        .I2(n22__2_n_0),
        .I3(n22__0_carry_i_18__0_n_0),
        .I4(n22__1_n_0),
        .I5(DOUTADOUT[0]),
        .O(n22__0_carry_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__0_carry_i_11__0
       (.I0(n22__0_carry_i_4__0_n_0),
        .I1(DOUTADOUT[1]),
        .I2(n22__3_n_0),
        .I3(n22__0_carry_i_19__0_n_0),
        .I4(n22__2_n_0),
        .I5(DOUTADOUT[0]),
        .O(n22__0_carry_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n22__0_carry_i_12__0
       (.I0(n22__4_n_0),
        .I1(n22__0_carry_i_20__0_n_0),
        .I2(n22__5_n_0),
        .I3(DOUTADOUT[1]),
        .I4(n22__6_n_0),
        .I5(DOUTADOUT[2]),
        .O(n22__0_carry_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n22__0_carry_i_13__0
       (.I0(n22__6_n_0),
        .I1(DOUTADOUT[2]),
        .I2(n22__5_n_0),
        .I3(DOUTADOUT[1]),
        .I4(DOUTADOUT[0]),
        .I5(n22__4_n_0),
        .O(n22__0_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__0_carry_i_14__0
       (.I0(DOUTADOUT[0]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[1]),
        .I3(n22__6_n_0),
        .O(n22__0_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__0_carry_i_15__0
       (.I0(n22__6_n_0),
        .I1(DOUTADOUT[0]),
        .O(n22__0_carry_i_15__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_16__0
       (.I0(n22__1_n_0),
        .I1(DOUTADOUT[2]),
        .O(n22__0_carry_i_16__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_17__0
       (.I0(n22__2_n_0),
        .I1(DOUTADOUT[2]),
        .O(n22__0_carry_i_17__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_18__0
       (.I0(n22__3_n_0),
        .I1(DOUTADOUT[2]),
        .O(n22__0_carry_i_18__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_19__0
       (.I0(n22__4_n_0),
        .I1(DOUTADOUT[2]),
        .O(n22__0_carry_i_19__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__0_carry_i_1__0
       (.I0(DOUTADOUT[2]),
        .I1(n22__2_n_0),
        .I2(DOUTADOUT[1]),
        .I3(n22__1_n_0),
        .I4(DOUTADOUT[0]),
        .I5(n22__0_n_0),
        .O(n22__0_carry_i_1__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_20__0
       (.I0(n22__3_n_0),
        .I1(DOUTADOUT[0]),
        .O(n22__0_carry_i_20__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__0_carry_i_2__0
       (.I0(DOUTADOUT[2]),
        .I1(n22__3_n_0),
        .I2(DOUTADOUT[1]),
        .I3(n22__2_n_0),
        .I4(DOUTADOUT[0]),
        .I5(n22__1_n_0),
        .O(n22__0_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__0_carry_i_3__0
       (.I0(DOUTADOUT[2]),
        .I1(n22__4_n_0),
        .I2(DOUTADOUT[1]),
        .I3(n22__3_n_0),
        .I4(DOUTADOUT[0]),
        .I5(n22__2_n_0),
        .O(n22__0_carry_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__0_carry_i_4__0
       (.I0(DOUTADOUT[2]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[1]),
        .I3(n22__4_n_0),
        .I4(DOUTADOUT[0]),
        .I5(n22__3_n_0),
        .O(n22__0_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n22__0_carry_i_5__0
       (.I0(DOUTADOUT[1]),
        .I1(n22__4_n_0),
        .I2(DOUTADOUT[2]),
        .I3(n22__5_n_0),
        .I4(n22__3_n_0),
        .I5(DOUTADOUT[0]),
        .O(n22__0_carry_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__0_carry_i_6__0
       (.I0(DOUTADOUT[1]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[2]),
        .I3(n22__6_n_0),
        .O(n22__0_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__0_carry_i_7__0
       (.I0(DOUTADOUT[0]),
        .I1(n22__5_n_0),
        .O(n22__0_carry_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n22__0_carry_i_8__0
       (.I0(n22__0_carry_i_1__0_n_0),
        .I1(DOUTADOUT[1]),
        .I2(n22__0_n_0),
        .I3(n22__0_carry_i_16__0_n_0),
        .I4(n22_n_0),
        .I5(DOUTADOUT[0]),
        .O(n22__0_carry_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__0_carry_i_9__0
       (.I0(n22__0_carry_i_2__0_n_0),
        .I1(DOUTADOUT[1]),
        .I2(n22__1_n_0),
        .I3(n22__0_carry_i_17__0_n_0),
        .I4(n22__0_n_0),
        .I5(DOUTADOUT[0]),
        .O(n22__0_carry_i_9__0_n_0));
  FDRE #(
    .INIT(1'b0)) 
    n22__1
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[13]),
        .Q(n22__1_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__2
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[12]),
        .Q(n22__2_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__27_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n22__27_carry_n_0,n22__27_carry_n_1,n22__27_carry_n_2,n22__27_carry_n_3,n22__27_carry_n_4,n22__27_carry_n_5,n22__27_carry_n_6,n22__27_carry_n_7}),
        .DI({n22__27_carry_i_1__0_n_0,n22__27_carry_i_2__0_n_0,n22__27_carry_i_3__0_n_0,n22__27_carry_i_4__0_n_0,n22__27_carry_i_5__0_n_0,n22__27_carry_i_6__0_n_0,n22__27_carry_i_7__0_n_0,1'b0}),
        .O({n22__27_carry_n_8,n22__27_carry_n_9,n22__27_carry_n_10,n22__27_carry_n_11,n22__27_carry_n_12,n22__27_carry_n_13,n22__27_carry_n_14,n22__27_carry_n_15}),
        .S({n22__27_carry_i_8__0_n_0,n22__27_carry_i_9__0_n_0,n22__27_carry_i_10__0_n_0,n22__27_carry_i_11__0_n_0,n22__27_carry_i_12__0_n_0,n22__27_carry_i_13__0_n_0,n22__27_carry_i_14__0_n_0,n22__27_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__27_carry__0
       (.CI(n22__27_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n22__27_carry__0_CO_UNCONNECTED[7:3],n22__27_carry__0_n_5,NLW_n22__27_carry__0_CO_UNCONNECTED[1],n22__27_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n22__27_carry__0_i_1__0_n_0,n22__27_carry__0_i_2__0_n_0}),
        .O({NLW_n22__27_carry__0_O_UNCONNECTED[7:2],n22__27_carry__0_n_14,n22__27_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n22__27_carry__0_i_3__0_n_0,n22__27_carry__0_i_4__0_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__27_carry__0_i_1__0
       (.I0(DOUTADOUT[4]),
        .I1(n22_n_0),
        .I2(DOUTADOUT[5]),
        .I3(n22__0_n_0),
        .O(n22__27_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n22__27_carry__0_i_2__0
       (.I0(DOUTADOUT[5]),
        .I1(n22__1_n_0),
        .I2(DOUTADOUT[4]),
        .I3(n22__0_n_0),
        .I4(DOUTADOUT[3]),
        .I5(n22_n_0),
        .O(n22__27_carry__0_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n22__27_carry__0_i_3__0
       (.I0(n22__0_n_0),
        .I1(DOUTADOUT[4]),
        .I2(DOUTADOUT[5]),
        .I3(n22_n_0),
        .O(n22__27_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n22__27_carry__0_i_4__0
       (.I0(DOUTADOUT[3]),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(DOUTADOUT[5]),
        .I4(n22_n_0),
        .I5(DOUTADOUT[4]),
        .O(n22__27_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__27_carry_i_10__0
       (.I0(n22__27_carry_i_3__0_n_0),
        .I1(DOUTADOUT[4]),
        .I2(n22__2_n_0),
        .I3(n22__27_carry_i_18__0_n_0),
        .I4(n22__1_n_0),
        .I5(DOUTADOUT[3]),
        .O(n22__27_carry_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__27_carry_i_11__0
       (.I0(n22__27_carry_i_4__0_n_0),
        .I1(DOUTADOUT[4]),
        .I2(n22__3_n_0),
        .I3(n22__27_carry_i_19__0_n_0),
        .I4(n22__2_n_0),
        .I5(DOUTADOUT[3]),
        .O(n22__27_carry_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n22__27_carry_i_12__0
       (.I0(n22__4_n_0),
        .I1(n22__27_carry_i_20__0_n_0),
        .I2(n22__5_n_0),
        .I3(DOUTADOUT[4]),
        .I4(n22__6_n_0),
        .I5(DOUTADOUT[5]),
        .O(n22__27_carry_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n22__27_carry_i_13__0
       (.I0(n22__6_n_0),
        .I1(DOUTADOUT[5]),
        .I2(n22__5_n_0),
        .I3(DOUTADOUT[4]),
        .I4(DOUTADOUT[3]),
        .I5(n22__4_n_0),
        .O(n22__27_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__27_carry_i_14__0
       (.I0(DOUTADOUT[3]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[4]),
        .I3(n22__6_n_0),
        .O(n22__27_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__27_carry_i_15__0
       (.I0(n22__6_n_0),
        .I1(DOUTADOUT[3]),
        .O(n22__27_carry_i_15__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_16__0
       (.I0(n22__1_n_0),
        .I1(DOUTADOUT[5]),
        .O(n22__27_carry_i_16__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_17__0
       (.I0(n22__2_n_0),
        .I1(DOUTADOUT[5]),
        .O(n22__27_carry_i_17__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_18__0
       (.I0(n22__3_n_0),
        .I1(DOUTADOUT[5]),
        .O(n22__27_carry_i_18__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_19__0
       (.I0(n22__4_n_0),
        .I1(DOUTADOUT[5]),
        .O(n22__27_carry_i_19__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__27_carry_i_1__0
       (.I0(DOUTADOUT[5]),
        .I1(n22__2_n_0),
        .I2(DOUTADOUT[4]),
        .I3(n22__1_n_0),
        .I4(DOUTADOUT[3]),
        .I5(n22__0_n_0),
        .O(n22__27_carry_i_1__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_20__0
       (.I0(n22__3_n_0),
        .I1(DOUTADOUT[3]),
        .O(n22__27_carry_i_20__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__27_carry_i_2__0
       (.I0(DOUTADOUT[5]),
        .I1(n22__3_n_0),
        .I2(DOUTADOUT[4]),
        .I3(n22__2_n_0),
        .I4(DOUTADOUT[3]),
        .I5(n22__1_n_0),
        .O(n22__27_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__27_carry_i_3__0
       (.I0(DOUTADOUT[5]),
        .I1(n22__4_n_0),
        .I2(DOUTADOUT[4]),
        .I3(n22__3_n_0),
        .I4(DOUTADOUT[3]),
        .I5(n22__2_n_0),
        .O(n22__27_carry_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__27_carry_i_4__0
       (.I0(DOUTADOUT[5]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[4]),
        .I3(n22__4_n_0),
        .I4(DOUTADOUT[3]),
        .I5(n22__3_n_0),
        .O(n22__27_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n22__27_carry_i_5__0
       (.I0(DOUTADOUT[4]),
        .I1(n22__4_n_0),
        .I2(DOUTADOUT[5]),
        .I3(n22__5_n_0),
        .I4(n22__3_n_0),
        .I5(DOUTADOUT[3]),
        .O(n22__27_carry_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__27_carry_i_6__0
       (.I0(DOUTADOUT[4]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[5]),
        .I3(n22__6_n_0),
        .O(n22__27_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__27_carry_i_7__0
       (.I0(DOUTADOUT[3]),
        .I1(n22__5_n_0),
        .O(n22__27_carry_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n22__27_carry_i_8__0
       (.I0(n22__27_carry_i_1__0_n_0),
        .I1(DOUTADOUT[4]),
        .I2(n22__0_n_0),
        .I3(n22__27_carry_i_16__0_n_0),
        .I4(n22_n_0),
        .I5(DOUTADOUT[3]),
        .O(n22__27_carry_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__27_carry_i_9__0
       (.I0(n22__27_carry_i_2__0_n_0),
        .I1(DOUTADOUT[4]),
        .I2(n22__1_n_0),
        .I3(n22__27_carry_i_17__0_n_0),
        .I4(n22__0_n_0),
        .I5(DOUTADOUT[3]),
        .O(n22__27_carry_i_9__0_n_0));
  FDRE #(
    .INIT(1'b0)) 
    n22__3
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[11]),
        .Q(n22__3_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__4
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[10]),
        .Q(n22__4_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__5
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[9]),
        .Q(n22__5_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__56_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n22__56_carry_n_0,n22__56_carry_n_1,n22__56_carry_n_2,n22__56_carry_n_3,n22__56_carry_n_4,n22__56_carry_n_5,n22__56_carry_n_6,n22__56_carry_n_7}),
        .DI({n22__56_carry_i_1__0_n_0,n22__56_carry_i_2__0_n_0,n22__56_carry_i_3__0_n_0,n22__56_carry_i_4__0_n_0,n22__56_carry_i_5__0_n_0,n22__56_carry_i_6__0_n_0,n22__56_carry_i_7__0_n_0,1'b0}),
        .O({n22__56_carry_n_8,n22__56_carry_n_9,n22__56_carry_n_10,n22__56_carry_n_11,n22__56_carry_n_12,n22__56_carry_n_13,n22__56_carry_n_14,n22__56_carry_n_15}),
        .S({n22__56_carry_i_8__0_n_0,n22__56_carry_i_9__0_n_0,n22__56_carry_i_10__0_n_0,n22__56_carry_i_11__0_n_0,n22__56_carry_i_12__0_n_0,n22__56_carry_i_13__0_n_0,n22__56_carry_i_14__0_n_0,n22__56_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__56_carry__0
       (.CI(n22__56_carry_n_0),
        .CI_TOP(1'b0),
        .CO(NLW_n22__56_carry__0_CO_UNCONNECTED[7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_n22__56_carry__0_O_UNCONNECTED[7:1],n22__56_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n22__56_carry__0_i_1__0_n_0}));
  LUT4 #(
    .INIT(16'hE53F)) 
    n22__56_carry__0_i_1__0
       (.I0(DOUTADOUT[6]),
        .I1(n22__0_n_0),
        .I2(DOUTADOUT[7]),
        .I3(n22_n_0),
        .O(n22__56_carry__0_i_1__0_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n22__56_carry_i_10__0
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(DOUTADOUT[7]),
        .I3(n22__1_n_0),
        .I4(DOUTADOUT[6]),
        .O(n22__56_carry_i_10__0_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n22__56_carry_i_11__0
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(DOUTADOUT[7]),
        .I3(n22__2_n_0),
        .I4(DOUTADOUT[6]),
        .O(n22__56_carry_i_11__0_n_0));
  LUT5 #(
    .INIT(32'h9F606060)) 
    n22__56_carry_i_12__0
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(DOUTADOUT[7]),
        .I3(n22__3_n_0),
        .I4(DOUTADOUT[6]),
        .O(n22__56_carry_i_12__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__56_carry_i_13__0
       (.I0(DOUTADOUT[7]),
        .I1(n22__5_n_0),
        .I2(DOUTADOUT[6]),
        .I3(n22__4_n_0),
        .O(n22__56_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h8777)) 
    n22__56_carry_i_14__0
       (.I0(DOUTADOUT[7]),
        .I1(n22__6_n_0),
        .I2(DOUTADOUT[6]),
        .I3(n22__5_n_0),
        .O(n22__56_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__56_carry_i_15__0
       (.I0(n22__6_n_0),
        .I1(DOUTADOUT[6]),
        .O(n22__56_carry_i_15__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__56_carry_i_1__0
       (.I0(DOUTADOUT[7]),
        .I1(n22__1_n_0),
        .I2(DOUTADOUT[6]),
        .I3(n22__0_n_0),
        .O(n22__56_carry_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__56_carry_i_2__0
       (.I0(DOUTADOUT[7]),
        .I1(n22__2_n_0),
        .I2(DOUTADOUT[6]),
        .I3(n22__1_n_0),
        .O(n22__56_carry_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__56_carry_i_3__0
       (.I0(DOUTADOUT[7]),
        .I1(n22__3_n_0),
        .I2(DOUTADOUT[6]),
        .I3(n22__2_n_0),
        .O(n22__56_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__56_carry_i_4__0
       (.I0(DOUTADOUT[7]),
        .I1(n22__4_n_0),
        .I2(DOUTADOUT[6]),
        .I3(n22__3_n_0),
        .O(n22__56_carry_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n22__56_carry_i_5__0
       (.I0(n22__5_n_0),
        .I1(DOUTADOUT[7]),
        .O(n22__56_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__56_carry_i_6__0
       (.I0(DOUTADOUT[7]),
        .I1(n22__5_n_0),
        .O(n22__56_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n22__56_carry_i_7__0
       (.I0(n22__6_n_0),
        .I1(DOUTADOUT[7]),
        .O(n22__56_carry_i_7__0_n_0));
  LUT5 #(
    .INIT(32'h738CC0C0)) 
    n22__56_carry_i_8__0
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(DOUTADOUT[7]),
        .I3(n22_n_0),
        .I4(DOUTADOUT[6]),
        .O(n22__56_carry_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n22__56_carry_i_9__0
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(DOUTADOUT[7]),
        .I3(n22__0_n_0),
        .I4(DOUTADOUT[6]),
        .O(n22__56_carry_i_9__0_n_0));
  FDRE #(
    .INIT(1'b0)) 
    n22__6
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[8]),
        .Q(n22__6_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__81_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n22__81_carry_n_0,n22__81_carry_n_1,n22__81_carry_n_2,n22__81_carry_n_3,n22__81_carry_n_4,n22__81_carry_n_5,n22__81_carry_n_6,n22__81_carry_n_7}),
        .DI({n22__81_carry_i_1__0_n_0,n22__81_carry_i_2__0_n_0,n22__81_carry_i_3__0_n_0,n22__81_carry_i_4__0_n_0,n22__81_carry_i_5__0_n_0,n22__81_carry_i_6__0_n_0,n22__81_carry_i_7__0_n_0,1'b0}),
        .O({n23[3:0],NLW_n22__81_carry_O_UNCONNECTED[3:0]}),
        .S({n22__81_carry_i_8__0_n_0,n22__81_carry_i_9__0_n_0,n22__81_carry_i_10__0_n_0,n22__81_carry_i_11__0_n_0,n22__81_carry_i_12__0_n_0,n22__81_carry_i_13__0_n_0,n22__81_carry_i_14__0_n_0,n22__81_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__81_carry__0
       (.CI(n22__81_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n22__81_carry__0_CO_UNCONNECTED[7:3],n22__81_carry__0_n_5,n22__81_carry__0_n_6,n22__81_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n22__81_carry__0_i_1__0_n_0,n22__81_carry__0_i_2__0_n_0,n22__81_carry__0_i_3__0_n_0}),
        .O({NLW_n22__81_carry__0_O_UNCONNECTED[7:4],n23[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n22__81_carry__0_i_4__0_n_0,n22__81_carry__0_i_5__0_n_0,n22__81_carry__0_i_6__0_n_0,n22__81_carry__0_i_7__0_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry__0_i_1__0
       (.I0(n22__27_carry__0_n_14),
        .I1(n22__56_carry_n_9),
        .O(n22__81_carry__0_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry__0_i_2__0
       (.I0(n22__27_carry__0_n_15),
        .I1(n22__56_carry_n_10),
        .O(n22__81_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry__0_i_3__0
       (.I0(n22__56_carry_n_11),
        .I1(n22__27_carry_n_8),
        .I2(n22__0_carry__0_n_5),
        .O(n22__81_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n22__81_carry__0_i_4__0
       (.I0(n22__27_carry__0_n_5),
        .I1(n22__56_carry_n_8),
        .I2(n22__56_carry__0_n_15),
        .O(n22__81_carry__0_i_4__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n22__81_carry__0_i_5__0
       (.I0(n22__27_carry__0_n_14),
        .I1(n22__56_carry_n_9),
        .I2(n22__56_carry_n_8),
        .I3(n22__27_carry__0_n_5),
        .O(n22__81_carry__0_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n22__81_carry__0_i_6__0
       (.I0(n22__27_carry__0_n_15),
        .I1(n22__56_carry_n_10),
        .I2(n22__56_carry_n_9),
        .I3(n22__27_carry__0_n_14),
        .O(n22__81_carry__0_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n22__81_carry__0_i_7__0
       (.I0(n22__0_carry__0_n_5),
        .I1(n22__27_carry_n_8),
        .I2(n22__56_carry_n_11),
        .I3(n22__56_carry_n_10),
        .I4(n22__27_carry__0_n_15),
        .O(n22__81_carry__0_i_7__0_n_0));
  (* HLUTNM = "lutpair6" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_10__0
       (.I0(n22__56_carry_n_13),
        .I1(n22__27_carry_n_10),
        .I2(n22__0_carry__0_n_15),
        .I3(n22__81_carry_i_3__0_n_0),
        .O(n22__81_carry_i_10__0_n_0));
  (* HLUTNM = "lutpair5" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_11__0
       (.I0(n22__56_carry_n_14),
        .I1(n22__27_carry_n_11),
        .I2(n22__0_carry_n_8),
        .I3(n22__81_carry_i_4__0_n_0),
        .O(n22__81_carry_i_11__0_n_0));
  (* HLUTNM = "lutpair4" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_12__0
       (.I0(n22__56_carry_n_15),
        .I1(n22__27_carry_n_12),
        .I2(n22__0_carry_n_9),
        .I3(n22__81_carry_i_5__0_n_0),
        .O(n22__81_carry_i_12__0_n_0));
  (* HLUTNM = "lutpair81" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n22__81_carry_i_13__0
       (.I0(n22__27_carry_n_13),
        .I1(n22__0_carry_n_10),
        .I2(n22__0_carry_n_11),
        .I3(n22__27_carry_n_14),
        .O(n22__81_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n22__81_carry_i_14__0
       (.I0(n22__0_carry_n_12),
        .I1(n22__27_carry_n_15),
        .I2(n22__27_carry_n_14),
        .I3(n22__0_carry_n_11),
        .O(n22__81_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n22__81_carry_i_15__0
       (.I0(n22__0_carry_n_12),
        .I1(n22__27_carry_n_15),
        .O(n22__81_carry_i_15__0_n_0));
  (* HLUTNM = "lutpair7" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry_i_1__0
       (.I0(n22__56_carry_n_12),
        .I1(n22__27_carry_n_9),
        .I2(n22__0_carry__0_n_14),
        .O(n22__81_carry_i_1__0_n_0));
  (* HLUTNM = "lutpair6" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry_i_2__0
       (.I0(n22__56_carry_n_13),
        .I1(n22__27_carry_n_10),
        .I2(n22__0_carry__0_n_15),
        .O(n22__81_carry_i_2__0_n_0));
  (* HLUTNM = "lutpair5" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry_i_3__0
       (.I0(n22__56_carry_n_14),
        .I1(n22__27_carry_n_11),
        .I2(n22__0_carry_n_8),
        .O(n22__81_carry_i_3__0_n_0));
  (* HLUTNM = "lutpair4" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry_i_4__0
       (.I0(n22__56_carry_n_15),
        .I1(n22__27_carry_n_12),
        .I2(n22__0_carry_n_9),
        .O(n22__81_carry_i_4__0_n_0));
  (* HLUTNM = "lutpair81" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry_i_5__0
       (.I0(n22__27_carry_n_13),
        .I1(n22__0_carry_n_10),
        .O(n22__81_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry_i_6__0
       (.I0(n22__0_carry_n_11),
        .I1(n22__27_carry_n_14),
        .O(n22__81_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry_i_7__0
       (.I0(n22__0_carry_n_12),
        .I1(n22__27_carry_n_15),
        .O(n22__81_carry_i_7__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_8__0
       (.I0(n22__81_carry_i_1__0_n_0),
        .I1(n22__27_carry_n_8),
        .I2(n22__56_carry_n_11),
        .I3(n22__0_carry__0_n_5),
        .O(n22__81_carry_i_8__0_n_0));
  (* HLUTNM = "lutpair7" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_9__0
       (.I0(n22__56_carry_n_12),
        .I1(n22__27_carry_n_9),
        .I2(n22__0_carry__0_n_14),
        .I3(n22__81_carry_i_2__0_n_0),
        .O(n22__81_carry_i_9__0_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[0]),
        .Q(n24[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[1]),
        .Q(n24[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[2]),
        .Q(n24[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[3]),
        .Q(n24[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[4]),
        .Q(n24[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[5]),
        .Q(n24[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[6]),
        .Q(n24[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[7]),
        .Q(n24[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__0_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__0_carry_n_0,n25__0_carry_n_1,n25__0_carry_n_2,n25__0_carry_n_3,n25__0_carry_n_4,n25__0_carry_n_5,n25__0_carry_n_6,n25__0_carry_n_7}),
        .DI({n25__0_carry_i_1__0_n_0,n25__0_carry_i_2__0_n_0,n25__0_carry_i_3__0_n_0,n25__0_carry_i_4__0_n_0,n25__0_carry_i_5__0_n_0,n25__0_carry_i_6__0_n_0,n25__0_carry_i_7__0_n_0,1'b0}),
        .O({n25__0_carry_n_8,n25__0_carry_n_9,n25__0_carry_n_10,n25__0_carry_n_11,n25__0_carry_n_12,NLW_n25__0_carry_O_UNCONNECTED[2:0]}),
        .S({n25__0_carry_i_8__0_n_0,n25__0_carry_i_9__0_n_0,n25__0_carry_i_10__0_n_0,n25__0_carry_i_11__0_n_0,n25__0_carry_i_12__0_n_0,n25__0_carry_i_13__0_n_0,n25__0_carry_i_14__0_n_0,n25__0_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__0_carry__0
       (.CI(n25__0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__0_carry__0_CO_UNCONNECTED[7:3],n25__0_carry__0_n_5,NLW_n25__0_carry__0_CO_UNCONNECTED[1],n25__0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25__0_carry__0_i_1__0_n_0,n25__0_carry__0_i_2__0_n_0}),
        .O({NLW_n25__0_carry__0_O_UNCONNECTED[7:2],n25__0_carry__0_n_14,n25__0_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n25__0_carry__0_i_3__0_n_0,n25__0_carry__0_i_4__0_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__0_carry__0_i_1__0
       (.I0(DOUTADOUT[9]),
        .I1(n4[7]),
        .I2(DOUTADOUT[10]),
        .I3(n4[6]),
        .O(n25__0_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n25__0_carry__0_i_2__0
       (.I0(DOUTADOUT[10]),
        .I1(n4[5]),
        .I2(DOUTADOUT[9]),
        .I3(n4[6]),
        .I4(DOUTADOUT[8]),
        .I5(n4[7]),
        .O(n25__0_carry__0_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n25__0_carry__0_i_3__0
       (.I0(n4[6]),
        .I1(DOUTADOUT[9]),
        .I2(DOUTADOUT[10]),
        .I3(n4[7]),
        .O(n25__0_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n25__0_carry__0_i_4__0
       (.I0(DOUTADOUT[8]),
        .I1(n4[5]),
        .I2(n4[6]),
        .I3(DOUTADOUT[10]),
        .I4(n4[7]),
        .I5(DOUTADOUT[9]),
        .O(n25__0_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__0_carry_i_10__0
       (.I0(n25__0_carry_i_3__0_n_0),
        .I1(DOUTADOUT[9]),
        .I2(n4[4]),
        .I3(n25__0_carry_i_19__0_n_0),
        .I4(n4[5]),
        .I5(DOUTADOUT[8]),
        .O(n25__0_carry_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__0_carry_i_11__0
       (.I0(n25__0_carry_i_4__0_n_0),
        .I1(DOUTADOUT[9]),
        .I2(n4[3]),
        .I3(n25__0_carry_i_20__0_n_0),
        .I4(n4[4]),
        .I5(DOUTADOUT[8]),
        .O(n25__0_carry_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n25__0_carry_i_12__0
       (.I0(n4[2]),
        .I1(n25__0_carry_i_21_n_0),
        .I2(n4[1]),
        .I3(DOUTADOUT[9]),
        .I4(n4[0]),
        .I5(DOUTADOUT[10]),
        .O(n25__0_carry_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n25__0_carry_i_13__0
       (.I0(n4[0]),
        .I1(DOUTADOUT[10]),
        .I2(n4[1]),
        .I3(DOUTADOUT[9]),
        .I4(DOUTADOUT[8]),
        .I5(n4[2]),
        .O(n25__0_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__0_carry_i_14__0
       (.I0(DOUTADOUT[8]),
        .I1(n4[1]),
        .I2(DOUTADOUT[9]),
        .I3(n4[0]),
        .O(n25__0_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__0_carry_i_15__0
       (.I0(n4[0]),
        .I1(DOUTADOUT[8]),
        .O(n25__0_carry_i_15__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_17__0
       (.I0(n4[5]),
        .I1(DOUTADOUT[10]),
        .O(n25__0_carry_i_17__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_18__0
       (.I0(n4[4]),
        .I1(DOUTADOUT[10]),
        .O(n25__0_carry_i_18__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_19__0
       (.I0(n4[3]),
        .I1(DOUTADOUT[10]),
        .O(n25__0_carry_i_19__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__0_carry_i_1__0
       (.I0(DOUTADOUT[10]),
        .I1(n4[4]),
        .I2(DOUTADOUT[9]),
        .I3(n4[5]),
        .I4(DOUTADOUT[8]),
        .I5(n4[6]),
        .O(n25__0_carry_i_1__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_20__0
       (.I0(n4[2]),
        .I1(DOUTADOUT[10]),
        .O(n25__0_carry_i_20__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_21
       (.I0(n4[3]),
        .I1(DOUTADOUT[8]),
        .O(n25__0_carry_i_21_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__0_carry_i_2__0
       (.I0(DOUTADOUT[10]),
        .I1(n4[3]),
        .I2(DOUTADOUT[9]),
        .I3(n4[4]),
        .I4(DOUTADOUT[8]),
        .I5(n4[5]),
        .O(n25__0_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__0_carry_i_3__0
       (.I0(DOUTADOUT[10]),
        .I1(n4[2]),
        .I2(DOUTADOUT[9]),
        .I3(n4[3]),
        .I4(DOUTADOUT[8]),
        .I5(n4[4]),
        .O(n25__0_carry_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__0_carry_i_4__0
       (.I0(DOUTADOUT[10]),
        .I1(n4[1]),
        .I2(DOUTADOUT[9]),
        .I3(n4[2]),
        .I4(DOUTADOUT[8]),
        .I5(n4[3]),
        .O(n25__0_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n25__0_carry_i_5__0
       (.I0(DOUTADOUT[9]),
        .I1(n4[2]),
        .I2(DOUTADOUT[10]),
        .I3(n4[1]),
        .I4(n4[3]),
        .I5(DOUTADOUT[8]),
        .O(n25__0_carry_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__0_carry_i_6__0
       (.I0(DOUTADOUT[9]),
        .I1(n4[1]),
        .I2(DOUTADOUT[10]),
        .I3(n4[0]),
        .O(n25__0_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__0_carry_i_7__0
       (.I0(DOUTADOUT[8]),
        .I1(n4[1]),
        .O(n25__0_carry_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n25__0_carry_i_8__0
       (.I0(n25__0_carry_i_1__0_n_0),
        .I1(DOUTADOUT[9]),
        .I2(n4[6]),
        .I3(n25__0_carry_i_17__0_n_0),
        .I4(n4[7]),
        .I5(DOUTADOUT[8]),
        .O(n25__0_carry_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__0_carry_i_9__0
       (.I0(n25__0_carry_i_2__0_n_0),
        .I1(DOUTADOUT[9]),
        .I2(n4[5]),
        .I3(n25__0_carry_i_18__0_n_0),
        .I4(n4[6]),
        .I5(DOUTADOUT[8]),
        .O(n25__0_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__27_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__27_carry_n_0,n25__27_carry_n_1,n25__27_carry_n_2,n25__27_carry_n_3,n25__27_carry_n_4,n25__27_carry_n_5,n25__27_carry_n_6,n25__27_carry_n_7}),
        .DI({n25__27_carry_i_1__0_n_0,n25__27_carry_i_2__0_n_0,n25__27_carry_i_3__0_n_0,n25__27_carry_i_4__0_n_0,n25__27_carry_i_5__0_n_0,n25__27_carry_i_6__0_n_0,n25__27_carry_i_7__0_n_0,1'b0}),
        .O({n25__27_carry_n_8,n25__27_carry_n_9,n25__27_carry_n_10,n25__27_carry_n_11,n25__27_carry_n_12,n25__27_carry_n_13,n25__27_carry_n_14,n25__27_carry_n_15}),
        .S({n25__27_carry_i_8__0_n_0,n25__27_carry_i_9__0_n_0,n25__27_carry_i_10__0_n_0,n25__27_carry_i_11__0_n_0,n25__27_carry_i_12__0_n_0,n25__27_carry_i_13__0_n_0,n25__27_carry_i_14__0_n_0,n25__27_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__27_carry__0
       (.CI(n25__27_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__27_carry__0_CO_UNCONNECTED[7:3],n25__27_carry__0_n_5,NLW_n25__27_carry__0_CO_UNCONNECTED[1],n25__27_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25__27_carry__0_i_1__0_n_0,n25__27_carry__0_i_2__0_n_0}),
        .O({NLW_n25__27_carry__0_O_UNCONNECTED[7:2],n25__27_carry__0_n_14,n25__27_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n25__27_carry__0_i_3__0_n_0,n25__27_carry__0_i_4__0_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__27_carry__0_i_1__0
       (.I0(DOUTADOUT[12]),
        .I1(n4[7]),
        .I2(DOUTADOUT[13]),
        .I3(n4[6]),
        .O(n25__27_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n25__27_carry__0_i_2__0
       (.I0(DOUTADOUT[13]),
        .I1(n4[5]),
        .I2(DOUTADOUT[12]),
        .I3(n4[6]),
        .I4(DOUTADOUT[11]),
        .I5(n4[7]),
        .O(n25__27_carry__0_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n25__27_carry__0_i_3__0
       (.I0(n4[6]),
        .I1(DOUTADOUT[12]),
        .I2(DOUTADOUT[13]),
        .I3(n4[7]),
        .O(n25__27_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n25__27_carry__0_i_4__0
       (.I0(DOUTADOUT[11]),
        .I1(n4[5]),
        .I2(n4[6]),
        .I3(DOUTADOUT[13]),
        .I4(n4[7]),
        .I5(DOUTADOUT[12]),
        .O(n25__27_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__27_carry_i_10__0
       (.I0(n25__27_carry_i_3__0_n_0),
        .I1(DOUTADOUT[12]),
        .I2(n4[4]),
        .I3(n25__27_carry_i_18__0_n_0),
        .I4(n4[5]),
        .I5(DOUTADOUT[11]),
        .O(n25__27_carry_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__27_carry_i_11__0
       (.I0(n25__27_carry_i_4__0_n_0),
        .I1(DOUTADOUT[12]),
        .I2(n4[3]),
        .I3(n25__27_carry_i_19__0_n_0),
        .I4(n4[4]),
        .I5(DOUTADOUT[11]),
        .O(n25__27_carry_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n25__27_carry_i_12__0
       (.I0(n4[2]),
        .I1(n25__27_carry_i_20__0_n_0),
        .I2(n4[1]),
        .I3(DOUTADOUT[12]),
        .I4(n4[0]),
        .I5(DOUTADOUT[13]),
        .O(n25__27_carry_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n25__27_carry_i_13__0
       (.I0(n4[0]),
        .I1(DOUTADOUT[13]),
        .I2(n4[1]),
        .I3(DOUTADOUT[12]),
        .I4(DOUTADOUT[11]),
        .I5(n4[2]),
        .O(n25__27_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__27_carry_i_14__0
       (.I0(DOUTADOUT[11]),
        .I1(n4[1]),
        .I2(DOUTADOUT[12]),
        .I3(n4[0]),
        .O(n25__27_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__27_carry_i_15__0
       (.I0(n4[0]),
        .I1(DOUTADOUT[11]),
        .O(n25__27_carry_i_15__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_16__0
       (.I0(n4[5]),
        .I1(DOUTADOUT[13]),
        .O(n25__27_carry_i_16__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_17__0
       (.I0(n4[4]),
        .I1(DOUTADOUT[13]),
        .O(n25__27_carry_i_17__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_18__0
       (.I0(n4[3]),
        .I1(DOUTADOUT[13]),
        .O(n25__27_carry_i_18__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_19__0
       (.I0(n4[2]),
        .I1(DOUTADOUT[13]),
        .O(n25__27_carry_i_19__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__27_carry_i_1__0
       (.I0(DOUTADOUT[13]),
        .I1(n4[4]),
        .I2(DOUTADOUT[12]),
        .I3(n4[5]),
        .I4(DOUTADOUT[11]),
        .I5(n4[6]),
        .O(n25__27_carry_i_1__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_20__0
       (.I0(n4[3]),
        .I1(DOUTADOUT[11]),
        .O(n25__27_carry_i_20__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__27_carry_i_2__0
       (.I0(DOUTADOUT[13]),
        .I1(n4[3]),
        .I2(DOUTADOUT[12]),
        .I3(n4[4]),
        .I4(DOUTADOUT[11]),
        .I5(n4[5]),
        .O(n25__27_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__27_carry_i_3__0
       (.I0(DOUTADOUT[13]),
        .I1(n4[2]),
        .I2(DOUTADOUT[12]),
        .I3(n4[3]),
        .I4(DOUTADOUT[11]),
        .I5(n4[4]),
        .O(n25__27_carry_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__27_carry_i_4__0
       (.I0(DOUTADOUT[13]),
        .I1(n4[1]),
        .I2(DOUTADOUT[12]),
        .I3(n4[2]),
        .I4(DOUTADOUT[11]),
        .I5(n4[3]),
        .O(n25__27_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n25__27_carry_i_5__0
       (.I0(DOUTADOUT[12]),
        .I1(n4[2]),
        .I2(DOUTADOUT[13]),
        .I3(n4[1]),
        .I4(n4[3]),
        .I5(DOUTADOUT[11]),
        .O(n25__27_carry_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__27_carry_i_6__0
       (.I0(DOUTADOUT[12]),
        .I1(n4[1]),
        .I2(DOUTADOUT[13]),
        .I3(n4[0]),
        .O(n25__27_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__27_carry_i_7__0
       (.I0(DOUTADOUT[11]),
        .I1(n4[1]),
        .O(n25__27_carry_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n25__27_carry_i_8__0
       (.I0(n25__27_carry_i_1__0_n_0),
        .I1(DOUTADOUT[12]),
        .I2(n4[6]),
        .I3(n25__27_carry_i_16__0_n_0),
        .I4(n4[7]),
        .I5(DOUTADOUT[11]),
        .O(n25__27_carry_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__27_carry_i_9__0
       (.I0(n25__27_carry_i_2__0_n_0),
        .I1(DOUTADOUT[12]),
        .I2(n4[5]),
        .I3(n25__27_carry_i_17__0_n_0),
        .I4(n4[6]),
        .I5(DOUTADOUT[11]),
        .O(n25__27_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__56_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__56_carry_n_0,n25__56_carry_n_1,n25__56_carry_n_2,n25__56_carry_n_3,n25__56_carry_n_4,n25__56_carry_n_5,n25__56_carry_n_6,n25__56_carry_n_7}),
        .DI({n25__56_carry_i_1__0_n_0,n25__56_carry_i_2__0_n_0,n25__56_carry_i_3__0_n_0,n25__56_carry_i_4__0_n_0,n25__56_carry_i_5__0_n_0,n25__56_carry_i_6__0_n_0,n25__56_carry_i_7__0_n_0,1'b0}),
        .O({n25__56_carry_n_8,n25__56_carry_n_9,n25__56_carry_n_10,n25__56_carry_n_11,n25__56_carry_n_12,n25__56_carry_n_13,n25__56_carry_n_14,n25__56_carry_n_15}),
        .S({n25__56_carry_i_8__0_n_0,n25__56_carry_i_9__0_n_0,n25__56_carry_i_10__0_n_0,n25__56_carry_i_11__0_n_0,n25__56_carry_i_12__0_n_0,n25__56_carry_i_13__0_n_0,n25__56_carry_i_14__0_n_0,n25__56_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__56_carry__0
       (.CI(n25__56_carry_n_0),
        .CI_TOP(1'b0),
        .CO(NLW_n25__56_carry__0_CO_UNCONNECTED[7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_n25__56_carry__0_O_UNCONNECTED[7:1],n25__56_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25__56_carry__0_i_1__0_n_0}));
  LUT4 #(
    .INIT(16'hE53F)) 
    n25__56_carry__0_i_1__0
       (.I0(DOUTADOUT[14]),
        .I1(n4[6]),
        .I2(DOUTADOUT[15]),
        .I3(n4[7]),
        .O(n25__56_carry__0_i_1__0_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n25__56_carry_i_10__0
       (.I0(n4[3]),
        .I1(n4[4]),
        .I2(DOUTADOUT[15]),
        .I3(n4[5]),
        .I4(DOUTADOUT[14]),
        .O(n25__56_carry_i_10__0_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n25__56_carry_i_11__0
       (.I0(n4[2]),
        .I1(n4[3]),
        .I2(DOUTADOUT[15]),
        .I3(n4[4]),
        .I4(DOUTADOUT[14]),
        .O(n25__56_carry_i_11__0_n_0));
  LUT5 #(
    .INIT(32'h9F606060)) 
    n25__56_carry_i_12__0
       (.I0(n4[1]),
        .I1(n4[2]),
        .I2(DOUTADOUT[15]),
        .I3(n4[3]),
        .I4(DOUTADOUT[14]),
        .O(n25__56_carry_i_12__0_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__56_carry_i_13__0
       (.I0(DOUTADOUT[15]),
        .I1(n4[1]),
        .I2(DOUTADOUT[14]),
        .I3(n4[2]),
        .O(n25__56_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h8777)) 
    n25__56_carry_i_14__0
       (.I0(DOUTADOUT[15]),
        .I1(n4[0]),
        .I2(DOUTADOUT[14]),
        .I3(n4[1]),
        .O(n25__56_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__56_carry_i_15__0
       (.I0(n4[0]),
        .I1(DOUTADOUT[14]),
        .O(n25__56_carry_i_15__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__56_carry_i_1__0
       (.I0(DOUTADOUT[15]),
        .I1(n4[5]),
        .I2(DOUTADOUT[14]),
        .I3(n4[6]),
        .O(n25__56_carry_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__56_carry_i_2__0
       (.I0(DOUTADOUT[15]),
        .I1(n4[4]),
        .I2(DOUTADOUT[14]),
        .I3(n4[5]),
        .O(n25__56_carry_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__56_carry_i_3__0
       (.I0(DOUTADOUT[15]),
        .I1(n4[3]),
        .I2(DOUTADOUT[14]),
        .I3(n4[4]),
        .O(n25__56_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__56_carry_i_4__0
       (.I0(DOUTADOUT[15]),
        .I1(n4[2]),
        .I2(DOUTADOUT[14]),
        .I3(n4[3]),
        .O(n25__56_carry_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n25__56_carry_i_5__0
       (.I0(n4[1]),
        .I1(DOUTADOUT[15]),
        .O(n25__56_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__56_carry_i_6__0
       (.I0(DOUTADOUT[15]),
        .I1(n4[1]),
        .O(n25__56_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n25__56_carry_i_7__0
       (.I0(n4[0]),
        .I1(DOUTADOUT[15]),
        .O(n25__56_carry_i_7__0_n_0));
  LUT5 #(
    .INIT(32'h738CC0C0)) 
    n25__56_carry_i_8__0
       (.I0(n4[5]),
        .I1(n4[6]),
        .I2(DOUTADOUT[15]),
        .I3(n4[7]),
        .I4(DOUTADOUT[14]),
        .O(n25__56_carry_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n25__56_carry_i_9__0
       (.I0(n4[4]),
        .I1(n4[5]),
        .I2(DOUTADOUT[15]),
        .I3(n4[6]),
        .I4(DOUTADOUT[14]),
        .O(n25__56_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__81_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__81_carry_n_0,n25__81_carry_n_1,n25__81_carry_n_2,n25__81_carry_n_3,n25__81_carry_n_4,n25__81_carry_n_5,n25__81_carry_n_6,n25__81_carry_n_7}),
        .DI({n25__81_carry_i_1__0_n_0,n25__81_carry_i_2__0_n_0,n25__81_carry_i_3__0_n_0,n25__81_carry_i_4__0_n_0,n25__81_carry_i_5__0_n_0,n25__81_carry_i_6__0_n_0,n25__81_carry_i_7__0_n_0,1'b0}),
        .O({n26[3:0],NLW_n25__81_carry_O_UNCONNECTED[3:0]}),
        .S({n25__81_carry_i_8__0_n_0,n25__81_carry_i_9__0_n_0,n25__81_carry_i_10__0_n_0,n25__81_carry_i_11__0_n_0,n25__81_carry_i_12__0_n_0,n25__81_carry_i_13__0_n_0,n25__81_carry_i_14__0_n_0,n25__81_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__81_carry__0
       (.CI(n25__81_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__81_carry__0_CO_UNCONNECTED[7:3],n25__81_carry__0_n_5,n25__81_carry__0_n_6,n25__81_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n25__81_carry__0_i_1__0_n_0,n25__81_carry__0_i_2__0_n_0,n25__81_carry__0_i_3__0_n_0}),
        .O({NLW_n25__81_carry__0_O_UNCONNECTED[7:4],n26[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n25__81_carry__0_i_4__0_n_0,n25__81_carry__0_i_5__0_n_0,n25__81_carry__0_i_6__0_n_0,n25__81_carry__0_i_7__0_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry__0_i_1__0
       (.I0(n25__27_carry__0_n_14),
        .I1(n25__56_carry_n_9),
        .O(n25__81_carry__0_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry__0_i_2__0
       (.I0(n25__27_carry__0_n_15),
        .I1(n25__56_carry_n_10),
        .O(n25__81_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry__0_i_3__0
       (.I0(n25__56_carry_n_11),
        .I1(n25__27_carry_n_8),
        .I2(n25__0_carry__0_n_5),
        .O(n25__81_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n25__81_carry__0_i_4__0
       (.I0(n25__27_carry__0_n_5),
        .I1(n25__56_carry_n_8),
        .I2(n25__56_carry__0_n_15),
        .O(n25__81_carry__0_i_4__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__81_carry__0_i_5__0
       (.I0(n25__27_carry__0_n_14),
        .I1(n25__56_carry_n_9),
        .I2(n25__56_carry_n_8),
        .I3(n25__27_carry__0_n_5),
        .O(n25__81_carry__0_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__81_carry__0_i_6__0
       (.I0(n25__27_carry__0_n_15),
        .I1(n25__56_carry_n_10),
        .I2(n25__56_carry_n_9),
        .I3(n25__27_carry__0_n_14),
        .O(n25__81_carry__0_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n25__81_carry__0_i_7__0
       (.I0(n25__0_carry__0_n_5),
        .I1(n25__27_carry_n_8),
        .I2(n25__56_carry_n_11),
        .I3(n25__56_carry_n_10),
        .I4(n25__27_carry__0_n_15),
        .O(n25__81_carry__0_i_7__0_n_0));
  (* HLUTNM = "lutpair2" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_10__0
       (.I0(n25__56_carry_n_13),
        .I1(n25__27_carry_n_10),
        .I2(n25__0_carry__0_n_15),
        .I3(n25__81_carry_i_3__0_n_0),
        .O(n25__81_carry_i_10__0_n_0));
  (* HLUTNM = "lutpair1" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_11__0
       (.I0(n25__56_carry_n_14),
        .I1(n25__27_carry_n_11),
        .I2(n25__0_carry_n_8),
        .I3(n25__81_carry_i_4__0_n_0),
        .O(n25__81_carry_i_11__0_n_0));
  (* HLUTNM = "lutpair0" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_12__0
       (.I0(n25__56_carry_n_15),
        .I1(n25__27_carry_n_12),
        .I2(n25__0_carry_n_9),
        .I3(n25__81_carry_i_5__0_n_0),
        .O(n25__81_carry_i_12__0_n_0));
  (* HLUTNM = "lutpair80" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n25__81_carry_i_13__0
       (.I0(n25__27_carry_n_13),
        .I1(n25__0_carry_n_10),
        .I2(n25__0_carry_n_11),
        .I3(n25__27_carry_n_14),
        .O(n25__81_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__81_carry_i_14__0
       (.I0(n25__0_carry_n_12),
        .I1(n25__27_carry_n_15),
        .I2(n25__27_carry_n_14),
        .I3(n25__0_carry_n_11),
        .O(n25__81_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n25__81_carry_i_15__0
       (.I0(n25__0_carry_n_12),
        .I1(n25__27_carry_n_15),
        .O(n25__81_carry_i_15__0_n_0));
  (* HLUTNM = "lutpair3" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry_i_1__0
       (.I0(n25__56_carry_n_12),
        .I1(n25__27_carry_n_9),
        .I2(n25__0_carry__0_n_14),
        .O(n25__81_carry_i_1__0_n_0));
  (* HLUTNM = "lutpair2" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry_i_2__0
       (.I0(n25__56_carry_n_13),
        .I1(n25__27_carry_n_10),
        .I2(n25__0_carry__0_n_15),
        .O(n25__81_carry_i_2__0_n_0));
  (* HLUTNM = "lutpair1" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry_i_3__0
       (.I0(n25__56_carry_n_14),
        .I1(n25__27_carry_n_11),
        .I2(n25__0_carry_n_8),
        .O(n25__81_carry_i_3__0_n_0));
  (* HLUTNM = "lutpair0" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry_i_4__0
       (.I0(n25__56_carry_n_15),
        .I1(n25__27_carry_n_12),
        .I2(n25__0_carry_n_9),
        .O(n25__81_carry_i_4__0_n_0));
  (* HLUTNM = "lutpair80" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry_i_5__0
       (.I0(n25__27_carry_n_13),
        .I1(n25__0_carry_n_10),
        .O(n25__81_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry_i_6__0
       (.I0(n25__0_carry_n_11),
        .I1(n25__27_carry_n_14),
        .O(n25__81_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry_i_7__0
       (.I0(n25__0_carry_n_12),
        .I1(n25__27_carry_n_15),
        .O(n25__81_carry_i_7__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_8__0
       (.I0(n25__81_carry_i_1__0_n_0),
        .I1(n25__27_carry_n_8),
        .I2(n25__56_carry_n_11),
        .I3(n25__0_carry__0_n_5),
        .O(n25__81_carry_i_8__0_n_0));
  (* HLUTNM = "lutpair3" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_9__0
       (.I0(n25__56_carry_n_12),
        .I1(n25__27_carry_n_9),
        .I2(n25__0_carry__0_n_14),
        .I3(n25__81_carry_i_2__0_n_0),
        .O(n25__81_carry_i_9__0_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[0]),
        .Q(n27[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[1]),
        .Q(n27[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[2]),
        .Q(n27[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[3]),
        .Q(n27[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[4]),
        .Q(n27[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[5]),
        .Q(n27[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[6]),
        .Q(n27[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[7]),
        .Q(n27[7]),
        .R(rst_i));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_2 
       (.I0(n24[7]),
        .I1(n27[7]),
        .O(\n29[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_3 
       (.I0(n24[6]),
        .I1(n27[6]),
        .O(\n29[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_4 
       (.I0(n24[5]),
        .I1(n27[5]),
        .O(\n29[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_5 
       (.I0(n24[4]),
        .I1(n27[4]),
        .O(\n29[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_6 
       (.I0(n24[3]),
        .I1(n27[3]),
        .O(\n29[7]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_7 
       (.I0(n24[2]),
        .I1(n27[2]),
        .O(\n29[7]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_8 
       (.I0(n24[1]),
        .I1(n27[1]),
        .O(\n29[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_9 
       (.I0(n24[0]),
        .I1(n27[0]),
        .O(\n29[7]_i_9_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[0]),
        .Q(n29[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[1]),
        .Q(n29[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[2]),
        .Q(n29[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[3]),
        .Q(n29[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[4]),
        .Q(n29[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[5]),
        .Q(n29[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[6]),
        .Q(n29[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[7]),
        .Q(n29[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n29_reg[7]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\NLW_n29_reg[7]_i_1_CO_UNCONNECTED [7],\n29_reg[7]_i_1_n_1 ,\n29_reg[7]_i_1_n_2 ,\n29_reg[7]_i_1_n_3 ,\n29_reg[7]_i_1_n_4 ,\n29_reg[7]_i_1_n_5 ,\n29_reg[7]_i_1_n_6 ,\n29_reg[7]_i_1_n_7 }),
        .DI({1'b0,n24[6:0]}),
        .O(n28),
        .S({\n29[7]_i_2_n_0 ,\n29[7]_i_3_n_0 ,\n29[7]_i_4_n_0 ,\n29[7]_i_5_n_0 ,\n29[7]_i_6_n_0 ,\n29[7]_i_7_n_0 ,\n29[7]_i_8_n_0 ,\n29[7]_i_9_n_0 }));
  LUT2 #(
    .INIT(4'h6)) 
    \n33[0]_i_1__0 
       (.I0(n29[0]),
        .I1(n10[0]),
        .O(n31[0]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[10]_i_1__0 
       (.I0(n21[2]),
        .I1(\n8_reg_n_0_[2] ),
        .I2(\n8_reg_n_0_[1] ),
        .I3(n21[1]),
        .I4(\n8_reg_n_0_[0] ),
        .I5(n21[0]),
        .O(\n33[10]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[11]_i_1__0 
       (.I0(n21[3]),
        .I1(\n8_reg_n_0_[3] ),
        .I2(\n33[12]_i_2__0_n_0 ),
        .O(\n33[11]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[12]_i_1__0 
       (.I0(n21[4]),
        .I1(\n8_reg_n_0_[4] ),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[3]),
        .I4(\n33[12]_i_2__0_n_0 ),
        .O(\n33[12]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[12]_i_2__0 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n33[12]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[13]_i_1__0 
       (.I0(n21[5]),
        .I1(\n8_reg_n_0_[5] ),
        .I2(\n33[14]_i_2__0_n_0 ),
        .O(\n33[13]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[14]_i_1__0 
       (.I0(n21[6]),
        .I1(\n8_reg_n_0_[6] ),
        .I2(\n8_reg_n_0_[5] ),
        .I3(n21[5]),
        .I4(\n33[14]_i_2__0_n_0 ),
        .O(\n33[14]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[14]_i_2__0 
       (.I0(\n33[12]_i_2__0_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n33[14]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[15]_i_1__0 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n33[15]_i_2__0_n_0 ),
        .O(n30[7]));
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[15]_i_2__0 
       (.I0(\n33[14]_i_2__0_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n33[15]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[1]_i_1__0 
       (.I0(n29[1]),
        .I1(n10[1]),
        .I2(n10[0]),
        .I3(n29[0]),
        .O(n31[1]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[2]_i_1__0 
       (.I0(n29[2]),
        .I1(n10[2]),
        .I2(n10[1]),
        .I3(n29[1]),
        .I4(n10[0]),
        .I5(n29[0]),
        .O(\n33[2]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[3]_i_1__0 
       (.I0(n29[3]),
        .I1(n10[3]),
        .I2(\n33[4]_i_2__0_n_0 ),
        .O(\n33[3]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[4]_i_1__0 
       (.I0(n29[4]),
        .I1(n10[4]),
        .I2(n10[3]),
        .I3(n29[3]),
        .I4(\n33[4]_i_2__0_n_0 ),
        .O(\n33[4]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[4]_i_2__0 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n33[4]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[5]_i_1__0 
       (.I0(n29[5]),
        .I1(n10[5]),
        .I2(\n33[6]_i_2__0_n_0 ),
        .O(\n33[5]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[6]_i_1__0 
       (.I0(n29[6]),
        .I1(n10[6]),
        .I2(n10[5]),
        .I3(n29[5]),
        .I4(\n33[6]_i_2__0_n_0 ),
        .O(\n33[6]_i_1__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[6]_i_2__0 
       (.I0(\n33[4]_i_2__0_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n33[6]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[7]_i_1__0 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n33[7]_i_2__0_n_0 ),
        .O(n31[7]));
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[7]_i_2__0 
       (.I0(\n33[6]_i_2__0_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n33[7]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n33[8]_i_1 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .O(n30[0]));
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[9]_i_1__0 
       (.I0(n21[1]),
        .I1(\n8_reg_n_0_[1] ),
        .I2(\n8_reg_n_0_[0] ),
        .I3(n21[0]),
        .O(\n33[9]_i_1__0_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[0]),
        .Q(i1[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[10]_i_1__0_n_0 ),
        .Q(i1[24]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[11]_i_1__0_n_0 ),
        .Q(i1[25]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[12]_i_1__0_n_0 ),
        .Q(i1[26]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[13]_i_1__0_n_0 ),
        .Q(i1[27]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[14]_i_1__0_n_0 ),
        .Q(i1[28]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n30[7]),
        .Q(i1[29]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[1]),
        .Q(i1[15]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[2]_i_1__0_n_0 ),
        .Q(i1[16]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[3]_i_1__0_n_0 ),
        .Q(i1[17]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[4]_i_1__0_n_0 ),
        .Q(i1[18]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[5]_i_1__0_n_0 ),
        .Q(i1[19]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[6]_i_1__0_n_0 ),
        .Q(i1[20]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[7]),
        .Q(i1[21]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n30[0]),
        .Q(i1[22]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[9]_i_1__0_n_0 ),
        .Q(i1[23]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[10]_i_1__0 
       (.I0(\n8_reg_n_0_[1] ),
        .I1(n21[1]),
        .I2(n21[0]),
        .I3(\n8_reg_n_0_[0] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(n341_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[11]_i_1__0 
       (.I0(\n37[12]_i_2__0_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .O(n341_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[12]_i_1__0 
       (.I0(\n8_reg_n_0_[3] ),
        .I1(n21[3]),
        .I2(\n37[12]_i_2__0_n_0 ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(n341_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[12]_i_2__0 
       (.I0(\n8_reg_n_0_[0] ),
        .I1(n21[0]),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n37[12]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[13]_i_1__0 
       (.I0(\n37[14]_i_2__0_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(n341_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[14]_i_1__0 
       (.I0(\n8_reg_n_0_[5] ),
        .I1(n21[5]),
        .I2(\n37[14]_i_2__0_n_0 ),
        .I3(n21[6]),
        .I4(\n8_reg_n_0_[6] ),
        .O(n341_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[14]_i_2__0 
       (.I0(\n37[12]_i_2__0_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n37[14]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[15]_i_1__0 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n37[15]_i_2__0_n_0 ),
        .O(n341_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[15]_i_2__0 
       (.I0(\n37[14]_i_2__0_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n37[15]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[1]_i_1__0 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .O(n350_out[1]));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[2]_i_1__0 
       (.I0(n10[1]),
        .I1(n29[1]),
        .I2(n29[0]),
        .I3(n10[0]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(n350_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[3]_i_1__0 
       (.I0(\n37[4]_i_2__0_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .O(n350_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[4]_i_1__0 
       (.I0(n10[3]),
        .I1(n29[3]),
        .I2(\n37[4]_i_2__0_n_0 ),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(n350_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[4]_i_2__0 
       (.I0(n10[0]),
        .I1(n29[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n37[4]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[5]_i_1__0 
       (.I0(\n37[6]_i_2__0_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(n350_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[6]_i_1__0 
       (.I0(n10[5]),
        .I1(n29[5]),
        .I2(\n37[6]_i_2__0_n_0 ),
        .I3(n29[6]),
        .I4(n10[6]),
        .O(n350_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[6]_i_2__0 
       (.I0(\n37[4]_i_2__0_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n37[6]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[7]_i_1__0 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n37[7]_i_2__0_n_0 ),
        .O(n350_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[7]_i_2__0 
       (.I0(\n37[6]_i_2__0_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n37[7]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[9]_i_1__0 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .O(n341_out[1]));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[2]),
        .Q(i1[9]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[3]),
        .Q(i1[10]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[4]),
        .Q(i1[11]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[5]),
        .Q(i1[12]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[6]),
        .Q(i1[13]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[7]),
        .Q(i1[14]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[1]),
        .Q(i1[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[2]),
        .Q(i1[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[3]),
        .Q(i1[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[4]),
        .Q(i1[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[5]),
        .Q(i1[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[6]),
        .Q(i1[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[7]),
        .Q(i1[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[1]),
        .Q(i1[8]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[0]),
        .Q(n4[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[1]),
        .Q(n4[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[2]),
        .Q(n4[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[3]),
        .Q(n4[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[4]),
        .Q(n4[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[5]),
        .Q(n4[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[6]),
        .Q(n4[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s3_3[7]),
        .Q(n4[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[0]),
        .Q(\n7_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[1]),
        .Q(\n7_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[2]),
        .Q(\n7_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[3]),
        .Q(\n7_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[4]),
        .Q(\n7_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[5]),
        .Q(\n7_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[6]),
        .Q(\n7_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[7]),
        .Q(\n7_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[0] ),
        .Q(\n8_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[1] ),
        .Q(\n8_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[2] ),
        .Q(\n8_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[3] ),
        .Q(\n8_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[4] ),
        .Q(\n8_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[5] ),
        .Q(\n8_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[6] ),
        .Q(\n8_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[7] ),
        .Q(\n8_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[0] ),
        .Q(\n9_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[1] ),
        .Q(\n9_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[2] ),
        .Q(\n9_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[3] ),
        .Q(\n9_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[4] ),
        .Q(\n9_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[5] ),
        .Q(\n9_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[6] ),
        .Q(\n9_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[7] ),
        .Q(\n9_reg_n_0_[7] ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_19" *) 
module switch_elements_cf_fft_512_8_19
   (p_6_out,
    inf4_s,
    enable_s,
    rst_i,
    enable_i,
    clk_i,
    s2_3,
    D);
  output [31:0]p_6_out;
  output [31:0]inf4_s;
  input [31:0]enable_s;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]s2_3;
  input [15:0]D;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [31:0]enable_s;
  wire [0:0]i8;
  wire [31:0]inf4_s;
  wire n12;
  wire [15:0]n33;
  wire [15:1]n37;
  wire n4;
  wire [31:0]p_6_out;
  wire rst_i;
  wire [15:0]s2_3;

  switch_elements_cf_fft_512_8_20 s25
       (.D(D),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .rst_i(rst_i),
        .s2_3(s2_3));
  switch_elements_cf_fft_512_8_31_19 s26
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i8(i8),
        .n4(n4),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_27_20 s27
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .enable_s({enable_s[31:28],enable_s[15:12],enable_s[7:0]}),
        .i1({n33[15:9],n33[7:0],n37}),
        .i8(i8),
        .inf4_s(inf4_s[31:16]),
        .\info_o_reg[27] (inf4_s[7:0]),
        .n12(n12),
        .p_6_out(p_6_out[27:16]),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_26_21 s28
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .enable_s(enable_s[27:0]),
        .i1({n33[15:9],n37[8],n33[7:0],n37[15:9],n37[7:1]}),
        .i8(i8),
        .inf4_s({inf4_s[31:28],inf4_s[19:16]}),
        .n12(n12),
        .\n12_reg[0]_0 (inf4_s[15:0]),
        .n4(n4),
        .p_6_out({p_6_out[31:28],p_6_out[15:0]}),
        .rst_i(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_2" *) 
module switch_elements_cf_fft_512_8_2
   (\n5_reg[0] ,
    \n5_reg[0]_0 ,
    \n5_reg[0]_1 ,
    rst_i,
    enable_i,
    clk_i,
    i2,
    n22);
  output [15:0]\n5_reg[0] ;
  output [7:0]\n5_reg[0]_0 ;
  output [7:0]\n5_reg[0]_1 ;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [31:0]i2;
  input n22;

  wire clk_i;
  wire [0:0]enable_i;
  wire [31:0]i2;
  wire [0:0]i8;
  wire n22;
  wire n4;
  wire [15:0]\n5_reg[0] ;
  wire [7:0]\n5_reg[0]_0 ;
  wire [7:0]\n5_reg[0]_1 ;
  wire rst_i;

  switch_elements_cf_fft_512_8_31 s13
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i8(i8),
        .n4(n4),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_4 s14
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i2(i2),
        .i8(i8),
        .n22(n22),
        .\n5_reg[0] (\n5_reg[0]_0 ),
        .\n5_reg[0]_0 (\n5_reg[0]_1 ),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_3 s15
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i2(i2),
        .i8(i8),
        .\n1_reg[15] (n22),
        .n4(n4),
        .\n5_reg[0] (\n5_reg[0] ),
        .rst_i(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_20" *) 
module switch_elements_cf_fft_512_8_20
   (i1,
    clk_i,
    enable_i,
    rst_i,
    s2_3,
    D);
  output [29:0]i1;
  input clk_i;
  input [0:0]enable_i;
  input rst_i;
  input [15:0]s2_3;
  input [15:0]D;

  wire [7:0]B;
  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [7:0]n10;
  wire n11_reg_n_40;
  wire n11_reg_n_41;
  wire n11_reg_n_42;
  wire n11_reg_n_43;
  wire n11_reg_n_44;
  wire n11_reg_n_45;
  wire n11_reg_n_46;
  wire n11_reg_n_47;
  wire n14__0_carry__0_i_1_n_0;
  wire n14__0_carry__0_i_2_n_0;
  wire n14__0_carry__0_i_3_n_0;
  wire n14__0_carry__0_i_4_n_0;
  wire n14__0_carry__0_n_14;
  wire n14__0_carry__0_n_15;
  wire n14__0_carry__0_n_5;
  wire n14__0_carry__0_n_7;
  wire n14__0_carry_i_10_n_0;
  wire n14__0_carry_i_11_n_0;
  wire n14__0_carry_i_12_n_0;
  wire n14__0_carry_i_13_n_0;
  wire n14__0_carry_i_14_n_0;
  wire n14__0_carry_i_15_n_0;
  wire n14__0_carry_i_16_n_0;
  wire n14__0_carry_i_17_n_0;
  wire n14__0_carry_i_18_n_0;
  wire n14__0_carry_i_19_n_0;
  wire n14__0_carry_i_1_n_0;
  wire n14__0_carry_i_20_n_0;
  wire n14__0_carry_i_2_n_0;
  wire n14__0_carry_i_3_n_0;
  wire n14__0_carry_i_4_n_0;
  wire n14__0_carry_i_5_n_0;
  wire n14__0_carry_i_6_n_0;
  wire n14__0_carry_i_7_n_0;
  wire n14__0_carry_i_8_n_0;
  wire n14__0_carry_i_9_n_0;
  wire n14__0_carry_n_0;
  wire n14__0_carry_n_1;
  wire n14__0_carry_n_10;
  wire n14__0_carry_n_11;
  wire n14__0_carry_n_12;
  wire n14__0_carry_n_2;
  wire n14__0_carry_n_3;
  wire n14__0_carry_n_4;
  wire n14__0_carry_n_5;
  wire n14__0_carry_n_6;
  wire n14__0_carry_n_7;
  wire n14__0_carry_n_8;
  wire n14__0_carry_n_9;
  wire n14__27_carry__0_i_1_n_0;
  wire n14__27_carry__0_i_2_n_0;
  wire n14__27_carry__0_i_3_n_0;
  wire n14__27_carry__0_i_4_n_0;
  wire n14__27_carry__0_n_14;
  wire n14__27_carry__0_n_15;
  wire n14__27_carry__0_n_5;
  wire n14__27_carry__0_n_7;
  wire n14__27_carry_i_10_n_0;
  wire n14__27_carry_i_11_n_0;
  wire n14__27_carry_i_12_n_0;
  wire n14__27_carry_i_13_n_0;
  wire n14__27_carry_i_14_n_0;
  wire n14__27_carry_i_15_n_0;
  wire n14__27_carry_i_16_n_0;
  wire n14__27_carry_i_17_n_0;
  wire n14__27_carry_i_18_n_0;
  wire n14__27_carry_i_19_n_0;
  wire n14__27_carry_i_1_n_0;
  wire n14__27_carry_i_20_n_0;
  wire n14__27_carry_i_2_n_0;
  wire n14__27_carry_i_3_n_0;
  wire n14__27_carry_i_4_n_0;
  wire n14__27_carry_i_5_n_0;
  wire n14__27_carry_i_6_n_0;
  wire n14__27_carry_i_7_n_0;
  wire n14__27_carry_i_8_n_0;
  wire n14__27_carry_i_9_n_0;
  wire n14__27_carry_n_0;
  wire n14__27_carry_n_1;
  wire n14__27_carry_n_10;
  wire n14__27_carry_n_11;
  wire n14__27_carry_n_12;
  wire n14__27_carry_n_13;
  wire n14__27_carry_n_14;
  wire n14__27_carry_n_15;
  wire n14__27_carry_n_2;
  wire n14__27_carry_n_3;
  wire n14__27_carry_n_4;
  wire n14__27_carry_n_5;
  wire n14__27_carry_n_6;
  wire n14__27_carry_n_7;
  wire n14__27_carry_n_8;
  wire n14__27_carry_n_9;
  wire n14__56_carry__0_i_1_n_0;
  wire n14__56_carry__0_n_15;
  wire n14__56_carry_i_10_n_0;
  wire n14__56_carry_i_11_n_0;
  wire n14__56_carry_i_12_n_0;
  wire n14__56_carry_i_13_n_0;
  wire n14__56_carry_i_14_n_0;
  wire n14__56_carry_i_15_n_0;
  wire n14__56_carry_i_1_n_0;
  wire n14__56_carry_i_2_n_0;
  wire n14__56_carry_i_3_n_0;
  wire n14__56_carry_i_4_n_0;
  wire n14__56_carry_i_5_n_0;
  wire n14__56_carry_i_6_n_0;
  wire n14__56_carry_i_7_n_0;
  wire n14__56_carry_i_8_n_0;
  wire n14__56_carry_i_9_n_0;
  wire n14__56_carry_n_0;
  wire n14__56_carry_n_1;
  wire n14__56_carry_n_10;
  wire n14__56_carry_n_11;
  wire n14__56_carry_n_12;
  wire n14__56_carry_n_13;
  wire n14__56_carry_n_14;
  wire n14__56_carry_n_15;
  wire n14__56_carry_n_2;
  wire n14__56_carry_n_3;
  wire n14__56_carry_n_4;
  wire n14__56_carry_n_5;
  wire n14__56_carry_n_6;
  wire n14__56_carry_n_7;
  wire n14__56_carry_n_8;
  wire n14__56_carry_n_9;
  wire n14__81_carry__0_i_1_n_0;
  wire n14__81_carry__0_i_2_n_0;
  wire n14__81_carry__0_i_3_n_0;
  wire n14__81_carry__0_i_4_n_0;
  wire n14__81_carry__0_i_5_n_0;
  wire n14__81_carry__0_i_6_n_0;
  wire n14__81_carry__0_i_7_n_0;
  wire n14__81_carry__0_n_5;
  wire n14__81_carry__0_n_6;
  wire n14__81_carry__0_n_7;
  wire n14__81_carry_i_10_n_0;
  wire n14__81_carry_i_11_n_0;
  wire n14__81_carry_i_12_n_0;
  wire n14__81_carry_i_13_n_0;
  wire n14__81_carry_i_14_n_0;
  wire n14__81_carry_i_15_n_0;
  wire n14__81_carry_i_1_n_0;
  wire n14__81_carry_i_2_n_0;
  wire n14__81_carry_i_3_n_0;
  wire n14__81_carry_i_4_n_0;
  wire n14__81_carry_i_5_n_0;
  wire n14__81_carry_i_6_n_0;
  wire n14__81_carry_i_7_n_0;
  wire n14__81_carry_i_8_n_0;
  wire n14__81_carry_i_9_n_0;
  wire n14__81_carry_n_0;
  wire n14__81_carry_n_1;
  wire n14__81_carry_n_2;
  wire n14__81_carry_n_3;
  wire n14__81_carry_n_4;
  wire n14__81_carry_n_5;
  wire n14__81_carry_n_6;
  wire n14__81_carry_n_7;
  wire [7:0]n15;
  wire \n16_reg_n_0_[0] ;
  wire \n16_reg_n_0_[1] ;
  wire \n16_reg_n_0_[2] ;
  wire \n16_reg_n_0_[3] ;
  wire \n16_reg_n_0_[4] ;
  wire \n16_reg_n_0_[5] ;
  wire \n16_reg_n_0_[6] ;
  wire \n16_reg_n_0_[7] ;
  wire [14:7]n17;
  wire n17__0_carry__0_i_1_n_0;
  wire n17__0_carry__0_i_2_n_0;
  wire n17__0_carry__0_i_3_n_0;
  wire n17__0_carry__0_i_4_n_0;
  wire n17__0_carry__0_n_14;
  wire n17__0_carry__0_n_15;
  wire n17__0_carry__0_n_5;
  wire n17__0_carry__0_n_7;
  wire n17__0_carry_i_10_n_0;
  wire n17__0_carry_i_11_n_0;
  wire n17__0_carry_i_12_n_0;
  wire n17__0_carry_i_13_n_0;
  wire n17__0_carry_i_14_n_0;
  wire n17__0_carry_i_15_n_0;
  wire n17__0_carry_i_16_n_0;
  wire n17__0_carry_i_17_n_0;
  wire n17__0_carry_i_18_n_0;
  wire n17__0_carry_i_19_n_0;
  wire n17__0_carry_i_1_n_0;
  wire n17__0_carry_i_20_n_0;
  wire n17__0_carry_i_2_n_0;
  wire n17__0_carry_i_3_n_0;
  wire n17__0_carry_i_4_n_0;
  wire n17__0_carry_i_5_n_0;
  wire n17__0_carry_i_6_n_0;
  wire n17__0_carry_i_7_n_0;
  wire n17__0_carry_i_8_n_0;
  wire n17__0_carry_i_9_n_0;
  wire n17__0_carry_n_0;
  wire n17__0_carry_n_1;
  wire n17__0_carry_n_10;
  wire n17__0_carry_n_11;
  wire n17__0_carry_n_12;
  wire n17__0_carry_n_2;
  wire n17__0_carry_n_3;
  wire n17__0_carry_n_4;
  wire n17__0_carry_n_5;
  wire n17__0_carry_n_6;
  wire n17__0_carry_n_7;
  wire n17__0_carry_n_8;
  wire n17__0_carry_n_9;
  wire n17__27_carry__0_i_1_n_0;
  wire n17__27_carry__0_i_2_n_0;
  wire n17__27_carry__0_i_3_n_0;
  wire n17__27_carry__0_i_4_n_0;
  wire n17__27_carry__0_n_14;
  wire n17__27_carry__0_n_15;
  wire n17__27_carry__0_n_5;
  wire n17__27_carry__0_n_7;
  wire n17__27_carry_i_10_n_0;
  wire n17__27_carry_i_11_n_0;
  wire n17__27_carry_i_12_n_0;
  wire n17__27_carry_i_13_n_0;
  wire n17__27_carry_i_14_n_0;
  wire n17__27_carry_i_15_n_0;
  wire n17__27_carry_i_16_n_0;
  wire n17__27_carry_i_17_n_0;
  wire n17__27_carry_i_18_n_0;
  wire n17__27_carry_i_19_n_0;
  wire n17__27_carry_i_1_n_0;
  wire n17__27_carry_i_20_n_0;
  wire n17__27_carry_i_2_n_0;
  wire n17__27_carry_i_3_n_0;
  wire n17__27_carry_i_4_n_0;
  wire n17__27_carry_i_5_n_0;
  wire n17__27_carry_i_6_n_0;
  wire n17__27_carry_i_7_n_0;
  wire n17__27_carry_i_8_n_0;
  wire n17__27_carry_i_9_n_0;
  wire n17__27_carry_n_0;
  wire n17__27_carry_n_1;
  wire n17__27_carry_n_10;
  wire n17__27_carry_n_11;
  wire n17__27_carry_n_12;
  wire n17__27_carry_n_13;
  wire n17__27_carry_n_14;
  wire n17__27_carry_n_15;
  wire n17__27_carry_n_2;
  wire n17__27_carry_n_3;
  wire n17__27_carry_n_4;
  wire n17__27_carry_n_5;
  wire n17__27_carry_n_6;
  wire n17__27_carry_n_7;
  wire n17__27_carry_n_8;
  wire n17__27_carry_n_9;
  wire n17__56_carry__0_i_1_n_0;
  wire n17__56_carry__0_n_15;
  wire n17__56_carry_i_10_n_0;
  wire n17__56_carry_i_11_n_0;
  wire n17__56_carry_i_12_n_0;
  wire n17__56_carry_i_13_n_0;
  wire n17__56_carry_i_14_n_0;
  wire n17__56_carry_i_15_n_0;
  wire n17__56_carry_i_1_n_0;
  wire n17__56_carry_i_2_n_0;
  wire n17__56_carry_i_3_n_0;
  wire n17__56_carry_i_4_n_0;
  wire n17__56_carry_i_5_n_0;
  wire n17__56_carry_i_6_n_0;
  wire n17__56_carry_i_7_n_0;
  wire n17__56_carry_i_8_n_0;
  wire n17__56_carry_i_9_n_0;
  wire n17__56_carry_n_0;
  wire n17__56_carry_n_1;
  wire n17__56_carry_n_10;
  wire n17__56_carry_n_11;
  wire n17__56_carry_n_12;
  wire n17__56_carry_n_13;
  wire n17__56_carry_n_14;
  wire n17__56_carry_n_15;
  wire n17__56_carry_n_2;
  wire n17__56_carry_n_3;
  wire n17__56_carry_n_4;
  wire n17__56_carry_n_5;
  wire n17__56_carry_n_6;
  wire n17__56_carry_n_7;
  wire n17__56_carry_n_8;
  wire n17__56_carry_n_9;
  wire n17__81_carry__0_i_1_n_0;
  wire n17__81_carry__0_i_2_n_0;
  wire n17__81_carry__0_i_3_n_0;
  wire n17__81_carry__0_i_4_n_0;
  wire n17__81_carry__0_i_5_n_0;
  wire n17__81_carry__0_i_6_n_0;
  wire n17__81_carry__0_i_7_n_0;
  wire n17__81_carry__0_n_5;
  wire n17__81_carry__0_n_6;
  wire n17__81_carry__0_n_7;
  wire n17__81_carry_i_10_n_0;
  wire n17__81_carry_i_11_n_0;
  wire n17__81_carry_i_12_n_0;
  wire n17__81_carry_i_13_n_0;
  wire n17__81_carry_i_14_n_0;
  wire n17__81_carry_i_15_n_0;
  wire n17__81_carry_i_1_n_0;
  wire n17__81_carry_i_2_n_0;
  wire n17__81_carry_i_3_n_0;
  wire n17__81_carry_i_4_n_0;
  wire n17__81_carry_i_5_n_0;
  wire n17__81_carry_i_6_n_0;
  wire n17__81_carry_i_7_n_0;
  wire n17__81_carry_i_8_n_0;
  wire n17__81_carry_i_9_n_0;
  wire n17__81_carry_n_0;
  wire n17__81_carry_n_1;
  wire n17__81_carry_n_2;
  wire n17__81_carry_n_3;
  wire n17__81_carry_n_4;
  wire n17__81_carry_n_5;
  wire n17__81_carry_n_6;
  wire n17__81_carry_n_7;
  wire n19_reg__0_n_0;
  wire n19_reg__1_n_0;
  wire n19_reg__2_n_0;
  wire n19_reg__3_n_0;
  wire n19_reg__4_n_0;
  wire n19_reg__5_n_0;
  wire n19_reg__6_n_0;
  wire n19_reg_n_0;
  wire \n1_reg_n_0_[0] ;
  wire \n1_reg_n_0_[1] ;
  wire \n1_reg_n_0_[2] ;
  wire \n1_reg_n_0_[3] ;
  wire \n1_reg_n_0_[4] ;
  wire \n1_reg_n_0_[5] ;
  wire \n1_reg_n_0_[6] ;
  wire \n1_reg_n_0_[7] ;
  wire [7:0]n2;
  wire [7:0]n202_out;
  wire n20_carry_i_1__0_n_0;
  wire n20_carry_i_2__0_n_0;
  wire n20_carry_i_3__0_n_0;
  wire n20_carry_i_4__0_n_0;
  wire n20_carry_i_5__0_n_0;
  wire n20_carry_i_6__0_n_0;
  wire n20_carry_i_7__0_n_0;
  wire n20_carry_i_8__0_n_0;
  wire n20_carry_n_1;
  wire n20_carry_n_2;
  wire n20_carry_n_3;
  wire n20_carry_n_4;
  wire n20_carry_n_5;
  wire n20_carry_n_6;
  wire n20_carry_n_7;
  wire [7:0]n21;
  wire n22__0_carry__0_i_1_n_0;
  wire n22__0_carry__0_i_2_n_0;
  wire n22__0_carry__0_i_3_n_0;
  wire n22__0_carry__0_i_4_n_0;
  wire n22__0_carry__0_n_14;
  wire n22__0_carry__0_n_15;
  wire n22__0_carry__0_n_5;
  wire n22__0_carry__0_n_7;
  wire n22__0_carry_i_10_n_0;
  wire n22__0_carry_i_11_n_0;
  wire n22__0_carry_i_12_n_0;
  wire n22__0_carry_i_13_n_0;
  wire n22__0_carry_i_14_n_0;
  wire n22__0_carry_i_15_n_0;
  wire n22__0_carry_i_16_n_0;
  wire n22__0_carry_i_17_n_0;
  wire n22__0_carry_i_18_n_0;
  wire n22__0_carry_i_19_n_0;
  wire n22__0_carry_i_1_n_0;
  wire n22__0_carry_i_20_n_0;
  wire n22__0_carry_i_2_n_0;
  wire n22__0_carry_i_3_n_0;
  wire n22__0_carry_i_4_n_0;
  wire n22__0_carry_i_5_n_0;
  wire n22__0_carry_i_6_n_0;
  wire n22__0_carry_i_7_n_0;
  wire n22__0_carry_i_8_n_0;
  wire n22__0_carry_i_9_n_0;
  wire n22__0_carry_n_0;
  wire n22__0_carry_n_1;
  wire n22__0_carry_n_10;
  wire n22__0_carry_n_11;
  wire n22__0_carry_n_12;
  wire n22__0_carry_n_2;
  wire n22__0_carry_n_3;
  wire n22__0_carry_n_4;
  wire n22__0_carry_n_5;
  wire n22__0_carry_n_6;
  wire n22__0_carry_n_7;
  wire n22__0_carry_n_8;
  wire n22__0_carry_n_9;
  wire n22__0_n_0;
  wire n22__1_n_0;
  wire n22__27_carry__0_i_1_n_0;
  wire n22__27_carry__0_i_2_n_0;
  wire n22__27_carry__0_i_3_n_0;
  wire n22__27_carry__0_i_4_n_0;
  wire n22__27_carry__0_n_14;
  wire n22__27_carry__0_n_15;
  wire n22__27_carry__0_n_5;
  wire n22__27_carry__0_n_7;
  wire n22__27_carry_i_10_n_0;
  wire n22__27_carry_i_11_n_0;
  wire n22__27_carry_i_12_n_0;
  wire n22__27_carry_i_13_n_0;
  wire n22__27_carry_i_14_n_0;
  wire n22__27_carry_i_15_n_0;
  wire n22__27_carry_i_16_n_0;
  wire n22__27_carry_i_17_n_0;
  wire n22__27_carry_i_18_n_0;
  wire n22__27_carry_i_19_n_0;
  wire n22__27_carry_i_1_n_0;
  wire n22__27_carry_i_20_n_0;
  wire n22__27_carry_i_2_n_0;
  wire n22__27_carry_i_3_n_0;
  wire n22__27_carry_i_4_n_0;
  wire n22__27_carry_i_5_n_0;
  wire n22__27_carry_i_6_n_0;
  wire n22__27_carry_i_7_n_0;
  wire n22__27_carry_i_8_n_0;
  wire n22__27_carry_i_9_n_0;
  wire n22__27_carry_n_0;
  wire n22__27_carry_n_1;
  wire n22__27_carry_n_10;
  wire n22__27_carry_n_11;
  wire n22__27_carry_n_12;
  wire n22__27_carry_n_13;
  wire n22__27_carry_n_14;
  wire n22__27_carry_n_15;
  wire n22__27_carry_n_2;
  wire n22__27_carry_n_3;
  wire n22__27_carry_n_4;
  wire n22__27_carry_n_5;
  wire n22__27_carry_n_6;
  wire n22__27_carry_n_7;
  wire n22__27_carry_n_8;
  wire n22__27_carry_n_9;
  wire n22__2_n_0;
  wire n22__3_n_0;
  wire n22__4_n_0;
  wire n22__56_carry__0_i_1_n_0;
  wire n22__56_carry__0_n_15;
  wire n22__56_carry_i_10_n_0;
  wire n22__56_carry_i_11_n_0;
  wire n22__56_carry_i_12_n_0;
  wire n22__56_carry_i_13_n_0;
  wire n22__56_carry_i_14_n_0;
  wire n22__56_carry_i_15_n_0;
  wire n22__56_carry_i_1_n_0;
  wire n22__56_carry_i_2_n_0;
  wire n22__56_carry_i_3_n_0;
  wire n22__56_carry_i_4_n_0;
  wire n22__56_carry_i_5_n_0;
  wire n22__56_carry_i_6_n_0;
  wire n22__56_carry_i_7_n_0;
  wire n22__56_carry_i_8_n_0;
  wire n22__56_carry_i_9_n_0;
  wire n22__56_carry_n_0;
  wire n22__56_carry_n_1;
  wire n22__56_carry_n_10;
  wire n22__56_carry_n_11;
  wire n22__56_carry_n_12;
  wire n22__56_carry_n_13;
  wire n22__56_carry_n_14;
  wire n22__56_carry_n_15;
  wire n22__56_carry_n_2;
  wire n22__56_carry_n_3;
  wire n22__56_carry_n_4;
  wire n22__56_carry_n_5;
  wire n22__56_carry_n_6;
  wire n22__56_carry_n_7;
  wire n22__56_carry_n_8;
  wire n22__56_carry_n_9;
  wire n22__5_n_0;
  wire n22__6_n_0;
  wire n22__81_carry__0_i_1_n_0;
  wire n22__81_carry__0_i_2_n_0;
  wire n22__81_carry__0_i_3_n_0;
  wire n22__81_carry__0_i_4_n_0;
  wire n22__81_carry__0_i_5_n_0;
  wire n22__81_carry__0_i_6_n_0;
  wire n22__81_carry__0_i_7_n_0;
  wire n22__81_carry__0_n_5;
  wire n22__81_carry__0_n_6;
  wire n22__81_carry__0_n_7;
  wire n22__81_carry_i_10_n_0;
  wire n22__81_carry_i_11_n_0;
  wire n22__81_carry_i_12_n_0;
  wire n22__81_carry_i_13_n_0;
  wire n22__81_carry_i_14_n_0;
  wire n22__81_carry_i_15_n_0;
  wire n22__81_carry_i_1_n_0;
  wire n22__81_carry_i_2_n_0;
  wire n22__81_carry_i_3_n_0;
  wire n22__81_carry_i_4_n_0;
  wire n22__81_carry_i_5_n_0;
  wire n22__81_carry_i_6_n_0;
  wire n22__81_carry_i_7_n_0;
  wire n22__81_carry_i_8_n_0;
  wire n22__81_carry_i_9_n_0;
  wire n22__81_carry_n_0;
  wire n22__81_carry_n_1;
  wire n22__81_carry_n_2;
  wire n22__81_carry_n_3;
  wire n22__81_carry_n_4;
  wire n22__81_carry_n_5;
  wire n22__81_carry_n_6;
  wire n22__81_carry_n_7;
  wire n22_n_0;
  wire [7:0]n23;
  wire [7:0]n24;
  wire n25__0_carry__0_i_1_n_0;
  wire n25__0_carry__0_i_2_n_0;
  wire n25__0_carry__0_i_3_n_0;
  wire n25__0_carry__0_i_4_n_0;
  wire n25__0_carry__0_n_14;
  wire n25__0_carry__0_n_15;
  wire n25__0_carry__0_n_5;
  wire n25__0_carry__0_n_7;
  wire n25__0_carry_i_10_n_0;
  wire n25__0_carry_i_11_n_0;
  wire n25__0_carry_i_12_n_0;
  wire n25__0_carry_i_13_n_0;
  wire n25__0_carry_i_14_n_0;
  wire n25__0_carry_i_15_n_0;
  wire n25__0_carry_i_16_n_0;
  wire n25__0_carry_i_17_n_0;
  wire n25__0_carry_i_18_n_0;
  wire n25__0_carry_i_19_n_0;
  wire n25__0_carry_i_1_n_0;
  wire n25__0_carry_i_20_n_0;
  wire n25__0_carry_i_2_n_0;
  wire n25__0_carry_i_3_n_0;
  wire n25__0_carry_i_4_n_0;
  wire n25__0_carry_i_5_n_0;
  wire n25__0_carry_i_6_n_0;
  wire n25__0_carry_i_7_n_0;
  wire n25__0_carry_i_8_n_0;
  wire n25__0_carry_i_9_n_0;
  wire n25__0_carry_n_0;
  wire n25__0_carry_n_1;
  wire n25__0_carry_n_10;
  wire n25__0_carry_n_11;
  wire n25__0_carry_n_12;
  wire n25__0_carry_n_2;
  wire n25__0_carry_n_3;
  wire n25__0_carry_n_4;
  wire n25__0_carry_n_5;
  wire n25__0_carry_n_6;
  wire n25__0_carry_n_7;
  wire n25__0_carry_n_8;
  wire n25__0_carry_n_9;
  wire n25__27_carry__0_i_1_n_0;
  wire n25__27_carry__0_i_2_n_0;
  wire n25__27_carry__0_i_3_n_0;
  wire n25__27_carry__0_i_4_n_0;
  wire n25__27_carry__0_n_14;
  wire n25__27_carry__0_n_15;
  wire n25__27_carry__0_n_5;
  wire n25__27_carry__0_n_7;
  wire n25__27_carry_i_10_n_0;
  wire n25__27_carry_i_11_n_0;
  wire n25__27_carry_i_12_n_0;
  wire n25__27_carry_i_13_n_0;
  wire n25__27_carry_i_14_n_0;
  wire n25__27_carry_i_15_n_0;
  wire n25__27_carry_i_16_n_0;
  wire n25__27_carry_i_17_n_0;
  wire n25__27_carry_i_18_n_0;
  wire n25__27_carry_i_19_n_0;
  wire n25__27_carry_i_1_n_0;
  wire n25__27_carry_i_20_n_0;
  wire n25__27_carry_i_2_n_0;
  wire n25__27_carry_i_3_n_0;
  wire n25__27_carry_i_4_n_0;
  wire n25__27_carry_i_5_n_0;
  wire n25__27_carry_i_6_n_0;
  wire n25__27_carry_i_7_n_0;
  wire n25__27_carry_i_8_n_0;
  wire n25__27_carry_i_9_n_0;
  wire n25__27_carry_n_0;
  wire n25__27_carry_n_1;
  wire n25__27_carry_n_10;
  wire n25__27_carry_n_11;
  wire n25__27_carry_n_12;
  wire n25__27_carry_n_13;
  wire n25__27_carry_n_14;
  wire n25__27_carry_n_15;
  wire n25__27_carry_n_2;
  wire n25__27_carry_n_3;
  wire n25__27_carry_n_4;
  wire n25__27_carry_n_5;
  wire n25__27_carry_n_6;
  wire n25__27_carry_n_7;
  wire n25__27_carry_n_8;
  wire n25__27_carry_n_9;
  wire n25__56_carry__0_i_1_n_0;
  wire n25__56_carry__0_n_15;
  wire n25__56_carry_i_10_n_0;
  wire n25__56_carry_i_11_n_0;
  wire n25__56_carry_i_12_n_0;
  wire n25__56_carry_i_13_n_0;
  wire n25__56_carry_i_14_n_0;
  wire n25__56_carry_i_15_n_0;
  wire n25__56_carry_i_1_n_0;
  wire n25__56_carry_i_2_n_0;
  wire n25__56_carry_i_3_n_0;
  wire n25__56_carry_i_4_n_0;
  wire n25__56_carry_i_5_n_0;
  wire n25__56_carry_i_6_n_0;
  wire n25__56_carry_i_7_n_0;
  wire n25__56_carry_i_8_n_0;
  wire n25__56_carry_i_9_n_0;
  wire n25__56_carry_n_0;
  wire n25__56_carry_n_1;
  wire n25__56_carry_n_10;
  wire n25__56_carry_n_11;
  wire n25__56_carry_n_12;
  wire n25__56_carry_n_13;
  wire n25__56_carry_n_14;
  wire n25__56_carry_n_15;
  wire n25__56_carry_n_2;
  wire n25__56_carry_n_3;
  wire n25__56_carry_n_4;
  wire n25__56_carry_n_5;
  wire n25__56_carry_n_6;
  wire n25__56_carry_n_7;
  wire n25__56_carry_n_8;
  wire n25__56_carry_n_9;
  wire n25__81_carry__0_i_1_n_0;
  wire n25__81_carry__0_i_2_n_0;
  wire n25__81_carry__0_i_3_n_0;
  wire n25__81_carry__0_i_4_n_0;
  wire n25__81_carry__0_i_5_n_0;
  wire n25__81_carry__0_i_6_n_0;
  wire n25__81_carry__0_i_7_n_0;
  wire n25__81_carry__0_n_5;
  wire n25__81_carry__0_n_6;
  wire n25__81_carry__0_n_7;
  wire n25__81_carry_i_10_n_0;
  wire n25__81_carry_i_11_n_0;
  wire n25__81_carry_i_12_n_0;
  wire n25__81_carry_i_13_n_0;
  wire n25__81_carry_i_14_n_0;
  wire n25__81_carry_i_15_n_0;
  wire n25__81_carry_i_1_n_0;
  wire n25__81_carry_i_2_n_0;
  wire n25__81_carry_i_3_n_0;
  wire n25__81_carry_i_4_n_0;
  wire n25__81_carry_i_5_n_0;
  wire n25__81_carry_i_6_n_0;
  wire n25__81_carry_i_7_n_0;
  wire n25__81_carry_i_8_n_0;
  wire n25__81_carry_i_9_n_0;
  wire n25__81_carry_n_0;
  wire n25__81_carry_n_1;
  wire n25__81_carry_n_2;
  wire n25__81_carry_n_3;
  wire n25__81_carry_n_4;
  wire n25__81_carry_n_5;
  wire n25__81_carry_n_6;
  wire n25__81_carry_n_7;
  wire [7:0]n26;
  wire [7:0]n27;
  wire [7:0]n28;
  wire [7:0]n29;
  wire \n29[7]_i_2_n_0 ;
  wire \n29[7]_i_3_n_0 ;
  wire \n29[7]_i_4_n_0 ;
  wire \n29[7]_i_5_n_0 ;
  wire \n29[7]_i_6_n_0 ;
  wire \n29[7]_i_7_n_0 ;
  wire \n29[7]_i_8_n_0 ;
  wire \n29[7]_i_9_n_0 ;
  wire \n29_reg[7]_i_1_n_1 ;
  wire \n29_reg[7]_i_1_n_2 ;
  wire \n29_reg[7]_i_1_n_3 ;
  wire \n29_reg[7]_i_1_n_4 ;
  wire \n29_reg[7]_i_1_n_5 ;
  wire \n29_reg[7]_i_1_n_6 ;
  wire \n29_reg[7]_i_1_n_7 ;
  wire [7:7]n30;
  wire [7:0]n31;
  wire \n33[10]_i_1_n_0 ;
  wire \n33[11]_i_1_n_0 ;
  wire \n33[12]_i_1_n_0 ;
  wire \n33[12]_i_2_n_0 ;
  wire \n33[13]_i_1_n_0 ;
  wire \n33[14]_i_1_n_0 ;
  wire \n33[14]_i_2_n_0 ;
  wire \n33[15]_i_2_n_0 ;
  wire \n33[2]_i_1_n_0 ;
  wire \n33[3]_i_1_n_0 ;
  wire \n33[4]_i_1_n_0 ;
  wire \n33[4]_i_2_n_0 ;
  wire \n33[5]_i_1_n_0 ;
  wire \n33[6]_i_1_n_0 ;
  wire \n33[6]_i_2_n_0 ;
  wire \n33[7]_i_2_n_0 ;
  wire \n33[9]_i_1_n_0 ;
  wire [7:0]n341_out;
  wire [7:1]n350_out;
  wire \n37[12]_i_2_n_0 ;
  wire \n37[14]_i_2_n_0 ;
  wire \n37[15]_i_2_n_0 ;
  wire \n37[4]_i_2_n_0 ;
  wire \n37[6]_i_2_n_0 ;
  wire \n37[7]_i_2_n_0 ;
  wire [7:0]n4;
  wire \n7_reg_n_0_[0] ;
  wire \n7_reg_n_0_[1] ;
  wire \n7_reg_n_0_[2] ;
  wire \n7_reg_n_0_[3] ;
  wire \n7_reg_n_0_[4] ;
  wire \n7_reg_n_0_[5] ;
  wire \n7_reg_n_0_[6] ;
  wire \n7_reg_n_0_[7] ;
  wire \n8_reg_n_0_[0] ;
  wire \n8_reg_n_0_[1] ;
  wire \n8_reg_n_0_[2] ;
  wire \n8_reg_n_0_[3] ;
  wire \n8_reg_n_0_[4] ;
  wire \n8_reg_n_0_[5] ;
  wire \n8_reg_n_0_[6] ;
  wire \n8_reg_n_0_[7] ;
  wire \n9_reg_n_0_[0] ;
  wire \n9_reg_n_0_[1] ;
  wire \n9_reg_n_0_[2] ;
  wire \n9_reg_n_0_[3] ;
  wire \n9_reg_n_0_[4] ;
  wire \n9_reg_n_0_[5] ;
  wire \n9_reg_n_0_[6] ;
  wire \n9_reg_n_0_[7] ;
  wire rst_i;
  wire [15:0]s2_3;
  wire [15:0]NLW_n11_reg_CASDOUTA_UNCONNECTED;
  wire [15:0]NLW_n11_reg_CASDOUTB_UNCONNECTED;
  wire [1:0]NLW_n11_reg_CASDOUTPA_UNCONNECTED;
  wire [1:0]NLW_n11_reg_CASDOUTPB_UNCONNECTED;
  wire [15:0]NLW_n11_reg_DOUTBDOUT_UNCONNECTED;
  wire [1:0]NLW_n11_reg_DOUTPADOUTP_UNCONNECTED;
  wire [1:0]NLW_n11_reg_DOUTPBDOUTP_UNCONNECTED;
  wire [2:0]NLW_n14__0_carry_O_UNCONNECTED;
  wire [7:1]NLW_n14__0_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n14__0_carry__0_O_UNCONNECTED;
  wire [7:1]NLW_n14__27_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n14__27_carry__0_O_UNCONNECTED;
  wire [7:0]NLW_n14__56_carry__0_CO_UNCONNECTED;
  wire [7:1]NLW_n14__56_carry__0_O_UNCONNECTED;
  wire [3:0]NLW_n14__81_carry_O_UNCONNECTED;
  wire [7:3]NLW_n14__81_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n14__81_carry__0_O_UNCONNECTED;
  wire [2:0]NLW_n17__0_carry_O_UNCONNECTED;
  wire [7:1]NLW_n17__0_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n17__0_carry__0_O_UNCONNECTED;
  wire [7:1]NLW_n17__27_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n17__27_carry__0_O_UNCONNECTED;
  wire [7:0]NLW_n17__56_carry__0_CO_UNCONNECTED;
  wire [7:1]NLW_n17__56_carry__0_O_UNCONNECTED;
  wire [3:0]NLW_n17__81_carry_O_UNCONNECTED;
  wire [7:3]NLW_n17__81_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n17__81_carry__0_O_UNCONNECTED;
  wire [7:7]NLW_n20_carry_CO_UNCONNECTED;
  wire [2:0]NLW_n22__0_carry_O_UNCONNECTED;
  wire [7:1]NLW_n22__0_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n22__0_carry__0_O_UNCONNECTED;
  wire [7:1]NLW_n22__27_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n22__27_carry__0_O_UNCONNECTED;
  wire [7:0]NLW_n22__56_carry__0_CO_UNCONNECTED;
  wire [7:1]NLW_n22__56_carry__0_O_UNCONNECTED;
  wire [3:0]NLW_n22__81_carry_O_UNCONNECTED;
  wire [7:3]NLW_n22__81_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n22__81_carry__0_O_UNCONNECTED;
  wire [2:0]NLW_n25__0_carry_O_UNCONNECTED;
  wire [7:1]NLW_n25__0_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n25__0_carry__0_O_UNCONNECTED;
  wire [7:1]NLW_n25__27_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n25__27_carry__0_O_UNCONNECTED;
  wire [7:0]NLW_n25__56_carry__0_CO_UNCONNECTED;
  wire [7:1]NLW_n25__56_carry__0_O_UNCONNECTED;
  wire [3:0]NLW_n25__81_carry_O_UNCONNECTED;
  wire [7:3]NLW_n25__81_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n25__81_carry__0_O_UNCONNECTED;
  wire [7:7]\NLW_n29_reg[7]_i_1_CO_UNCONNECTED ;

  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[0] ),
        .Q(n10[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[1] ),
        .Q(n10[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[2] ),
        .Q(n10[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[3] ),
        .Q(n10[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[4] ),
        .Q(n10[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[5] ),
        .Q(n10[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[6] ),
        .Q(n10[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[7] ),
        .Q(n10[7]),
        .R(rst_i));
  (* \MEM.PORTA.DATA_BIT_LAYOUT  = "p0_d16" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RDADDR_COLLISION_HWCONFIG = "PERFORMANCE" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s25/n11" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "15" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "1023" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "15" *) 
  RAMB18E2 #(
    .CASCADE_ORDER_A("NONE"),
    .CASCADE_ORDER_B("NONE"),
    .CLOCK_DOMAINS("INDEPENDENT"),
    .DOA_REG(0),
    .DOB_REG(0),
    .ENADDRENA("FALSE"),
    .ENADDRENB("FALSE"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h7DE87EEA7EEB7EED7EEE7FF07FF17FF37FF57FF67FF87FF97FFB7FFC7FFE7F00),
    .INIT_01(256'h76D077D177D378D479D679D77AD97ADA7ADC7BDD7BDF7CE07CE27CE37DE57DE7),
    .INIT_02(256'h6BBA6CBB6CBC6DBE6EBF6FC070C270C371C572C673C773C974CA75CC75CD76CF),
    .INIT_03(256'h5BA65CA75DA85EAA5FAB60AC61AD62AE63B064B165B266B367B568B669B76AB8),
    .INIT_04(256'h489649974A984C994D9A4E9B4F9C519D529E539F54A055A157A258A359A45AA5),
    .INIT_05(256'h328A338A358B368C388C398D3A8E3C8F3D8F3F90409141924393449345944795),
    .INIT_06(256'h1A821C831D831F8320842284238525852685288629862B872C882E882F893089),
    .INIT_07(256'h0180038004800680078009800A800C800E800F80118112811481158117821882),
    .INIT_08(256'hE882EA81EB81ED81EE81F080F180F380F580F680F880F980FB80FC80FE800080),
    .INIT_09(256'hD089D188D388D487D686D786D985DA85DC85DD84DF84E083E283E383E582E782),
    .INIT_0A(256'hBA94BB93BC93BE92BF91C090C28FC38FC58EC68DC78CC98CCA8BCC8ACD8ACF89),
    .INIT_0B(256'hA6A4A7A3A8A2AAA1ABA0AC9FAD9EAE9DB09CB19BB29AB399B598B697B796B895),
    .INIT_0C(256'h96B797B698B599B39AB29BB19CB09DAE9EAD9FACA0ABA1AAA2A8A3A7A4A6A5A5),
    .INIT_0D(256'h8ACD8ACC8BCA8CC98CC78DC68EC58FC38FC290C091BF92BE93BC93BB94BA95B8),
    .INIT_0E(256'h82E583E383E283E084DF84DD85DC85DA85D986D786D687D488D388D189D089CF),
    .INIT_0F(256'h80FE80FC80FB80F980F880F680F580F380F180F081EE81ED81EB81EA82E882E7),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .RDADDRCHANGEA("FALSE"),
    .RDADDRCHANGEB("FALSE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(0),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SLEEP_ASYNC("FALSE"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    n11_reg
       (.ADDRARDADDR({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .ADDRBWRADDR({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .ADDRENA(1'b0),
        .ADDRENB(1'b0),
        .CASDIMUXA(1'b0),
        .CASDIMUXB(1'b0),
        .CASDINA({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .CASDINB({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .CASDINPA({1'b0,1'b0}),
        .CASDINPB({1'b0,1'b0}),
        .CASDOMUXA(1'b0),
        .CASDOMUXB(1'b0),
        .CASDOMUXEN_A(1'b1),
        .CASDOMUXEN_B(1'b1),
        .CASDOUTA(NLW_n11_reg_CASDOUTA_UNCONNECTED[15:0]),
        .CASDOUTB(NLW_n11_reg_CASDOUTB_UNCONNECTED[15:0]),
        .CASDOUTPA(NLW_n11_reg_CASDOUTPA_UNCONNECTED[1:0]),
        .CASDOUTPB(NLW_n11_reg_CASDOUTPB_UNCONNECTED[1:0]),
        .CASOREGIMUXA(1'b0),
        .CASOREGIMUXB(1'b0),
        .CASOREGIMUXEN_A(1'b1),
        .CASOREGIMUXEN_B(1'b1),
        .CLKARDCLK(clk_i),
        .CLKBWRCLK(1'b0),
        .DINADIN({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DINBDIN({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DINPADINP({1'b0,1'b0}),
        .DINPBDINP({1'b1,1'b1}),
        .DOUTADOUT({B,n11_reg_n_40,n11_reg_n_41,n11_reg_n_42,n11_reg_n_43,n11_reg_n_44,n11_reg_n_45,n11_reg_n_46,n11_reg_n_47}),
        .DOUTBDOUT(NLW_n11_reg_DOUTBDOUT_UNCONNECTED[15:0]),
        .DOUTPADOUTP(NLW_n11_reg_DOUTPADOUTP_UNCONNECTED[1:0]),
        .DOUTPBDOUTP(NLW_n11_reg_DOUTPBDOUTP_UNCONNECTED[1:0]),
        .ENARDEN(enable_i),
        .ENBWREN(1'b0),
        .REGCEAREGCE(1'b1),
        .REGCEB(1'b1),
        .RSTRAMARSTRAM(1'b0),
        .RSTRAMB(1'b0),
        .RSTREGARSTREG(1'b0),
        .RSTREGB(1'b0),
        .SLEEP(1'b0),
        .WEA({1'b0,1'b0}),
        .WEBWE({1'b0,1'b0,1'b0,1'b0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__0_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__0_carry_n_0,n14__0_carry_n_1,n14__0_carry_n_2,n14__0_carry_n_3,n14__0_carry_n_4,n14__0_carry_n_5,n14__0_carry_n_6,n14__0_carry_n_7}),
        .DI({n14__0_carry_i_1_n_0,n14__0_carry_i_2_n_0,n14__0_carry_i_3_n_0,n14__0_carry_i_4_n_0,n14__0_carry_i_5_n_0,n14__0_carry_i_6_n_0,n14__0_carry_i_7_n_0,1'b0}),
        .O({n14__0_carry_n_8,n14__0_carry_n_9,n14__0_carry_n_10,n14__0_carry_n_11,n14__0_carry_n_12,NLW_n14__0_carry_O_UNCONNECTED[2:0]}),
        .S({n14__0_carry_i_8_n_0,n14__0_carry_i_9_n_0,n14__0_carry_i_10_n_0,n14__0_carry_i_11_n_0,n14__0_carry_i_12_n_0,n14__0_carry_i_13_n_0,n14__0_carry_i_14_n_0,n14__0_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__0_carry__0
       (.CI(n14__0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__0_carry__0_CO_UNCONNECTED[7:3],n14__0_carry__0_n_5,NLW_n14__0_carry__0_CO_UNCONNECTED[1],n14__0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14__0_carry__0_i_1_n_0,n14__0_carry__0_i_2_n_0}),
        .O({NLW_n14__0_carry__0_O_UNCONNECTED[7:2],n14__0_carry__0_n_14,n14__0_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n14__0_carry__0_i_3_n_0,n14__0_carry__0_i_4_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__0_carry__0_i_1
       (.I0(B[1]),
        .I1(n22_n_0),
        .I2(B[2]),
        .I3(n22__0_n_0),
        .O(n14__0_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n14__0_carry__0_i_2
       (.I0(B[2]),
        .I1(n22__1_n_0),
        .I2(B[1]),
        .I3(n22__0_n_0),
        .I4(B[0]),
        .I5(n22_n_0),
        .O(n14__0_carry__0_i_2_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n14__0_carry__0_i_3
       (.I0(n22__0_n_0),
        .I1(B[1]),
        .I2(B[2]),
        .I3(n22_n_0),
        .O(n14__0_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n14__0_carry__0_i_4
       (.I0(B[0]),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(B[2]),
        .I4(n22_n_0),
        .I5(B[1]),
        .O(n14__0_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__0_carry_i_1
       (.I0(B[2]),
        .I1(n22__2_n_0),
        .I2(B[1]),
        .I3(n22__1_n_0),
        .I4(B[0]),
        .I5(n22__0_n_0),
        .O(n14__0_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__0_carry_i_10
       (.I0(n14__0_carry_i_3_n_0),
        .I1(B[1]),
        .I2(n22__2_n_0),
        .I3(n14__0_carry_i_18_n_0),
        .I4(n22__1_n_0),
        .I5(B[0]),
        .O(n14__0_carry_i_10_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__0_carry_i_11
       (.I0(n14__0_carry_i_4_n_0),
        .I1(B[1]),
        .I2(n22__3_n_0),
        .I3(n14__0_carry_i_19_n_0),
        .I4(n22__2_n_0),
        .I5(B[0]),
        .O(n14__0_carry_i_11_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n14__0_carry_i_12
       (.I0(n22__4_n_0),
        .I1(n14__0_carry_i_20_n_0),
        .I2(n22__5_n_0),
        .I3(B[1]),
        .I4(n22__6_n_0),
        .I5(B[2]),
        .O(n14__0_carry_i_12_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n14__0_carry_i_13
       (.I0(n22__6_n_0),
        .I1(B[2]),
        .I2(n22__5_n_0),
        .I3(B[1]),
        .I4(B[0]),
        .I5(n22__4_n_0),
        .O(n14__0_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__0_carry_i_14
       (.I0(B[0]),
        .I1(n22__5_n_0),
        .I2(B[1]),
        .I3(n22__6_n_0),
        .O(n14__0_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__0_carry_i_15
       (.I0(n22__6_n_0),
        .I1(B[0]),
        .O(n14__0_carry_i_15_n_0));
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_16
       (.I0(n22__1_n_0),
        .I1(B[2]),
        .O(n14__0_carry_i_16_n_0));
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_17
       (.I0(n22__2_n_0),
        .I1(B[2]),
        .O(n14__0_carry_i_17_n_0));
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_18
       (.I0(n22__3_n_0),
        .I1(B[2]),
        .O(n14__0_carry_i_18_n_0));
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_19
       (.I0(n22__4_n_0),
        .I1(B[2]),
        .O(n14__0_carry_i_19_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__0_carry_i_2
       (.I0(B[2]),
        .I1(n22__3_n_0),
        .I2(B[1]),
        .I3(n22__2_n_0),
        .I4(B[0]),
        .I5(n22__1_n_0),
        .O(n14__0_carry_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__0_carry_i_20
       (.I0(n22__3_n_0),
        .I1(B[0]),
        .O(n14__0_carry_i_20_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__0_carry_i_3
       (.I0(B[2]),
        .I1(n22__4_n_0),
        .I2(B[1]),
        .I3(n22__3_n_0),
        .I4(B[0]),
        .I5(n22__2_n_0),
        .O(n14__0_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__0_carry_i_4
       (.I0(B[2]),
        .I1(n22__5_n_0),
        .I2(B[1]),
        .I3(n22__4_n_0),
        .I4(B[0]),
        .I5(n22__3_n_0),
        .O(n14__0_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n14__0_carry_i_5
       (.I0(B[1]),
        .I1(n22__4_n_0),
        .I2(B[2]),
        .I3(n22__5_n_0),
        .I4(n22__3_n_0),
        .I5(B[0]),
        .O(n14__0_carry_i_5_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__0_carry_i_6
       (.I0(B[1]),
        .I1(n22__5_n_0),
        .I2(B[2]),
        .I3(n22__6_n_0),
        .O(n14__0_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__0_carry_i_7
       (.I0(B[0]),
        .I1(n22__5_n_0),
        .O(n14__0_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n14__0_carry_i_8
       (.I0(n14__0_carry_i_1_n_0),
        .I1(B[1]),
        .I2(n22__0_n_0),
        .I3(n14__0_carry_i_16_n_0),
        .I4(n22_n_0),
        .I5(B[0]),
        .O(n14__0_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__0_carry_i_9
       (.I0(n14__0_carry_i_2_n_0),
        .I1(B[1]),
        .I2(n22__1_n_0),
        .I3(n14__0_carry_i_17_n_0),
        .I4(n22__0_n_0),
        .I5(B[0]),
        .O(n14__0_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__27_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__27_carry_n_0,n14__27_carry_n_1,n14__27_carry_n_2,n14__27_carry_n_3,n14__27_carry_n_4,n14__27_carry_n_5,n14__27_carry_n_6,n14__27_carry_n_7}),
        .DI({n14__27_carry_i_1_n_0,n14__27_carry_i_2_n_0,n14__27_carry_i_3_n_0,n14__27_carry_i_4_n_0,n14__27_carry_i_5_n_0,n14__27_carry_i_6_n_0,n14__27_carry_i_7_n_0,1'b0}),
        .O({n14__27_carry_n_8,n14__27_carry_n_9,n14__27_carry_n_10,n14__27_carry_n_11,n14__27_carry_n_12,n14__27_carry_n_13,n14__27_carry_n_14,n14__27_carry_n_15}),
        .S({n14__27_carry_i_8_n_0,n14__27_carry_i_9_n_0,n14__27_carry_i_10_n_0,n14__27_carry_i_11_n_0,n14__27_carry_i_12_n_0,n14__27_carry_i_13_n_0,n14__27_carry_i_14_n_0,n14__27_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__27_carry__0
       (.CI(n14__27_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__27_carry__0_CO_UNCONNECTED[7:3],n14__27_carry__0_n_5,NLW_n14__27_carry__0_CO_UNCONNECTED[1],n14__27_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14__27_carry__0_i_1_n_0,n14__27_carry__0_i_2_n_0}),
        .O({NLW_n14__27_carry__0_O_UNCONNECTED[7:2],n14__27_carry__0_n_14,n14__27_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n14__27_carry__0_i_3_n_0,n14__27_carry__0_i_4_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__27_carry__0_i_1
       (.I0(B[4]),
        .I1(n22_n_0),
        .I2(B[5]),
        .I3(n22__0_n_0),
        .O(n14__27_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n14__27_carry__0_i_2
       (.I0(B[5]),
        .I1(n22__1_n_0),
        .I2(B[4]),
        .I3(n22__0_n_0),
        .I4(B[3]),
        .I5(n22_n_0),
        .O(n14__27_carry__0_i_2_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n14__27_carry__0_i_3
       (.I0(n22__0_n_0),
        .I1(B[4]),
        .I2(B[5]),
        .I3(n22_n_0),
        .O(n14__27_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n14__27_carry__0_i_4
       (.I0(B[3]),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(B[5]),
        .I4(n22_n_0),
        .I5(B[4]),
        .O(n14__27_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__27_carry_i_1
       (.I0(B[5]),
        .I1(n22__2_n_0),
        .I2(B[4]),
        .I3(n22__1_n_0),
        .I4(B[3]),
        .I5(n22__0_n_0),
        .O(n14__27_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__27_carry_i_10
       (.I0(n14__27_carry_i_3_n_0),
        .I1(B[4]),
        .I2(n22__2_n_0),
        .I3(n14__27_carry_i_18_n_0),
        .I4(n22__1_n_0),
        .I5(B[3]),
        .O(n14__27_carry_i_10_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__27_carry_i_11
       (.I0(n14__27_carry_i_4_n_0),
        .I1(B[4]),
        .I2(n22__3_n_0),
        .I3(n14__27_carry_i_19_n_0),
        .I4(n22__2_n_0),
        .I5(B[3]),
        .O(n14__27_carry_i_11_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n14__27_carry_i_12
       (.I0(n22__4_n_0),
        .I1(n14__27_carry_i_20_n_0),
        .I2(n22__5_n_0),
        .I3(B[4]),
        .I4(n22__6_n_0),
        .I5(B[5]),
        .O(n14__27_carry_i_12_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n14__27_carry_i_13
       (.I0(n22__6_n_0),
        .I1(B[5]),
        .I2(n22__5_n_0),
        .I3(B[4]),
        .I4(B[3]),
        .I5(n22__4_n_0),
        .O(n14__27_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__27_carry_i_14
       (.I0(B[3]),
        .I1(n22__5_n_0),
        .I2(B[4]),
        .I3(n22__6_n_0),
        .O(n14__27_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__27_carry_i_15
       (.I0(n22__6_n_0),
        .I1(B[3]),
        .O(n14__27_carry_i_15_n_0));
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_16
       (.I0(n22__1_n_0),
        .I1(B[5]),
        .O(n14__27_carry_i_16_n_0));
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_17
       (.I0(n22__2_n_0),
        .I1(B[5]),
        .O(n14__27_carry_i_17_n_0));
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_18
       (.I0(n22__3_n_0),
        .I1(B[5]),
        .O(n14__27_carry_i_18_n_0));
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_19
       (.I0(n22__4_n_0),
        .I1(B[5]),
        .O(n14__27_carry_i_19_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__27_carry_i_2
       (.I0(B[5]),
        .I1(n22__3_n_0),
        .I2(B[4]),
        .I3(n22__2_n_0),
        .I4(B[3]),
        .I5(n22__1_n_0),
        .O(n14__27_carry_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n14__27_carry_i_20
       (.I0(n22__3_n_0),
        .I1(B[3]),
        .O(n14__27_carry_i_20_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__27_carry_i_3
       (.I0(B[5]),
        .I1(n22__4_n_0),
        .I2(B[4]),
        .I3(n22__3_n_0),
        .I4(B[3]),
        .I5(n22__2_n_0),
        .O(n14__27_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n14__27_carry_i_4
       (.I0(B[5]),
        .I1(n22__5_n_0),
        .I2(B[4]),
        .I3(n22__4_n_0),
        .I4(B[3]),
        .I5(n22__3_n_0),
        .O(n14__27_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n14__27_carry_i_5
       (.I0(B[4]),
        .I1(n22__4_n_0),
        .I2(B[5]),
        .I3(n22__5_n_0),
        .I4(n22__3_n_0),
        .I5(B[3]),
        .O(n14__27_carry_i_5_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__27_carry_i_6
       (.I0(B[4]),
        .I1(n22__5_n_0),
        .I2(B[5]),
        .I3(n22__6_n_0),
        .O(n14__27_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__27_carry_i_7
       (.I0(B[3]),
        .I1(n22__5_n_0),
        .O(n14__27_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n14__27_carry_i_8
       (.I0(n14__27_carry_i_1_n_0),
        .I1(B[4]),
        .I2(n22__0_n_0),
        .I3(n14__27_carry_i_16_n_0),
        .I4(n22_n_0),
        .I5(B[3]),
        .O(n14__27_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n14__27_carry_i_9
       (.I0(n14__27_carry_i_2_n_0),
        .I1(B[4]),
        .I2(n22__1_n_0),
        .I3(n14__27_carry_i_17_n_0),
        .I4(n22__0_n_0),
        .I5(B[3]),
        .O(n14__27_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__56_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__56_carry_n_0,n14__56_carry_n_1,n14__56_carry_n_2,n14__56_carry_n_3,n14__56_carry_n_4,n14__56_carry_n_5,n14__56_carry_n_6,n14__56_carry_n_7}),
        .DI({n14__56_carry_i_1_n_0,n14__56_carry_i_2_n_0,n14__56_carry_i_3_n_0,n14__56_carry_i_4_n_0,n14__56_carry_i_5_n_0,n14__56_carry_i_6_n_0,n14__56_carry_i_7_n_0,1'b0}),
        .O({n14__56_carry_n_8,n14__56_carry_n_9,n14__56_carry_n_10,n14__56_carry_n_11,n14__56_carry_n_12,n14__56_carry_n_13,n14__56_carry_n_14,n14__56_carry_n_15}),
        .S({n14__56_carry_i_8_n_0,n14__56_carry_i_9_n_0,n14__56_carry_i_10_n_0,n14__56_carry_i_11_n_0,n14__56_carry_i_12_n_0,n14__56_carry_i_13_n_0,n14__56_carry_i_14_n_0,n14__56_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__56_carry__0
       (.CI(n14__56_carry_n_0),
        .CI_TOP(1'b0),
        .CO(NLW_n14__56_carry__0_CO_UNCONNECTED[7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_n14__56_carry__0_O_UNCONNECTED[7:1],n14__56_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14__56_carry__0_i_1_n_0}));
  LUT4 #(
    .INIT(16'hE53F)) 
    n14__56_carry__0_i_1
       (.I0(B[6]),
        .I1(n22__0_n_0),
        .I2(B[7]),
        .I3(n22_n_0),
        .O(n14__56_carry__0_i_1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__56_carry_i_1
       (.I0(B[7]),
        .I1(n22__1_n_0),
        .I2(B[6]),
        .I3(n22__0_n_0),
        .O(n14__56_carry_i_1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n14__56_carry_i_10
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(B[7]),
        .I3(n22__1_n_0),
        .I4(B[6]),
        .O(n14__56_carry_i_10_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n14__56_carry_i_11
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(B[7]),
        .I3(n22__2_n_0),
        .I4(B[6]),
        .O(n14__56_carry_i_11_n_0));
  LUT5 #(
    .INIT(32'h9F606060)) 
    n14__56_carry_i_12
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(B[7]),
        .I3(n22__3_n_0),
        .I4(B[6]),
        .O(n14__56_carry_i_12_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n14__56_carry_i_13
       (.I0(B[7]),
        .I1(n22__5_n_0),
        .I2(B[6]),
        .I3(n22__4_n_0),
        .O(n14__56_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h8777)) 
    n14__56_carry_i_14
       (.I0(B[7]),
        .I1(n22__6_n_0),
        .I2(B[6]),
        .I3(n22__5_n_0),
        .O(n14__56_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__56_carry_i_15
       (.I0(n22__6_n_0),
        .I1(B[6]),
        .O(n14__56_carry_i_15_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__56_carry_i_2
       (.I0(B[7]),
        .I1(n22__2_n_0),
        .I2(B[6]),
        .I3(n22__1_n_0),
        .O(n14__56_carry_i_2_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__56_carry_i_3
       (.I0(B[7]),
        .I1(n22__3_n_0),
        .I2(B[6]),
        .I3(n22__2_n_0),
        .O(n14__56_carry_i_3_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n14__56_carry_i_4
       (.I0(B[7]),
        .I1(n22__4_n_0),
        .I2(B[6]),
        .I3(n22__3_n_0),
        .O(n14__56_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n14__56_carry_i_5
       (.I0(n22__5_n_0),
        .I1(B[7]),
        .O(n14__56_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__56_carry_i_6
       (.I0(B[7]),
        .I1(n22__5_n_0),
        .O(n14__56_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n14__56_carry_i_7
       (.I0(n22__6_n_0),
        .I1(B[7]),
        .O(n14__56_carry_i_7_n_0));
  LUT5 #(
    .INIT(32'h738CC0C0)) 
    n14__56_carry_i_8
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(B[7]),
        .I3(n22_n_0),
        .I4(B[6]),
        .O(n14__56_carry_i_8_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n14__56_carry_i_9
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(B[7]),
        .I3(n22__0_n_0),
        .I4(B[6]),
        .O(n14__56_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__81_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__81_carry_n_0,n14__81_carry_n_1,n14__81_carry_n_2,n14__81_carry_n_3,n14__81_carry_n_4,n14__81_carry_n_5,n14__81_carry_n_6,n14__81_carry_n_7}),
        .DI({n14__81_carry_i_1_n_0,n14__81_carry_i_2_n_0,n14__81_carry_i_3_n_0,n14__81_carry_i_4_n_0,n14__81_carry_i_5_n_0,n14__81_carry_i_6_n_0,n14__81_carry_i_7_n_0,1'b0}),
        .O({n15[3:0],NLW_n14__81_carry_O_UNCONNECTED[3:0]}),
        .S({n14__81_carry_i_8_n_0,n14__81_carry_i_9_n_0,n14__81_carry_i_10_n_0,n14__81_carry_i_11_n_0,n14__81_carry_i_12_n_0,n14__81_carry_i_13_n_0,n14__81_carry_i_14_n_0,n14__81_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__81_carry__0
       (.CI(n14__81_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__81_carry__0_CO_UNCONNECTED[7:3],n14__81_carry__0_n_5,n14__81_carry__0_n_6,n14__81_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n14__81_carry__0_i_1_n_0,n14__81_carry__0_i_2_n_0,n14__81_carry__0_i_3_n_0}),
        .O({NLW_n14__81_carry__0_O_UNCONNECTED[7:4],n15[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n14__81_carry__0_i_4_n_0,n14__81_carry__0_i_5_n_0,n14__81_carry__0_i_6_n_0,n14__81_carry__0_i_7_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry__0_i_1
       (.I0(n14__27_carry__0_n_14),
        .I1(n14__56_carry_n_9),
        .O(n14__81_carry__0_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry__0_i_2
       (.I0(n14__27_carry__0_n_15),
        .I1(n14__56_carry_n_10),
        .O(n14__81_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry__0_i_3
       (.I0(n14__56_carry_n_11),
        .I1(n14__27_carry_n_8),
        .I2(n14__0_carry__0_n_5),
        .O(n14__81_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n14__81_carry__0_i_4
       (.I0(n14__27_carry__0_n_5),
        .I1(n14__56_carry_n_8),
        .I2(n14__56_carry__0_n_15),
        .O(n14__81_carry__0_i_4_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__81_carry__0_i_5
       (.I0(n14__27_carry__0_n_14),
        .I1(n14__56_carry_n_9),
        .I2(n14__56_carry_n_8),
        .I3(n14__27_carry__0_n_5),
        .O(n14__81_carry__0_i_5_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__81_carry__0_i_6
       (.I0(n14__27_carry__0_n_15),
        .I1(n14__56_carry_n_10),
        .I2(n14__56_carry_n_9),
        .I3(n14__27_carry__0_n_14),
        .O(n14__81_carry__0_i_6_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n14__81_carry__0_i_7
       (.I0(n14__0_carry__0_n_5),
        .I1(n14__27_carry_n_8),
        .I2(n14__56_carry_n_11),
        .I3(n14__56_carry_n_10),
        .I4(n14__27_carry__0_n_15),
        .O(n14__81_carry__0_i_7_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry_i_1
       (.I0(n14__56_carry_n_12),
        .I1(n14__27_carry_n_9),
        .I2(n14__0_carry__0_n_14),
        .O(n14__81_carry_i_1_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_10
       (.I0(n14__56_carry_n_13),
        .I1(n14__27_carry_n_10),
        .I2(n14__0_carry__0_n_15),
        .I3(n14__81_carry_i_3_n_0),
        .O(n14__81_carry_i_10_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_11
       (.I0(n14__56_carry_n_14),
        .I1(n14__27_carry_n_11),
        .I2(n14__0_carry_n_8),
        .I3(n14__81_carry_i_4_n_0),
        .O(n14__81_carry_i_11_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_12
       (.I0(n14__56_carry_n_15),
        .I1(n14__27_carry_n_12),
        .I2(n14__0_carry_n_9),
        .I3(n14__81_carry_i_5_n_0),
        .O(n14__81_carry_i_12_n_0));
  LUT4 #(
    .INIT(16'h9666)) 
    n14__81_carry_i_13
       (.I0(n14__27_carry_n_13),
        .I1(n14__0_carry_n_10),
        .I2(n14__0_carry_n_11),
        .I3(n14__27_carry_n_14),
        .O(n14__81_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__81_carry_i_14
       (.I0(n14__0_carry_n_12),
        .I1(n14__27_carry_n_15),
        .I2(n14__27_carry_n_14),
        .I3(n14__0_carry_n_11),
        .O(n14__81_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n14__81_carry_i_15
       (.I0(n14__0_carry_n_12),
        .I1(n14__27_carry_n_15),
        .O(n14__81_carry_i_15_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry_i_2
       (.I0(n14__56_carry_n_13),
        .I1(n14__27_carry_n_10),
        .I2(n14__0_carry__0_n_15),
        .O(n14__81_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry_i_3
       (.I0(n14__56_carry_n_14),
        .I1(n14__27_carry_n_11),
        .I2(n14__0_carry_n_8),
        .O(n14__81_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14__81_carry_i_4
       (.I0(n14__56_carry_n_15),
        .I1(n14__27_carry_n_12),
        .I2(n14__0_carry_n_9),
        .O(n14__81_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry_i_5
       (.I0(n14__27_carry_n_13),
        .I1(n14__0_carry_n_10),
        .O(n14__81_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry_i_6
       (.I0(n14__0_carry_n_11),
        .I1(n14__27_carry_n_14),
        .O(n14__81_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__81_carry_i_7
       (.I0(n14__0_carry_n_12),
        .I1(n14__27_carry_n_15),
        .O(n14__81_carry_i_7_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_8
       (.I0(n14__81_carry_i_1_n_0),
        .I1(n14__27_carry_n_8),
        .I2(n14__56_carry_n_11),
        .I3(n14__0_carry__0_n_5),
        .O(n14__81_carry_i_8_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n14__81_carry_i_9
       (.I0(n14__56_carry_n_12),
        .I1(n14__27_carry_n_9),
        .I2(n14__0_carry__0_n_14),
        .I3(n14__81_carry_i_2_n_0),
        .O(n14__81_carry_i_9_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[0]),
        .Q(\n16_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[1]),
        .Q(\n16_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[2]),
        .Q(\n16_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[3]),
        .Q(\n16_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[4]),
        .Q(\n16_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[5]),
        .Q(\n16_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[6]),
        .Q(\n16_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[7]),
        .Q(\n16_reg_n_0_[7] ),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__0_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n17__0_carry_n_0,n17__0_carry_n_1,n17__0_carry_n_2,n17__0_carry_n_3,n17__0_carry_n_4,n17__0_carry_n_5,n17__0_carry_n_6,n17__0_carry_n_7}),
        .DI({n17__0_carry_i_1_n_0,n17__0_carry_i_2_n_0,n17__0_carry_i_3_n_0,n17__0_carry_i_4_n_0,n17__0_carry_i_5_n_0,n17__0_carry_i_6_n_0,n17__0_carry_i_7_n_0,1'b0}),
        .O({n17__0_carry_n_8,n17__0_carry_n_9,n17__0_carry_n_10,n17__0_carry_n_11,n17__0_carry_n_12,NLW_n17__0_carry_O_UNCONNECTED[2:0]}),
        .S({n17__0_carry_i_8_n_0,n17__0_carry_i_9_n_0,n17__0_carry_i_10_n_0,n17__0_carry_i_11_n_0,n17__0_carry_i_12_n_0,n17__0_carry_i_13_n_0,n17__0_carry_i_14_n_0,n17__0_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__0_carry__0
       (.CI(n17__0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n17__0_carry__0_CO_UNCONNECTED[7:3],n17__0_carry__0_n_5,NLW_n17__0_carry__0_CO_UNCONNECTED[1],n17__0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n17__0_carry__0_i_1_n_0,n17__0_carry__0_i_2_n_0}),
        .O({NLW_n17__0_carry__0_O_UNCONNECTED[7:2],n17__0_carry__0_n_14,n17__0_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n17__0_carry__0_i_3_n_0,n17__0_carry__0_i_4_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__0_carry__0_i_1
       (.I0(n11_reg_n_46),
        .I1(n4[7]),
        .I2(n11_reg_n_45),
        .I3(n4[6]),
        .O(n17__0_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n17__0_carry__0_i_2
       (.I0(n11_reg_n_45),
        .I1(n4[5]),
        .I2(n11_reg_n_46),
        .I3(n4[6]),
        .I4(n11_reg_n_47),
        .I5(n4[7]),
        .O(n17__0_carry__0_i_2_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n17__0_carry__0_i_3
       (.I0(n4[6]),
        .I1(n11_reg_n_46),
        .I2(n11_reg_n_45),
        .I3(n4[7]),
        .O(n17__0_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n17__0_carry__0_i_4
       (.I0(n11_reg_n_47),
        .I1(n4[5]),
        .I2(n4[6]),
        .I3(n11_reg_n_45),
        .I4(n4[7]),
        .I5(n11_reg_n_46),
        .O(n17__0_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__0_carry_i_1
       (.I0(n11_reg_n_45),
        .I1(n4[4]),
        .I2(n11_reg_n_46),
        .I3(n4[5]),
        .I4(n11_reg_n_47),
        .I5(n4[6]),
        .O(n17__0_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__0_carry_i_10
       (.I0(n17__0_carry_i_3_n_0),
        .I1(n11_reg_n_46),
        .I2(n4[4]),
        .I3(n17__0_carry_i_18_n_0),
        .I4(n4[5]),
        .I5(n11_reg_n_47),
        .O(n17__0_carry_i_10_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__0_carry_i_11
       (.I0(n17__0_carry_i_4_n_0),
        .I1(n11_reg_n_46),
        .I2(n4[3]),
        .I3(n17__0_carry_i_19_n_0),
        .I4(n4[4]),
        .I5(n11_reg_n_47),
        .O(n17__0_carry_i_11_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n17__0_carry_i_12
       (.I0(n4[2]),
        .I1(n17__0_carry_i_20_n_0),
        .I2(n4[1]),
        .I3(n11_reg_n_46),
        .I4(n4[0]),
        .I5(n11_reg_n_45),
        .O(n17__0_carry_i_12_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n17__0_carry_i_13
       (.I0(n4[0]),
        .I1(n11_reg_n_45),
        .I2(n4[1]),
        .I3(n11_reg_n_46),
        .I4(n11_reg_n_47),
        .I5(n4[2]),
        .O(n17__0_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__0_carry_i_14
       (.I0(n11_reg_n_47),
        .I1(n4[1]),
        .I2(n11_reg_n_46),
        .I3(n4[0]),
        .O(n17__0_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__0_carry_i_15
       (.I0(n4[0]),
        .I1(n11_reg_n_47),
        .O(n17__0_carry_i_15_n_0));
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_16
       (.I0(n4[5]),
        .I1(n11_reg_n_45),
        .O(n17__0_carry_i_16_n_0));
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_17
       (.I0(n4[4]),
        .I1(n11_reg_n_45),
        .O(n17__0_carry_i_17_n_0));
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_18
       (.I0(n4[3]),
        .I1(n11_reg_n_45),
        .O(n17__0_carry_i_18_n_0));
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_19
       (.I0(n4[2]),
        .I1(n11_reg_n_45),
        .O(n17__0_carry_i_19_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__0_carry_i_2
       (.I0(n11_reg_n_45),
        .I1(n4[3]),
        .I2(n11_reg_n_46),
        .I3(n4[4]),
        .I4(n11_reg_n_47),
        .I5(n4[5]),
        .O(n17__0_carry_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__0_carry_i_20
       (.I0(n4[3]),
        .I1(n11_reg_n_47),
        .O(n17__0_carry_i_20_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__0_carry_i_3
       (.I0(n11_reg_n_45),
        .I1(n4[2]),
        .I2(n11_reg_n_46),
        .I3(n4[3]),
        .I4(n11_reg_n_47),
        .I5(n4[4]),
        .O(n17__0_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__0_carry_i_4
       (.I0(n11_reg_n_45),
        .I1(n4[1]),
        .I2(n11_reg_n_46),
        .I3(n4[2]),
        .I4(n11_reg_n_47),
        .I5(n4[3]),
        .O(n17__0_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n17__0_carry_i_5
       (.I0(n11_reg_n_46),
        .I1(n4[2]),
        .I2(n11_reg_n_45),
        .I3(n4[1]),
        .I4(n4[3]),
        .I5(n11_reg_n_47),
        .O(n17__0_carry_i_5_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__0_carry_i_6
       (.I0(n11_reg_n_46),
        .I1(n4[1]),
        .I2(n11_reg_n_45),
        .I3(n4[0]),
        .O(n17__0_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__0_carry_i_7
       (.I0(n11_reg_n_47),
        .I1(n4[1]),
        .O(n17__0_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n17__0_carry_i_8
       (.I0(n17__0_carry_i_1_n_0),
        .I1(n11_reg_n_46),
        .I2(n4[6]),
        .I3(n17__0_carry_i_16_n_0),
        .I4(n4[7]),
        .I5(n11_reg_n_47),
        .O(n17__0_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__0_carry_i_9
       (.I0(n17__0_carry_i_2_n_0),
        .I1(n11_reg_n_46),
        .I2(n4[5]),
        .I3(n17__0_carry_i_17_n_0),
        .I4(n4[6]),
        .I5(n11_reg_n_47),
        .O(n17__0_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__27_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n17__27_carry_n_0,n17__27_carry_n_1,n17__27_carry_n_2,n17__27_carry_n_3,n17__27_carry_n_4,n17__27_carry_n_5,n17__27_carry_n_6,n17__27_carry_n_7}),
        .DI({n17__27_carry_i_1_n_0,n17__27_carry_i_2_n_0,n17__27_carry_i_3_n_0,n17__27_carry_i_4_n_0,n17__27_carry_i_5_n_0,n17__27_carry_i_6_n_0,n17__27_carry_i_7_n_0,1'b0}),
        .O({n17__27_carry_n_8,n17__27_carry_n_9,n17__27_carry_n_10,n17__27_carry_n_11,n17__27_carry_n_12,n17__27_carry_n_13,n17__27_carry_n_14,n17__27_carry_n_15}),
        .S({n17__27_carry_i_8_n_0,n17__27_carry_i_9_n_0,n17__27_carry_i_10_n_0,n17__27_carry_i_11_n_0,n17__27_carry_i_12_n_0,n17__27_carry_i_13_n_0,n17__27_carry_i_14_n_0,n17__27_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__27_carry__0
       (.CI(n17__27_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n17__27_carry__0_CO_UNCONNECTED[7:3],n17__27_carry__0_n_5,NLW_n17__27_carry__0_CO_UNCONNECTED[1],n17__27_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n17__27_carry__0_i_1_n_0,n17__27_carry__0_i_2_n_0}),
        .O({NLW_n17__27_carry__0_O_UNCONNECTED[7:2],n17__27_carry__0_n_14,n17__27_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n17__27_carry__0_i_3_n_0,n17__27_carry__0_i_4_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__27_carry__0_i_1
       (.I0(n11_reg_n_43),
        .I1(n4[7]),
        .I2(n11_reg_n_42),
        .I3(n4[6]),
        .O(n17__27_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n17__27_carry__0_i_2
       (.I0(n11_reg_n_42),
        .I1(n4[5]),
        .I2(n11_reg_n_43),
        .I3(n4[6]),
        .I4(n11_reg_n_44),
        .I5(n4[7]),
        .O(n17__27_carry__0_i_2_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n17__27_carry__0_i_3
       (.I0(n4[6]),
        .I1(n11_reg_n_43),
        .I2(n11_reg_n_42),
        .I3(n4[7]),
        .O(n17__27_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n17__27_carry__0_i_4
       (.I0(n11_reg_n_44),
        .I1(n4[5]),
        .I2(n4[6]),
        .I3(n11_reg_n_42),
        .I4(n4[7]),
        .I5(n11_reg_n_43),
        .O(n17__27_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__27_carry_i_1
       (.I0(n11_reg_n_42),
        .I1(n4[4]),
        .I2(n11_reg_n_43),
        .I3(n4[5]),
        .I4(n11_reg_n_44),
        .I5(n4[6]),
        .O(n17__27_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__27_carry_i_10
       (.I0(n17__27_carry_i_3_n_0),
        .I1(n11_reg_n_43),
        .I2(n4[4]),
        .I3(n17__27_carry_i_18_n_0),
        .I4(n4[5]),
        .I5(n11_reg_n_44),
        .O(n17__27_carry_i_10_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__27_carry_i_11
       (.I0(n17__27_carry_i_4_n_0),
        .I1(n11_reg_n_43),
        .I2(n4[3]),
        .I3(n17__27_carry_i_19_n_0),
        .I4(n4[4]),
        .I5(n11_reg_n_44),
        .O(n17__27_carry_i_11_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n17__27_carry_i_12
       (.I0(n4[2]),
        .I1(n17__27_carry_i_20_n_0),
        .I2(n4[1]),
        .I3(n11_reg_n_43),
        .I4(n4[0]),
        .I5(n11_reg_n_42),
        .O(n17__27_carry_i_12_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n17__27_carry_i_13
       (.I0(n4[0]),
        .I1(n11_reg_n_42),
        .I2(n4[1]),
        .I3(n11_reg_n_43),
        .I4(n11_reg_n_44),
        .I5(n4[2]),
        .O(n17__27_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__27_carry_i_14
       (.I0(n11_reg_n_44),
        .I1(n4[1]),
        .I2(n11_reg_n_43),
        .I3(n4[0]),
        .O(n17__27_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__27_carry_i_15
       (.I0(n4[0]),
        .I1(n11_reg_n_44),
        .O(n17__27_carry_i_15_n_0));
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_16
       (.I0(n4[5]),
        .I1(n11_reg_n_42),
        .O(n17__27_carry_i_16_n_0));
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_17
       (.I0(n4[4]),
        .I1(n11_reg_n_42),
        .O(n17__27_carry_i_17_n_0));
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_18
       (.I0(n4[3]),
        .I1(n11_reg_n_42),
        .O(n17__27_carry_i_18_n_0));
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_19
       (.I0(n4[2]),
        .I1(n11_reg_n_42),
        .O(n17__27_carry_i_19_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__27_carry_i_2
       (.I0(n11_reg_n_42),
        .I1(n4[3]),
        .I2(n11_reg_n_43),
        .I3(n4[4]),
        .I4(n11_reg_n_44),
        .I5(n4[5]),
        .O(n17__27_carry_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n17__27_carry_i_20
       (.I0(n4[3]),
        .I1(n11_reg_n_44),
        .O(n17__27_carry_i_20_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__27_carry_i_3
       (.I0(n11_reg_n_42),
        .I1(n4[2]),
        .I2(n11_reg_n_43),
        .I3(n4[3]),
        .I4(n11_reg_n_44),
        .I5(n4[4]),
        .O(n17__27_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n17__27_carry_i_4
       (.I0(n11_reg_n_42),
        .I1(n4[1]),
        .I2(n11_reg_n_43),
        .I3(n4[2]),
        .I4(n11_reg_n_44),
        .I5(n4[3]),
        .O(n17__27_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n17__27_carry_i_5
       (.I0(n11_reg_n_43),
        .I1(n4[2]),
        .I2(n11_reg_n_42),
        .I3(n4[1]),
        .I4(n4[3]),
        .I5(n11_reg_n_44),
        .O(n17__27_carry_i_5_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__27_carry_i_6
       (.I0(n11_reg_n_43),
        .I1(n4[1]),
        .I2(n11_reg_n_42),
        .I3(n4[0]),
        .O(n17__27_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__27_carry_i_7
       (.I0(n11_reg_n_44),
        .I1(n4[1]),
        .O(n17__27_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n17__27_carry_i_8
       (.I0(n17__27_carry_i_1_n_0),
        .I1(n11_reg_n_43),
        .I2(n4[6]),
        .I3(n17__27_carry_i_16_n_0),
        .I4(n4[7]),
        .I5(n11_reg_n_44),
        .O(n17__27_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n17__27_carry_i_9
       (.I0(n17__27_carry_i_2_n_0),
        .I1(n11_reg_n_43),
        .I2(n4[5]),
        .I3(n17__27_carry_i_17_n_0),
        .I4(n4[6]),
        .I5(n11_reg_n_44),
        .O(n17__27_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__56_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n17__56_carry_n_0,n17__56_carry_n_1,n17__56_carry_n_2,n17__56_carry_n_3,n17__56_carry_n_4,n17__56_carry_n_5,n17__56_carry_n_6,n17__56_carry_n_7}),
        .DI({n17__56_carry_i_1_n_0,n17__56_carry_i_2_n_0,n17__56_carry_i_3_n_0,n17__56_carry_i_4_n_0,n17__56_carry_i_5_n_0,n17__56_carry_i_6_n_0,n17__56_carry_i_7_n_0,1'b0}),
        .O({n17__56_carry_n_8,n17__56_carry_n_9,n17__56_carry_n_10,n17__56_carry_n_11,n17__56_carry_n_12,n17__56_carry_n_13,n17__56_carry_n_14,n17__56_carry_n_15}),
        .S({n17__56_carry_i_8_n_0,n17__56_carry_i_9_n_0,n17__56_carry_i_10_n_0,n17__56_carry_i_11_n_0,n17__56_carry_i_12_n_0,n17__56_carry_i_13_n_0,n17__56_carry_i_14_n_0,n17__56_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__56_carry__0
       (.CI(n17__56_carry_n_0),
        .CI_TOP(1'b0),
        .CO(NLW_n17__56_carry__0_CO_UNCONNECTED[7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_n17__56_carry__0_O_UNCONNECTED[7:1],n17__56_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n17__56_carry__0_i_1_n_0}));
  LUT4 #(
    .INIT(16'hE53F)) 
    n17__56_carry__0_i_1
       (.I0(n11_reg_n_41),
        .I1(n4[6]),
        .I2(n11_reg_n_40),
        .I3(n4[7]),
        .O(n17__56_carry__0_i_1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__56_carry_i_1
       (.I0(n11_reg_n_40),
        .I1(n4[5]),
        .I2(n11_reg_n_41),
        .I3(n4[6]),
        .O(n17__56_carry_i_1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n17__56_carry_i_10
       (.I0(n4[3]),
        .I1(n4[4]),
        .I2(n11_reg_n_40),
        .I3(n4[5]),
        .I4(n11_reg_n_41),
        .O(n17__56_carry_i_10_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n17__56_carry_i_11
       (.I0(n4[2]),
        .I1(n4[3]),
        .I2(n11_reg_n_40),
        .I3(n4[4]),
        .I4(n11_reg_n_41),
        .O(n17__56_carry_i_11_n_0));
  LUT5 #(
    .INIT(32'h9F606060)) 
    n17__56_carry_i_12
       (.I0(n4[1]),
        .I1(n4[2]),
        .I2(n11_reg_n_40),
        .I3(n4[3]),
        .I4(n11_reg_n_41),
        .O(n17__56_carry_i_12_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n17__56_carry_i_13
       (.I0(n11_reg_n_40),
        .I1(n4[1]),
        .I2(n11_reg_n_41),
        .I3(n4[2]),
        .O(n17__56_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h8777)) 
    n17__56_carry_i_14
       (.I0(n11_reg_n_40),
        .I1(n4[0]),
        .I2(n11_reg_n_41),
        .I3(n4[1]),
        .O(n17__56_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__56_carry_i_15
       (.I0(n4[0]),
        .I1(n11_reg_n_41),
        .O(n17__56_carry_i_15_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__56_carry_i_2
       (.I0(n11_reg_n_40),
        .I1(n4[4]),
        .I2(n11_reg_n_41),
        .I3(n4[5]),
        .O(n17__56_carry_i_2_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__56_carry_i_3
       (.I0(n11_reg_n_40),
        .I1(n4[3]),
        .I2(n11_reg_n_41),
        .I3(n4[4]),
        .O(n17__56_carry_i_3_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n17__56_carry_i_4
       (.I0(n11_reg_n_40),
        .I1(n4[2]),
        .I2(n11_reg_n_41),
        .I3(n4[3]),
        .O(n17__56_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n17__56_carry_i_5
       (.I0(n4[1]),
        .I1(n11_reg_n_40),
        .O(n17__56_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__56_carry_i_6
       (.I0(n11_reg_n_40),
        .I1(n4[1]),
        .O(n17__56_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n17__56_carry_i_7
       (.I0(n4[0]),
        .I1(n11_reg_n_40),
        .O(n17__56_carry_i_7_n_0));
  LUT5 #(
    .INIT(32'h738CC0C0)) 
    n17__56_carry_i_8
       (.I0(n4[5]),
        .I1(n4[6]),
        .I2(n11_reg_n_40),
        .I3(n4[7]),
        .I4(n11_reg_n_41),
        .O(n17__56_carry_i_8_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n17__56_carry_i_9
       (.I0(n4[4]),
        .I1(n4[5]),
        .I2(n11_reg_n_40),
        .I3(n4[6]),
        .I4(n11_reg_n_41),
        .O(n17__56_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__81_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n17__81_carry_n_0,n17__81_carry_n_1,n17__81_carry_n_2,n17__81_carry_n_3,n17__81_carry_n_4,n17__81_carry_n_5,n17__81_carry_n_6,n17__81_carry_n_7}),
        .DI({n17__81_carry_i_1_n_0,n17__81_carry_i_2_n_0,n17__81_carry_i_3_n_0,n17__81_carry_i_4_n_0,n17__81_carry_i_5_n_0,n17__81_carry_i_6_n_0,n17__81_carry_i_7_n_0,1'b0}),
        .O({n17[10:7],NLW_n17__81_carry_O_UNCONNECTED[3:0]}),
        .S({n17__81_carry_i_8_n_0,n17__81_carry_i_9_n_0,n17__81_carry_i_10_n_0,n17__81_carry_i_11_n_0,n17__81_carry_i_12_n_0,n17__81_carry_i_13_n_0,n17__81_carry_i_14_n_0,n17__81_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n17__81_carry__0
       (.CI(n17__81_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n17__81_carry__0_CO_UNCONNECTED[7:3],n17__81_carry__0_n_5,n17__81_carry__0_n_6,n17__81_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n17__81_carry__0_i_1_n_0,n17__81_carry__0_i_2_n_0,n17__81_carry__0_i_3_n_0}),
        .O({NLW_n17__81_carry__0_O_UNCONNECTED[7:4],n17[14:11]}),
        .S({1'b0,1'b0,1'b0,1'b0,n17__81_carry__0_i_4_n_0,n17__81_carry__0_i_5_n_0,n17__81_carry__0_i_6_n_0,n17__81_carry__0_i_7_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry__0_i_1
       (.I0(n17__27_carry__0_n_14),
        .I1(n17__56_carry_n_9),
        .O(n17__81_carry__0_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry__0_i_2
       (.I0(n17__27_carry__0_n_15),
        .I1(n17__56_carry_n_10),
        .O(n17__81_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry__0_i_3
       (.I0(n17__56_carry_n_11),
        .I1(n17__27_carry_n_8),
        .I2(n17__0_carry__0_n_5),
        .O(n17__81_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n17__81_carry__0_i_4
       (.I0(n17__27_carry__0_n_5),
        .I1(n17__56_carry_n_8),
        .I2(n17__56_carry__0_n_15),
        .O(n17__81_carry__0_i_4_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n17__81_carry__0_i_5
       (.I0(n17__27_carry__0_n_14),
        .I1(n17__56_carry_n_9),
        .I2(n17__56_carry_n_8),
        .I3(n17__27_carry__0_n_5),
        .O(n17__81_carry__0_i_5_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n17__81_carry__0_i_6
       (.I0(n17__27_carry__0_n_15),
        .I1(n17__56_carry_n_10),
        .I2(n17__56_carry_n_9),
        .I3(n17__27_carry__0_n_14),
        .O(n17__81_carry__0_i_6_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n17__81_carry__0_i_7
       (.I0(n17__0_carry__0_n_5),
        .I1(n17__27_carry_n_8),
        .I2(n17__56_carry_n_11),
        .I3(n17__56_carry_n_10),
        .I4(n17__27_carry__0_n_15),
        .O(n17__81_carry__0_i_7_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry_i_1
       (.I0(n17__56_carry_n_12),
        .I1(n17__27_carry_n_9),
        .I2(n17__0_carry__0_n_14),
        .O(n17__81_carry_i_1_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_10
       (.I0(n17__56_carry_n_13),
        .I1(n17__27_carry_n_10),
        .I2(n17__0_carry__0_n_15),
        .I3(n17__81_carry_i_3_n_0),
        .O(n17__81_carry_i_10_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_11
       (.I0(n17__56_carry_n_14),
        .I1(n17__27_carry_n_11),
        .I2(n17__0_carry_n_8),
        .I3(n17__81_carry_i_4_n_0),
        .O(n17__81_carry_i_11_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_12
       (.I0(n17__56_carry_n_15),
        .I1(n17__27_carry_n_12),
        .I2(n17__0_carry_n_9),
        .I3(n17__81_carry_i_5_n_0),
        .O(n17__81_carry_i_12_n_0));
  LUT4 #(
    .INIT(16'h9666)) 
    n17__81_carry_i_13
       (.I0(n17__27_carry_n_13),
        .I1(n17__0_carry_n_10),
        .I2(n17__0_carry_n_11),
        .I3(n17__27_carry_n_14),
        .O(n17__81_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n17__81_carry_i_14
       (.I0(n17__0_carry_n_12),
        .I1(n17__27_carry_n_15),
        .I2(n17__27_carry_n_14),
        .I3(n17__0_carry_n_11),
        .O(n17__81_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n17__81_carry_i_15
       (.I0(n17__0_carry_n_12),
        .I1(n17__27_carry_n_15),
        .O(n17__81_carry_i_15_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry_i_2
       (.I0(n17__56_carry_n_13),
        .I1(n17__27_carry_n_10),
        .I2(n17__0_carry__0_n_15),
        .O(n17__81_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry_i_3
       (.I0(n17__56_carry_n_14),
        .I1(n17__27_carry_n_11),
        .I2(n17__0_carry_n_8),
        .O(n17__81_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n17__81_carry_i_4
       (.I0(n17__56_carry_n_15),
        .I1(n17__27_carry_n_12),
        .I2(n17__0_carry_n_9),
        .O(n17__81_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry_i_5
       (.I0(n17__27_carry_n_13),
        .I1(n17__0_carry_n_10),
        .O(n17__81_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry_i_6
       (.I0(n17__0_carry_n_11),
        .I1(n17__27_carry_n_14),
        .O(n17__81_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n17__81_carry_i_7
       (.I0(n17__0_carry_n_12),
        .I1(n17__27_carry_n_15),
        .O(n17__81_carry_i_7_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_8
       (.I0(n17__81_carry_i_1_n_0),
        .I1(n17__27_carry_n_8),
        .I2(n17__56_carry_n_11),
        .I3(n17__0_carry__0_n_5),
        .O(n17__81_carry_i_8_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n17__81_carry_i_9
       (.I0(n17__56_carry_n_12),
        .I1(n17__27_carry_n_9),
        .I2(n17__0_carry__0_n_14),
        .I3(n17__81_carry_i_2_n_0),
        .O(n17__81_carry_i_9_n_0));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[14]),
        .Q(n19_reg_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__0
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[13]),
        .Q(n19_reg__0_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__1
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[12]),
        .Q(n19_reg__1_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__2
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[11]),
        .Q(n19_reg__2_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__3
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[10]),
        .Q(n19_reg__3_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__4
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[9]),
        .Q(n19_reg__4_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__5
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[8]),
        .Q(n19_reg__5_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n19_reg__6
       (.C(clk_i),
        .CE(enable_i),
        .D(n17[7]),
        .Q(n19_reg__6_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[0]),
        .Q(\n1_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[10]),
        .Q(n2[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[11]),
        .Q(n2[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[12]),
        .Q(n2[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[13]),
        .Q(n2[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[14]),
        .Q(n2[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[15]),
        .Q(n2[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[1]),
        .Q(\n1_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[2]),
        .Q(\n1_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[3]),
        .Q(\n1_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[4]),
        .Q(\n1_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[5]),
        .Q(\n1_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[6]),
        .Q(\n1_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[7]),
        .Q(\n1_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[8]),
        .Q(n2[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[9]),
        .Q(n2[1]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n20_carry
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({NLW_n20_carry_CO_UNCONNECTED[7],n20_carry_n_1,n20_carry_n_2,n20_carry_n_3,n20_carry_n_4,n20_carry_n_5,n20_carry_n_6,n20_carry_n_7}),
        .DI({1'b0,\n16_reg_n_0_[6] ,\n16_reg_n_0_[5] ,\n16_reg_n_0_[4] ,\n16_reg_n_0_[3] ,\n16_reg_n_0_[2] ,\n16_reg_n_0_[1] ,\n16_reg_n_0_[0] }),
        .O(n202_out),
        .S({n20_carry_i_1__0_n_0,n20_carry_i_2__0_n_0,n20_carry_i_3__0_n_0,n20_carry_i_4__0_n_0,n20_carry_i_5__0_n_0,n20_carry_i_6__0_n_0,n20_carry_i_7__0_n_0,n20_carry_i_8__0_n_0}));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_1__0
       (.I0(\n16_reg_n_0_[7] ),
        .I1(n19_reg_n_0),
        .O(n20_carry_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_2__0
       (.I0(\n16_reg_n_0_[6] ),
        .I1(n19_reg__0_n_0),
        .O(n20_carry_i_2__0_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_3__0
       (.I0(\n16_reg_n_0_[5] ),
        .I1(n19_reg__1_n_0),
        .O(n20_carry_i_3__0_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_4__0
       (.I0(\n16_reg_n_0_[4] ),
        .I1(n19_reg__2_n_0),
        .O(n20_carry_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_5__0
       (.I0(\n16_reg_n_0_[3] ),
        .I1(n19_reg__3_n_0),
        .O(n20_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_6__0
       (.I0(\n16_reg_n_0_[2] ),
        .I1(n19_reg__4_n_0),
        .O(n20_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_7__0
       (.I0(\n16_reg_n_0_[1] ),
        .I1(n19_reg__5_n_0),
        .O(n20_carry_i_7__0_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    n20_carry_i_8__0
       (.I0(\n16_reg_n_0_[0] ),
        .I1(n19_reg__6_n_0),
        .O(n20_carry_i_8__0_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[0]),
        .Q(n21[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[1]),
        .Q(n21[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[2]),
        .Q(n21[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[3]),
        .Q(n21[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[4]),
        .Q(n21[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[5]),
        .Q(n21[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[6]),
        .Q(n21[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[7]),
        .Q(n21[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[15]),
        .Q(n22_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__0
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[14]),
        .Q(n22__0_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__0_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n22__0_carry_n_0,n22__0_carry_n_1,n22__0_carry_n_2,n22__0_carry_n_3,n22__0_carry_n_4,n22__0_carry_n_5,n22__0_carry_n_6,n22__0_carry_n_7}),
        .DI({n22__0_carry_i_1_n_0,n22__0_carry_i_2_n_0,n22__0_carry_i_3_n_0,n22__0_carry_i_4_n_0,n22__0_carry_i_5_n_0,n22__0_carry_i_6_n_0,n22__0_carry_i_7_n_0,1'b0}),
        .O({n22__0_carry_n_8,n22__0_carry_n_9,n22__0_carry_n_10,n22__0_carry_n_11,n22__0_carry_n_12,NLW_n22__0_carry_O_UNCONNECTED[2:0]}),
        .S({n22__0_carry_i_8_n_0,n22__0_carry_i_9_n_0,n22__0_carry_i_10_n_0,n22__0_carry_i_11_n_0,n22__0_carry_i_12_n_0,n22__0_carry_i_13_n_0,n22__0_carry_i_14_n_0,n22__0_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__0_carry__0
       (.CI(n22__0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n22__0_carry__0_CO_UNCONNECTED[7:3],n22__0_carry__0_n_5,NLW_n22__0_carry__0_CO_UNCONNECTED[1],n22__0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n22__0_carry__0_i_1_n_0,n22__0_carry__0_i_2_n_0}),
        .O({NLW_n22__0_carry__0_O_UNCONNECTED[7:2],n22__0_carry__0_n_14,n22__0_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n22__0_carry__0_i_3_n_0,n22__0_carry__0_i_4_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__0_carry__0_i_1
       (.I0(n11_reg_n_46),
        .I1(n22_n_0),
        .I2(n11_reg_n_45),
        .I3(n22__0_n_0),
        .O(n22__0_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n22__0_carry__0_i_2
       (.I0(n11_reg_n_45),
        .I1(n22__1_n_0),
        .I2(n11_reg_n_46),
        .I3(n22__0_n_0),
        .I4(n11_reg_n_47),
        .I5(n22_n_0),
        .O(n22__0_carry__0_i_2_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n22__0_carry__0_i_3
       (.I0(n22__0_n_0),
        .I1(n11_reg_n_46),
        .I2(n11_reg_n_45),
        .I3(n22_n_0),
        .O(n22__0_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n22__0_carry__0_i_4
       (.I0(n11_reg_n_47),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(n11_reg_n_45),
        .I4(n22_n_0),
        .I5(n11_reg_n_46),
        .O(n22__0_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__0_carry_i_1
       (.I0(n11_reg_n_45),
        .I1(n22__2_n_0),
        .I2(n11_reg_n_46),
        .I3(n22__1_n_0),
        .I4(n11_reg_n_47),
        .I5(n22__0_n_0),
        .O(n22__0_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__0_carry_i_10
       (.I0(n22__0_carry_i_3_n_0),
        .I1(n11_reg_n_46),
        .I2(n22__2_n_0),
        .I3(n22__0_carry_i_18_n_0),
        .I4(n22__1_n_0),
        .I5(n11_reg_n_47),
        .O(n22__0_carry_i_10_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__0_carry_i_11
       (.I0(n22__0_carry_i_4_n_0),
        .I1(n11_reg_n_46),
        .I2(n22__3_n_0),
        .I3(n22__0_carry_i_19_n_0),
        .I4(n22__2_n_0),
        .I5(n11_reg_n_47),
        .O(n22__0_carry_i_11_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n22__0_carry_i_12
       (.I0(n22__4_n_0),
        .I1(n22__0_carry_i_20_n_0),
        .I2(n22__5_n_0),
        .I3(n11_reg_n_46),
        .I4(n22__6_n_0),
        .I5(n11_reg_n_45),
        .O(n22__0_carry_i_12_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n22__0_carry_i_13
       (.I0(n22__6_n_0),
        .I1(n11_reg_n_45),
        .I2(n22__5_n_0),
        .I3(n11_reg_n_46),
        .I4(n11_reg_n_47),
        .I5(n22__4_n_0),
        .O(n22__0_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__0_carry_i_14
       (.I0(n11_reg_n_47),
        .I1(n22__5_n_0),
        .I2(n11_reg_n_46),
        .I3(n22__6_n_0),
        .O(n22__0_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__0_carry_i_15
       (.I0(n22__6_n_0),
        .I1(n11_reg_n_47),
        .O(n22__0_carry_i_15_n_0));
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_16
       (.I0(n22__1_n_0),
        .I1(n11_reg_n_45),
        .O(n22__0_carry_i_16_n_0));
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_17
       (.I0(n22__2_n_0),
        .I1(n11_reg_n_45),
        .O(n22__0_carry_i_17_n_0));
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_18
       (.I0(n22__3_n_0),
        .I1(n11_reg_n_45),
        .O(n22__0_carry_i_18_n_0));
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_19
       (.I0(n22__4_n_0),
        .I1(n11_reg_n_45),
        .O(n22__0_carry_i_19_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__0_carry_i_2
       (.I0(n11_reg_n_45),
        .I1(n22__3_n_0),
        .I2(n11_reg_n_46),
        .I3(n22__2_n_0),
        .I4(n11_reg_n_47),
        .I5(n22__1_n_0),
        .O(n22__0_carry_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__0_carry_i_20
       (.I0(n22__3_n_0),
        .I1(n11_reg_n_47),
        .O(n22__0_carry_i_20_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__0_carry_i_3
       (.I0(n11_reg_n_45),
        .I1(n22__4_n_0),
        .I2(n11_reg_n_46),
        .I3(n22__3_n_0),
        .I4(n11_reg_n_47),
        .I5(n22__2_n_0),
        .O(n22__0_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__0_carry_i_4
       (.I0(n11_reg_n_45),
        .I1(n22__5_n_0),
        .I2(n11_reg_n_46),
        .I3(n22__4_n_0),
        .I4(n11_reg_n_47),
        .I5(n22__3_n_0),
        .O(n22__0_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n22__0_carry_i_5
       (.I0(n11_reg_n_46),
        .I1(n22__4_n_0),
        .I2(n11_reg_n_45),
        .I3(n22__5_n_0),
        .I4(n22__3_n_0),
        .I5(n11_reg_n_47),
        .O(n22__0_carry_i_5_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__0_carry_i_6
       (.I0(n11_reg_n_46),
        .I1(n22__5_n_0),
        .I2(n11_reg_n_45),
        .I3(n22__6_n_0),
        .O(n22__0_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__0_carry_i_7
       (.I0(n11_reg_n_47),
        .I1(n22__5_n_0),
        .O(n22__0_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n22__0_carry_i_8
       (.I0(n22__0_carry_i_1_n_0),
        .I1(n11_reg_n_46),
        .I2(n22__0_n_0),
        .I3(n22__0_carry_i_16_n_0),
        .I4(n22_n_0),
        .I5(n11_reg_n_47),
        .O(n22__0_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__0_carry_i_9
       (.I0(n22__0_carry_i_2_n_0),
        .I1(n11_reg_n_46),
        .I2(n22__1_n_0),
        .I3(n22__0_carry_i_17_n_0),
        .I4(n22__0_n_0),
        .I5(n11_reg_n_47),
        .O(n22__0_carry_i_9_n_0));
  FDRE #(
    .INIT(1'b0)) 
    n22__1
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[13]),
        .Q(n22__1_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__2
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[12]),
        .Q(n22__2_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__27_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n22__27_carry_n_0,n22__27_carry_n_1,n22__27_carry_n_2,n22__27_carry_n_3,n22__27_carry_n_4,n22__27_carry_n_5,n22__27_carry_n_6,n22__27_carry_n_7}),
        .DI({n22__27_carry_i_1_n_0,n22__27_carry_i_2_n_0,n22__27_carry_i_3_n_0,n22__27_carry_i_4_n_0,n22__27_carry_i_5_n_0,n22__27_carry_i_6_n_0,n22__27_carry_i_7_n_0,1'b0}),
        .O({n22__27_carry_n_8,n22__27_carry_n_9,n22__27_carry_n_10,n22__27_carry_n_11,n22__27_carry_n_12,n22__27_carry_n_13,n22__27_carry_n_14,n22__27_carry_n_15}),
        .S({n22__27_carry_i_8_n_0,n22__27_carry_i_9_n_0,n22__27_carry_i_10_n_0,n22__27_carry_i_11_n_0,n22__27_carry_i_12_n_0,n22__27_carry_i_13_n_0,n22__27_carry_i_14_n_0,n22__27_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__27_carry__0
       (.CI(n22__27_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n22__27_carry__0_CO_UNCONNECTED[7:3],n22__27_carry__0_n_5,NLW_n22__27_carry__0_CO_UNCONNECTED[1],n22__27_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n22__27_carry__0_i_1_n_0,n22__27_carry__0_i_2_n_0}),
        .O({NLW_n22__27_carry__0_O_UNCONNECTED[7:2],n22__27_carry__0_n_14,n22__27_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n22__27_carry__0_i_3_n_0,n22__27_carry__0_i_4_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__27_carry__0_i_1
       (.I0(n11_reg_n_43),
        .I1(n22_n_0),
        .I2(n11_reg_n_42),
        .I3(n22__0_n_0),
        .O(n22__27_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n22__27_carry__0_i_2
       (.I0(n11_reg_n_42),
        .I1(n22__1_n_0),
        .I2(n11_reg_n_43),
        .I3(n22__0_n_0),
        .I4(n11_reg_n_44),
        .I5(n22_n_0),
        .O(n22__27_carry__0_i_2_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n22__27_carry__0_i_3
       (.I0(n22__0_n_0),
        .I1(n11_reg_n_43),
        .I2(n11_reg_n_42),
        .I3(n22_n_0),
        .O(n22__27_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n22__27_carry__0_i_4
       (.I0(n11_reg_n_44),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(n11_reg_n_42),
        .I4(n22_n_0),
        .I5(n11_reg_n_43),
        .O(n22__27_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__27_carry_i_1
       (.I0(n11_reg_n_42),
        .I1(n22__2_n_0),
        .I2(n11_reg_n_43),
        .I3(n22__1_n_0),
        .I4(n11_reg_n_44),
        .I5(n22__0_n_0),
        .O(n22__27_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__27_carry_i_10
       (.I0(n22__27_carry_i_3_n_0),
        .I1(n11_reg_n_43),
        .I2(n22__2_n_0),
        .I3(n22__27_carry_i_18_n_0),
        .I4(n22__1_n_0),
        .I5(n11_reg_n_44),
        .O(n22__27_carry_i_10_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__27_carry_i_11
       (.I0(n22__27_carry_i_4_n_0),
        .I1(n11_reg_n_43),
        .I2(n22__3_n_0),
        .I3(n22__27_carry_i_19_n_0),
        .I4(n22__2_n_0),
        .I5(n11_reg_n_44),
        .O(n22__27_carry_i_11_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n22__27_carry_i_12
       (.I0(n22__4_n_0),
        .I1(n22__27_carry_i_20_n_0),
        .I2(n22__5_n_0),
        .I3(n11_reg_n_43),
        .I4(n22__6_n_0),
        .I5(n11_reg_n_42),
        .O(n22__27_carry_i_12_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n22__27_carry_i_13
       (.I0(n22__6_n_0),
        .I1(n11_reg_n_42),
        .I2(n22__5_n_0),
        .I3(n11_reg_n_43),
        .I4(n11_reg_n_44),
        .I5(n22__4_n_0),
        .O(n22__27_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__27_carry_i_14
       (.I0(n11_reg_n_44),
        .I1(n22__5_n_0),
        .I2(n11_reg_n_43),
        .I3(n22__6_n_0),
        .O(n22__27_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__27_carry_i_15
       (.I0(n22__6_n_0),
        .I1(n11_reg_n_44),
        .O(n22__27_carry_i_15_n_0));
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_16
       (.I0(n22__1_n_0),
        .I1(n11_reg_n_42),
        .O(n22__27_carry_i_16_n_0));
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_17
       (.I0(n22__2_n_0),
        .I1(n11_reg_n_42),
        .O(n22__27_carry_i_17_n_0));
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_18
       (.I0(n22__3_n_0),
        .I1(n11_reg_n_42),
        .O(n22__27_carry_i_18_n_0));
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_19
       (.I0(n22__4_n_0),
        .I1(n11_reg_n_42),
        .O(n22__27_carry_i_19_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__27_carry_i_2
       (.I0(n11_reg_n_42),
        .I1(n22__3_n_0),
        .I2(n11_reg_n_43),
        .I3(n22__2_n_0),
        .I4(n11_reg_n_44),
        .I5(n22__1_n_0),
        .O(n22__27_carry_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n22__27_carry_i_20
       (.I0(n22__3_n_0),
        .I1(n11_reg_n_44),
        .O(n22__27_carry_i_20_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__27_carry_i_3
       (.I0(n11_reg_n_42),
        .I1(n22__4_n_0),
        .I2(n11_reg_n_43),
        .I3(n22__3_n_0),
        .I4(n11_reg_n_44),
        .I5(n22__2_n_0),
        .O(n22__27_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n22__27_carry_i_4
       (.I0(n11_reg_n_42),
        .I1(n22__5_n_0),
        .I2(n11_reg_n_43),
        .I3(n22__4_n_0),
        .I4(n11_reg_n_44),
        .I5(n22__3_n_0),
        .O(n22__27_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n22__27_carry_i_5
       (.I0(n11_reg_n_43),
        .I1(n22__4_n_0),
        .I2(n11_reg_n_42),
        .I3(n22__5_n_0),
        .I4(n22__3_n_0),
        .I5(n11_reg_n_44),
        .O(n22__27_carry_i_5_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__27_carry_i_6
       (.I0(n11_reg_n_43),
        .I1(n22__5_n_0),
        .I2(n11_reg_n_42),
        .I3(n22__6_n_0),
        .O(n22__27_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__27_carry_i_7
       (.I0(n11_reg_n_44),
        .I1(n22__5_n_0),
        .O(n22__27_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n22__27_carry_i_8
       (.I0(n22__27_carry_i_1_n_0),
        .I1(n11_reg_n_43),
        .I2(n22__0_n_0),
        .I3(n22__27_carry_i_16_n_0),
        .I4(n22_n_0),
        .I5(n11_reg_n_44),
        .O(n22__27_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n22__27_carry_i_9
       (.I0(n22__27_carry_i_2_n_0),
        .I1(n11_reg_n_43),
        .I2(n22__1_n_0),
        .I3(n22__27_carry_i_17_n_0),
        .I4(n22__0_n_0),
        .I5(n11_reg_n_44),
        .O(n22__27_carry_i_9_n_0));
  FDRE #(
    .INIT(1'b0)) 
    n22__3
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[11]),
        .Q(n22__3_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__4
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[10]),
        .Q(n22__4_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__5
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[9]),
        .Q(n22__5_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__56_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n22__56_carry_n_0,n22__56_carry_n_1,n22__56_carry_n_2,n22__56_carry_n_3,n22__56_carry_n_4,n22__56_carry_n_5,n22__56_carry_n_6,n22__56_carry_n_7}),
        .DI({n22__56_carry_i_1_n_0,n22__56_carry_i_2_n_0,n22__56_carry_i_3_n_0,n22__56_carry_i_4_n_0,n22__56_carry_i_5_n_0,n22__56_carry_i_6_n_0,n22__56_carry_i_7_n_0,1'b0}),
        .O({n22__56_carry_n_8,n22__56_carry_n_9,n22__56_carry_n_10,n22__56_carry_n_11,n22__56_carry_n_12,n22__56_carry_n_13,n22__56_carry_n_14,n22__56_carry_n_15}),
        .S({n22__56_carry_i_8_n_0,n22__56_carry_i_9_n_0,n22__56_carry_i_10_n_0,n22__56_carry_i_11_n_0,n22__56_carry_i_12_n_0,n22__56_carry_i_13_n_0,n22__56_carry_i_14_n_0,n22__56_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__56_carry__0
       (.CI(n22__56_carry_n_0),
        .CI_TOP(1'b0),
        .CO(NLW_n22__56_carry__0_CO_UNCONNECTED[7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_n22__56_carry__0_O_UNCONNECTED[7:1],n22__56_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n22__56_carry__0_i_1_n_0}));
  LUT4 #(
    .INIT(16'hE53F)) 
    n22__56_carry__0_i_1
       (.I0(n11_reg_n_41),
        .I1(n22__0_n_0),
        .I2(n11_reg_n_40),
        .I3(n22_n_0),
        .O(n22__56_carry__0_i_1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__56_carry_i_1
       (.I0(n11_reg_n_40),
        .I1(n22__1_n_0),
        .I2(n11_reg_n_41),
        .I3(n22__0_n_0),
        .O(n22__56_carry_i_1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n22__56_carry_i_10
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(n11_reg_n_40),
        .I3(n22__1_n_0),
        .I4(n11_reg_n_41),
        .O(n22__56_carry_i_10_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n22__56_carry_i_11
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n11_reg_n_40),
        .I3(n22__2_n_0),
        .I4(n11_reg_n_41),
        .O(n22__56_carry_i_11_n_0));
  LUT5 #(
    .INIT(32'h9F606060)) 
    n22__56_carry_i_12
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(n11_reg_n_40),
        .I3(n22__3_n_0),
        .I4(n11_reg_n_41),
        .O(n22__56_carry_i_12_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n22__56_carry_i_13
       (.I0(n11_reg_n_40),
        .I1(n22__5_n_0),
        .I2(n11_reg_n_41),
        .I3(n22__4_n_0),
        .O(n22__56_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h8777)) 
    n22__56_carry_i_14
       (.I0(n11_reg_n_40),
        .I1(n22__6_n_0),
        .I2(n11_reg_n_41),
        .I3(n22__5_n_0),
        .O(n22__56_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__56_carry_i_15
       (.I0(n22__6_n_0),
        .I1(n11_reg_n_41),
        .O(n22__56_carry_i_15_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__56_carry_i_2
       (.I0(n11_reg_n_40),
        .I1(n22__2_n_0),
        .I2(n11_reg_n_41),
        .I3(n22__1_n_0),
        .O(n22__56_carry_i_2_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__56_carry_i_3
       (.I0(n11_reg_n_40),
        .I1(n22__3_n_0),
        .I2(n11_reg_n_41),
        .I3(n22__2_n_0),
        .O(n22__56_carry_i_3_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n22__56_carry_i_4
       (.I0(n11_reg_n_40),
        .I1(n22__4_n_0),
        .I2(n11_reg_n_41),
        .I3(n22__3_n_0),
        .O(n22__56_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n22__56_carry_i_5
       (.I0(n22__5_n_0),
        .I1(n11_reg_n_40),
        .O(n22__56_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__56_carry_i_6
       (.I0(n11_reg_n_40),
        .I1(n22__5_n_0),
        .O(n22__56_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n22__56_carry_i_7
       (.I0(n22__6_n_0),
        .I1(n11_reg_n_40),
        .O(n22__56_carry_i_7_n_0));
  LUT5 #(
    .INIT(32'h738CC0C0)) 
    n22__56_carry_i_8
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n11_reg_n_40),
        .I3(n22_n_0),
        .I4(n11_reg_n_41),
        .O(n22__56_carry_i_8_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n22__56_carry_i_9
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(n11_reg_n_40),
        .I3(n22__0_n_0),
        .I4(n11_reg_n_41),
        .O(n22__56_carry_i_9_n_0));
  FDRE #(
    .INIT(1'b0)) 
    n22__6
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[8]),
        .Q(n22__6_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__81_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n22__81_carry_n_0,n22__81_carry_n_1,n22__81_carry_n_2,n22__81_carry_n_3,n22__81_carry_n_4,n22__81_carry_n_5,n22__81_carry_n_6,n22__81_carry_n_7}),
        .DI({n22__81_carry_i_1_n_0,n22__81_carry_i_2_n_0,n22__81_carry_i_3_n_0,n22__81_carry_i_4_n_0,n22__81_carry_i_5_n_0,n22__81_carry_i_6_n_0,n22__81_carry_i_7_n_0,1'b0}),
        .O({n23[3:0],NLW_n22__81_carry_O_UNCONNECTED[3:0]}),
        .S({n22__81_carry_i_8_n_0,n22__81_carry_i_9_n_0,n22__81_carry_i_10_n_0,n22__81_carry_i_11_n_0,n22__81_carry_i_12_n_0,n22__81_carry_i_13_n_0,n22__81_carry_i_14_n_0,n22__81_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n22__81_carry__0
       (.CI(n22__81_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n22__81_carry__0_CO_UNCONNECTED[7:3],n22__81_carry__0_n_5,n22__81_carry__0_n_6,n22__81_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n22__81_carry__0_i_1_n_0,n22__81_carry__0_i_2_n_0,n22__81_carry__0_i_3_n_0}),
        .O({NLW_n22__81_carry__0_O_UNCONNECTED[7:4],n23[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n22__81_carry__0_i_4_n_0,n22__81_carry__0_i_5_n_0,n22__81_carry__0_i_6_n_0,n22__81_carry__0_i_7_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry__0_i_1
       (.I0(n22__27_carry__0_n_14),
        .I1(n22__56_carry_n_9),
        .O(n22__81_carry__0_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry__0_i_2
       (.I0(n22__27_carry__0_n_15),
        .I1(n22__56_carry_n_10),
        .O(n22__81_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry__0_i_3
       (.I0(n22__56_carry_n_11),
        .I1(n22__27_carry_n_8),
        .I2(n22__0_carry__0_n_5),
        .O(n22__81_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n22__81_carry__0_i_4
       (.I0(n22__27_carry__0_n_5),
        .I1(n22__56_carry_n_8),
        .I2(n22__56_carry__0_n_15),
        .O(n22__81_carry__0_i_4_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n22__81_carry__0_i_5
       (.I0(n22__27_carry__0_n_14),
        .I1(n22__56_carry_n_9),
        .I2(n22__56_carry_n_8),
        .I3(n22__27_carry__0_n_5),
        .O(n22__81_carry__0_i_5_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n22__81_carry__0_i_6
       (.I0(n22__27_carry__0_n_15),
        .I1(n22__56_carry_n_10),
        .I2(n22__56_carry_n_9),
        .I3(n22__27_carry__0_n_14),
        .O(n22__81_carry__0_i_6_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n22__81_carry__0_i_7
       (.I0(n22__0_carry__0_n_5),
        .I1(n22__27_carry_n_8),
        .I2(n22__56_carry_n_11),
        .I3(n22__56_carry_n_10),
        .I4(n22__27_carry__0_n_15),
        .O(n22__81_carry__0_i_7_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry_i_1
       (.I0(n22__56_carry_n_12),
        .I1(n22__27_carry_n_9),
        .I2(n22__0_carry__0_n_14),
        .O(n22__81_carry_i_1_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_10
       (.I0(n22__56_carry_n_13),
        .I1(n22__27_carry_n_10),
        .I2(n22__0_carry__0_n_15),
        .I3(n22__81_carry_i_3_n_0),
        .O(n22__81_carry_i_10_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_11
       (.I0(n22__56_carry_n_14),
        .I1(n22__27_carry_n_11),
        .I2(n22__0_carry_n_8),
        .I3(n22__81_carry_i_4_n_0),
        .O(n22__81_carry_i_11_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_12
       (.I0(n22__56_carry_n_15),
        .I1(n22__27_carry_n_12),
        .I2(n22__0_carry_n_9),
        .I3(n22__81_carry_i_5_n_0),
        .O(n22__81_carry_i_12_n_0));
  LUT4 #(
    .INIT(16'h9666)) 
    n22__81_carry_i_13
       (.I0(n22__27_carry_n_13),
        .I1(n22__0_carry_n_10),
        .I2(n22__0_carry_n_11),
        .I3(n22__27_carry_n_14),
        .O(n22__81_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n22__81_carry_i_14
       (.I0(n22__0_carry_n_12),
        .I1(n22__27_carry_n_15),
        .I2(n22__27_carry_n_14),
        .I3(n22__0_carry_n_11),
        .O(n22__81_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n22__81_carry_i_15
       (.I0(n22__0_carry_n_12),
        .I1(n22__27_carry_n_15),
        .O(n22__81_carry_i_15_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry_i_2
       (.I0(n22__56_carry_n_13),
        .I1(n22__27_carry_n_10),
        .I2(n22__0_carry__0_n_15),
        .O(n22__81_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry_i_3
       (.I0(n22__56_carry_n_14),
        .I1(n22__27_carry_n_11),
        .I2(n22__0_carry_n_8),
        .O(n22__81_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n22__81_carry_i_4
       (.I0(n22__56_carry_n_15),
        .I1(n22__27_carry_n_12),
        .I2(n22__0_carry_n_9),
        .O(n22__81_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry_i_5
       (.I0(n22__27_carry_n_13),
        .I1(n22__0_carry_n_10),
        .O(n22__81_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry_i_6
       (.I0(n22__0_carry_n_11),
        .I1(n22__27_carry_n_14),
        .O(n22__81_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n22__81_carry_i_7
       (.I0(n22__0_carry_n_12),
        .I1(n22__27_carry_n_15),
        .O(n22__81_carry_i_7_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_8
       (.I0(n22__81_carry_i_1_n_0),
        .I1(n22__27_carry_n_8),
        .I2(n22__56_carry_n_11),
        .I3(n22__0_carry__0_n_5),
        .O(n22__81_carry_i_8_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n22__81_carry_i_9
       (.I0(n22__56_carry_n_12),
        .I1(n22__27_carry_n_9),
        .I2(n22__0_carry__0_n_14),
        .I3(n22__81_carry_i_2_n_0),
        .O(n22__81_carry_i_9_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[0]),
        .Q(n24[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[1]),
        .Q(n24[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[2]),
        .Q(n24[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[3]),
        .Q(n24[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[4]),
        .Q(n24[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[5]),
        .Q(n24[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[6]),
        .Q(n24[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n24_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n23[7]),
        .Q(n24[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__0_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__0_carry_n_0,n25__0_carry_n_1,n25__0_carry_n_2,n25__0_carry_n_3,n25__0_carry_n_4,n25__0_carry_n_5,n25__0_carry_n_6,n25__0_carry_n_7}),
        .DI({n25__0_carry_i_1_n_0,n25__0_carry_i_2_n_0,n25__0_carry_i_3_n_0,n25__0_carry_i_4_n_0,n25__0_carry_i_5_n_0,n25__0_carry_i_6_n_0,n25__0_carry_i_7_n_0,1'b0}),
        .O({n25__0_carry_n_8,n25__0_carry_n_9,n25__0_carry_n_10,n25__0_carry_n_11,n25__0_carry_n_12,NLW_n25__0_carry_O_UNCONNECTED[2:0]}),
        .S({n25__0_carry_i_8_n_0,n25__0_carry_i_9_n_0,n25__0_carry_i_10_n_0,n25__0_carry_i_11_n_0,n25__0_carry_i_12_n_0,n25__0_carry_i_13_n_0,n25__0_carry_i_14_n_0,n25__0_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__0_carry__0
       (.CI(n25__0_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__0_carry__0_CO_UNCONNECTED[7:3],n25__0_carry__0_n_5,NLW_n25__0_carry__0_CO_UNCONNECTED[1],n25__0_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25__0_carry__0_i_1_n_0,n25__0_carry__0_i_2_n_0}),
        .O({NLW_n25__0_carry__0_O_UNCONNECTED[7:2],n25__0_carry__0_n_14,n25__0_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n25__0_carry__0_i_3_n_0,n25__0_carry__0_i_4_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__0_carry__0_i_1
       (.I0(B[1]),
        .I1(n4[7]),
        .I2(B[2]),
        .I3(n4[6]),
        .O(n25__0_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n25__0_carry__0_i_2
       (.I0(B[2]),
        .I1(n4[5]),
        .I2(B[1]),
        .I3(n4[6]),
        .I4(B[0]),
        .I5(n4[7]),
        .O(n25__0_carry__0_i_2_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n25__0_carry__0_i_3
       (.I0(n4[6]),
        .I1(B[1]),
        .I2(B[2]),
        .I3(n4[7]),
        .O(n25__0_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n25__0_carry__0_i_4
       (.I0(B[0]),
        .I1(n4[5]),
        .I2(n4[6]),
        .I3(B[2]),
        .I4(n4[7]),
        .I5(B[1]),
        .O(n25__0_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__0_carry_i_1
       (.I0(B[2]),
        .I1(n4[4]),
        .I2(B[1]),
        .I3(n4[5]),
        .I4(B[0]),
        .I5(n4[6]),
        .O(n25__0_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__0_carry_i_10
       (.I0(n25__0_carry_i_3_n_0),
        .I1(B[1]),
        .I2(n4[4]),
        .I3(n25__0_carry_i_18_n_0),
        .I4(n4[5]),
        .I5(B[0]),
        .O(n25__0_carry_i_10_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__0_carry_i_11
       (.I0(n25__0_carry_i_4_n_0),
        .I1(B[1]),
        .I2(n4[3]),
        .I3(n25__0_carry_i_19_n_0),
        .I4(n4[4]),
        .I5(B[0]),
        .O(n25__0_carry_i_11_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n25__0_carry_i_12
       (.I0(n4[2]),
        .I1(n25__0_carry_i_20_n_0),
        .I2(n4[1]),
        .I3(B[1]),
        .I4(n4[0]),
        .I5(B[2]),
        .O(n25__0_carry_i_12_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n25__0_carry_i_13
       (.I0(n4[0]),
        .I1(B[2]),
        .I2(n4[1]),
        .I3(B[1]),
        .I4(B[0]),
        .I5(n4[2]),
        .O(n25__0_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__0_carry_i_14
       (.I0(B[0]),
        .I1(n4[1]),
        .I2(B[1]),
        .I3(n4[0]),
        .O(n25__0_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__0_carry_i_15
       (.I0(n4[0]),
        .I1(B[0]),
        .O(n25__0_carry_i_15_n_0));
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_16
       (.I0(n4[5]),
        .I1(B[2]),
        .O(n25__0_carry_i_16_n_0));
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_17
       (.I0(n4[4]),
        .I1(B[2]),
        .O(n25__0_carry_i_17_n_0));
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_18
       (.I0(n4[3]),
        .I1(B[2]),
        .O(n25__0_carry_i_18_n_0));
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_19
       (.I0(n4[2]),
        .I1(B[2]),
        .O(n25__0_carry_i_19_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__0_carry_i_2
       (.I0(B[2]),
        .I1(n4[3]),
        .I2(B[1]),
        .I3(n4[4]),
        .I4(B[0]),
        .I5(n4[5]),
        .O(n25__0_carry_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__0_carry_i_20
       (.I0(n4[3]),
        .I1(B[0]),
        .O(n25__0_carry_i_20_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__0_carry_i_3
       (.I0(B[2]),
        .I1(n4[2]),
        .I2(B[1]),
        .I3(n4[3]),
        .I4(B[0]),
        .I5(n4[4]),
        .O(n25__0_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__0_carry_i_4
       (.I0(B[2]),
        .I1(n4[1]),
        .I2(B[1]),
        .I3(n4[2]),
        .I4(B[0]),
        .I5(n4[3]),
        .O(n25__0_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n25__0_carry_i_5
       (.I0(B[1]),
        .I1(n4[2]),
        .I2(B[2]),
        .I3(n4[1]),
        .I4(n4[3]),
        .I5(B[0]),
        .O(n25__0_carry_i_5_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__0_carry_i_6
       (.I0(B[1]),
        .I1(n4[1]),
        .I2(B[2]),
        .I3(n4[0]),
        .O(n25__0_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__0_carry_i_7
       (.I0(B[0]),
        .I1(n4[1]),
        .O(n25__0_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n25__0_carry_i_8
       (.I0(n25__0_carry_i_1_n_0),
        .I1(B[1]),
        .I2(n4[6]),
        .I3(n25__0_carry_i_16_n_0),
        .I4(n4[7]),
        .I5(B[0]),
        .O(n25__0_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__0_carry_i_9
       (.I0(n25__0_carry_i_2_n_0),
        .I1(B[1]),
        .I2(n4[5]),
        .I3(n25__0_carry_i_17_n_0),
        .I4(n4[6]),
        .I5(B[0]),
        .O(n25__0_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__27_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__27_carry_n_0,n25__27_carry_n_1,n25__27_carry_n_2,n25__27_carry_n_3,n25__27_carry_n_4,n25__27_carry_n_5,n25__27_carry_n_6,n25__27_carry_n_7}),
        .DI({n25__27_carry_i_1_n_0,n25__27_carry_i_2_n_0,n25__27_carry_i_3_n_0,n25__27_carry_i_4_n_0,n25__27_carry_i_5_n_0,n25__27_carry_i_6_n_0,n25__27_carry_i_7_n_0,1'b0}),
        .O({n25__27_carry_n_8,n25__27_carry_n_9,n25__27_carry_n_10,n25__27_carry_n_11,n25__27_carry_n_12,n25__27_carry_n_13,n25__27_carry_n_14,n25__27_carry_n_15}),
        .S({n25__27_carry_i_8_n_0,n25__27_carry_i_9_n_0,n25__27_carry_i_10_n_0,n25__27_carry_i_11_n_0,n25__27_carry_i_12_n_0,n25__27_carry_i_13_n_0,n25__27_carry_i_14_n_0,n25__27_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__27_carry__0
       (.CI(n25__27_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__27_carry__0_CO_UNCONNECTED[7:3],n25__27_carry__0_n_5,NLW_n25__27_carry__0_CO_UNCONNECTED[1],n25__27_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25__27_carry__0_i_1_n_0,n25__27_carry__0_i_2_n_0}),
        .O({NLW_n25__27_carry__0_O_UNCONNECTED[7:2],n25__27_carry__0_n_14,n25__27_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n25__27_carry__0_i_3_n_0,n25__27_carry__0_i_4_n_0}));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__27_carry__0_i_1
       (.I0(B[4]),
        .I1(n4[7]),
        .I2(B[5]),
        .I3(n4[6]),
        .O(n25__27_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h8000F888F888F888)) 
    n25__27_carry__0_i_2
       (.I0(B[5]),
        .I1(n4[5]),
        .I2(B[4]),
        .I3(n4[6]),
        .I4(B[3]),
        .I5(n4[7]),
        .O(n25__27_carry__0_i_2_n_0));
  LUT4 #(
    .INIT(16'h2F5F)) 
    n25__27_carry__0_i_3
       (.I0(n4[6]),
        .I1(B[4]),
        .I2(B[5]),
        .I3(n4[7]),
        .O(n25__27_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h2450F30F4BFFC3FF)) 
    n25__27_carry__0_i_4
       (.I0(B[3]),
        .I1(n4[5]),
        .I2(n4[6]),
        .I3(B[5]),
        .I4(n4[7]),
        .I5(B[4]),
        .O(n25__27_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__27_carry_i_1
       (.I0(B[5]),
        .I1(n4[4]),
        .I2(B[4]),
        .I3(n4[5]),
        .I4(B[3]),
        .I5(n4[6]),
        .O(n25__27_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__27_carry_i_10
       (.I0(n25__27_carry_i_3_n_0),
        .I1(B[4]),
        .I2(n4[4]),
        .I3(n25__27_carry_i_18_n_0),
        .I4(n4[5]),
        .I5(B[3]),
        .O(n25__27_carry_i_10_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__27_carry_i_11
       (.I0(n25__27_carry_i_4_n_0),
        .I1(B[4]),
        .I2(n4[3]),
        .I3(n25__27_carry_i_19_n_0),
        .I4(n4[4]),
        .I5(B[3]),
        .O(n25__27_carry_i_11_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    n25__27_carry_i_12
       (.I0(n4[2]),
        .I1(n25__27_carry_i_20_n_0),
        .I2(n4[1]),
        .I3(B[4]),
        .I4(n4[0]),
        .I5(B[5]),
        .O(n25__27_carry_i_12_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n25__27_carry_i_13
       (.I0(n4[0]),
        .I1(B[5]),
        .I2(n4[1]),
        .I3(B[4]),
        .I4(B[3]),
        .I5(n4[2]),
        .O(n25__27_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__27_carry_i_14
       (.I0(B[3]),
        .I1(n4[1]),
        .I2(B[4]),
        .I3(n4[0]),
        .O(n25__27_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__27_carry_i_15
       (.I0(n4[0]),
        .I1(B[3]),
        .O(n25__27_carry_i_15_n_0));
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_16
       (.I0(n4[5]),
        .I1(B[5]),
        .O(n25__27_carry_i_16_n_0));
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_17
       (.I0(n4[4]),
        .I1(B[5]),
        .O(n25__27_carry_i_17_n_0));
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_18
       (.I0(n4[3]),
        .I1(B[5]),
        .O(n25__27_carry_i_18_n_0));
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_19
       (.I0(n4[2]),
        .I1(B[5]),
        .O(n25__27_carry_i_19_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__27_carry_i_2
       (.I0(B[5]),
        .I1(n4[3]),
        .I2(B[4]),
        .I3(n4[4]),
        .I4(B[3]),
        .I5(n4[5]),
        .O(n25__27_carry_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT2 #(
    .INIT(4'h7)) 
    n25__27_carry_i_20
       (.I0(n4[3]),
        .I1(B[3]),
        .O(n25__27_carry_i_20_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__27_carry_i_3
       (.I0(B[5]),
        .I1(n4[2]),
        .I2(B[4]),
        .I3(n4[3]),
        .I4(B[3]),
        .I5(n4[4]),
        .O(n25__27_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    n25__27_carry_i_4
       (.I0(B[5]),
        .I1(n4[1]),
        .I2(B[4]),
        .I3(n4[2]),
        .I4(B[3]),
        .I5(n4[3]),
        .O(n25__27_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    n25__27_carry_i_5
       (.I0(B[4]),
        .I1(n4[2]),
        .I2(B[5]),
        .I3(n4[1]),
        .I4(n4[3]),
        .I5(B[3]),
        .O(n25__27_carry_i_5_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__27_carry_i_6
       (.I0(B[4]),
        .I1(n4[1]),
        .I2(B[5]),
        .I3(n4[0]),
        .O(n25__27_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__27_carry_i_7
       (.I0(B[3]),
        .I1(n4[1]),
        .O(n25__27_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'h6A95956A956A956A)) 
    n25__27_carry_i_8
       (.I0(n25__27_carry_i_1_n_0),
        .I1(B[4]),
        .I2(n4[6]),
        .I3(n25__27_carry_i_16_n_0),
        .I4(n4[7]),
        .I5(B[3]),
        .O(n25__27_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    n25__27_carry_i_9
       (.I0(n25__27_carry_i_2_n_0),
        .I1(B[4]),
        .I2(n4[5]),
        .I3(n25__27_carry_i_17_n_0),
        .I4(n4[6]),
        .I5(B[3]),
        .O(n25__27_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__56_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__56_carry_n_0,n25__56_carry_n_1,n25__56_carry_n_2,n25__56_carry_n_3,n25__56_carry_n_4,n25__56_carry_n_5,n25__56_carry_n_6,n25__56_carry_n_7}),
        .DI({n25__56_carry_i_1_n_0,n25__56_carry_i_2_n_0,n25__56_carry_i_3_n_0,n25__56_carry_i_4_n_0,n25__56_carry_i_5_n_0,n25__56_carry_i_6_n_0,n25__56_carry_i_7_n_0,1'b0}),
        .O({n25__56_carry_n_8,n25__56_carry_n_9,n25__56_carry_n_10,n25__56_carry_n_11,n25__56_carry_n_12,n25__56_carry_n_13,n25__56_carry_n_14,n25__56_carry_n_15}),
        .S({n25__56_carry_i_8_n_0,n25__56_carry_i_9_n_0,n25__56_carry_i_10_n_0,n25__56_carry_i_11_n_0,n25__56_carry_i_12_n_0,n25__56_carry_i_13_n_0,n25__56_carry_i_14_n_0,n25__56_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__56_carry__0
       (.CI(n25__56_carry_n_0),
        .CI_TOP(1'b0),
        .CO(NLW_n25__56_carry__0_CO_UNCONNECTED[7:0]),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({NLW_n25__56_carry__0_O_UNCONNECTED[7:1],n25__56_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25__56_carry__0_i_1_n_0}));
  LUT4 #(
    .INIT(16'hE53F)) 
    n25__56_carry__0_i_1
       (.I0(B[6]),
        .I1(n4[6]),
        .I2(B[7]),
        .I3(n4[7]),
        .O(n25__56_carry__0_i_1_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__56_carry_i_1
       (.I0(B[7]),
        .I1(n4[5]),
        .I2(B[6]),
        .I3(n4[6]),
        .O(n25__56_carry_i_1_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n25__56_carry_i_10
       (.I0(n4[3]),
        .I1(n4[4]),
        .I2(B[7]),
        .I3(n4[5]),
        .I4(B[6]),
        .O(n25__56_carry_i_10_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n25__56_carry_i_11
       (.I0(n4[2]),
        .I1(n4[3]),
        .I2(B[7]),
        .I3(n4[4]),
        .I4(B[6]),
        .O(n25__56_carry_i_11_n_0));
  LUT5 #(
    .INIT(32'h9F606060)) 
    n25__56_carry_i_12
       (.I0(n4[1]),
        .I1(n4[2]),
        .I2(B[7]),
        .I3(n4[3]),
        .I4(B[6]),
        .O(n25__56_carry_i_12_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    n25__56_carry_i_13
       (.I0(B[7]),
        .I1(n4[1]),
        .I2(B[6]),
        .I3(n4[2]),
        .O(n25__56_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h8777)) 
    n25__56_carry_i_14
       (.I0(B[7]),
        .I1(n4[0]),
        .I2(B[6]),
        .I3(n4[1]),
        .O(n25__56_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__56_carry_i_15
       (.I0(n4[0]),
        .I1(B[6]),
        .O(n25__56_carry_i_15_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__56_carry_i_2
       (.I0(B[7]),
        .I1(n4[4]),
        .I2(B[6]),
        .I3(n4[5]),
        .O(n25__56_carry_i_2_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__56_carry_i_3
       (.I0(B[7]),
        .I1(n4[3]),
        .I2(B[6]),
        .I3(n4[4]),
        .O(n25__56_carry_i_3_n_0));
  LUT4 #(
    .INIT(16'h7000)) 
    n25__56_carry_i_4
       (.I0(B[7]),
        .I1(n4[2]),
        .I2(B[6]),
        .I3(n4[3]),
        .O(n25__56_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n25__56_carry_i_5
       (.I0(n4[1]),
        .I1(B[7]),
        .O(n25__56_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__56_carry_i_6
       (.I0(B[7]),
        .I1(n4[1]),
        .O(n25__56_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n25__56_carry_i_7
       (.I0(n4[0]),
        .I1(B[7]),
        .O(n25__56_carry_i_7_n_0));
  LUT5 #(
    .INIT(32'h738CC0C0)) 
    n25__56_carry_i_8
       (.I0(n4[5]),
        .I1(n4[6]),
        .I2(B[7]),
        .I3(n4[7]),
        .I4(B[6]),
        .O(n25__56_carry_i_8_n_0));
  LUT5 #(
    .INIT(32'h8C733F3F)) 
    n25__56_carry_i_9
       (.I0(n4[4]),
        .I1(n4[5]),
        .I2(B[7]),
        .I3(n4[6]),
        .I4(B[6]),
        .O(n25__56_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__81_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__81_carry_n_0,n25__81_carry_n_1,n25__81_carry_n_2,n25__81_carry_n_3,n25__81_carry_n_4,n25__81_carry_n_5,n25__81_carry_n_6,n25__81_carry_n_7}),
        .DI({n25__81_carry_i_1_n_0,n25__81_carry_i_2_n_0,n25__81_carry_i_3_n_0,n25__81_carry_i_4_n_0,n25__81_carry_i_5_n_0,n25__81_carry_i_6_n_0,n25__81_carry_i_7_n_0,1'b0}),
        .O({n26[3:0],NLW_n25__81_carry_O_UNCONNECTED[3:0]}),
        .S({n25__81_carry_i_8_n_0,n25__81_carry_i_9_n_0,n25__81_carry_i_10_n_0,n25__81_carry_i_11_n_0,n25__81_carry_i_12_n_0,n25__81_carry_i_13_n_0,n25__81_carry_i_14_n_0,n25__81_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__81_carry__0
       (.CI(n25__81_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__81_carry__0_CO_UNCONNECTED[7:3],n25__81_carry__0_n_5,n25__81_carry__0_n_6,n25__81_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n25__81_carry__0_i_1_n_0,n25__81_carry__0_i_2_n_0,n25__81_carry__0_i_3_n_0}),
        .O({NLW_n25__81_carry__0_O_UNCONNECTED[7:4],n26[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n25__81_carry__0_i_4_n_0,n25__81_carry__0_i_5_n_0,n25__81_carry__0_i_6_n_0,n25__81_carry__0_i_7_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry__0_i_1
       (.I0(n25__27_carry__0_n_14),
        .I1(n25__56_carry_n_9),
        .O(n25__81_carry__0_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry__0_i_2
       (.I0(n25__27_carry__0_n_15),
        .I1(n25__56_carry_n_10),
        .O(n25__81_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry__0_i_3
       (.I0(n25__56_carry_n_11),
        .I1(n25__27_carry_n_8),
        .I2(n25__0_carry__0_n_5),
        .O(n25__81_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n25__81_carry__0_i_4
       (.I0(n25__27_carry__0_n_5),
        .I1(n25__56_carry_n_8),
        .I2(n25__56_carry__0_n_15),
        .O(n25__81_carry__0_i_4_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__81_carry__0_i_5
       (.I0(n25__27_carry__0_n_14),
        .I1(n25__56_carry_n_9),
        .I2(n25__56_carry_n_8),
        .I3(n25__27_carry__0_n_5),
        .O(n25__81_carry__0_i_5_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__81_carry__0_i_6
       (.I0(n25__27_carry__0_n_15),
        .I1(n25__56_carry_n_10),
        .I2(n25__56_carry_n_9),
        .I3(n25__27_carry__0_n_14),
        .O(n25__81_carry__0_i_6_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n25__81_carry__0_i_7
       (.I0(n25__0_carry__0_n_5),
        .I1(n25__27_carry_n_8),
        .I2(n25__56_carry_n_11),
        .I3(n25__56_carry_n_10),
        .I4(n25__27_carry__0_n_15),
        .O(n25__81_carry__0_i_7_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry_i_1
       (.I0(n25__56_carry_n_12),
        .I1(n25__27_carry_n_9),
        .I2(n25__0_carry__0_n_14),
        .O(n25__81_carry_i_1_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_10
       (.I0(n25__56_carry_n_13),
        .I1(n25__27_carry_n_10),
        .I2(n25__0_carry__0_n_15),
        .I3(n25__81_carry_i_3_n_0),
        .O(n25__81_carry_i_10_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_11
       (.I0(n25__56_carry_n_14),
        .I1(n25__27_carry_n_11),
        .I2(n25__0_carry_n_8),
        .I3(n25__81_carry_i_4_n_0),
        .O(n25__81_carry_i_11_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_12
       (.I0(n25__56_carry_n_15),
        .I1(n25__27_carry_n_12),
        .I2(n25__0_carry_n_9),
        .I3(n25__81_carry_i_5_n_0),
        .O(n25__81_carry_i_12_n_0));
  LUT4 #(
    .INIT(16'h9666)) 
    n25__81_carry_i_13
       (.I0(n25__27_carry_n_13),
        .I1(n25__0_carry_n_10),
        .I2(n25__0_carry_n_11),
        .I3(n25__27_carry_n_14),
        .O(n25__81_carry_i_13_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__81_carry_i_14
       (.I0(n25__0_carry_n_12),
        .I1(n25__27_carry_n_15),
        .I2(n25__27_carry_n_14),
        .I3(n25__0_carry_n_11),
        .O(n25__81_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n25__81_carry_i_15
       (.I0(n25__0_carry_n_12),
        .I1(n25__27_carry_n_15),
        .O(n25__81_carry_i_15_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry_i_2
       (.I0(n25__56_carry_n_13),
        .I1(n25__27_carry_n_10),
        .I2(n25__0_carry__0_n_15),
        .O(n25__81_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry_i_3
       (.I0(n25__56_carry_n_14),
        .I1(n25__27_carry_n_11),
        .I2(n25__0_carry_n_8),
        .O(n25__81_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25__81_carry_i_4
       (.I0(n25__56_carry_n_15),
        .I1(n25__27_carry_n_12),
        .I2(n25__0_carry_n_9),
        .O(n25__81_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry_i_5
       (.I0(n25__27_carry_n_13),
        .I1(n25__0_carry_n_10),
        .O(n25__81_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry_i_6
       (.I0(n25__0_carry_n_11),
        .I1(n25__27_carry_n_14),
        .O(n25__81_carry_i_6_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__81_carry_i_7
       (.I0(n25__0_carry_n_12),
        .I1(n25__27_carry_n_15),
        .O(n25__81_carry_i_7_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_8
       (.I0(n25__81_carry_i_1_n_0),
        .I1(n25__27_carry_n_8),
        .I2(n25__56_carry_n_11),
        .I3(n25__0_carry__0_n_5),
        .O(n25__81_carry_i_8_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n25__81_carry_i_9
       (.I0(n25__56_carry_n_12),
        .I1(n25__27_carry_n_9),
        .I2(n25__0_carry__0_n_14),
        .I3(n25__81_carry_i_2_n_0),
        .O(n25__81_carry_i_9_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[0]),
        .Q(n27[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[1]),
        .Q(n27[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[2]),
        .Q(n27[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[3]),
        .Q(n27[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[4]),
        .Q(n27[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[5]),
        .Q(n27[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[6]),
        .Q(n27[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[7]),
        .Q(n27[7]),
        .R(rst_i));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_2 
       (.I0(n24[7]),
        .I1(n27[7]),
        .O(\n29[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_3 
       (.I0(n24[6]),
        .I1(n27[6]),
        .O(\n29[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_4 
       (.I0(n24[5]),
        .I1(n27[5]),
        .O(\n29[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_5 
       (.I0(n24[4]),
        .I1(n27[4]),
        .O(\n29[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_6 
       (.I0(n24[3]),
        .I1(n27[3]),
        .O(\n29[7]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_7 
       (.I0(n24[2]),
        .I1(n27[2]),
        .O(\n29[7]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_8 
       (.I0(n24[1]),
        .I1(n27[1]),
        .O(\n29[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n29[7]_i_9 
       (.I0(n24[0]),
        .I1(n27[0]),
        .O(\n29[7]_i_9_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[0]),
        .Q(n29[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[1]),
        .Q(n29[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[2]),
        .Q(n29[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[3]),
        .Q(n29[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[4]),
        .Q(n29[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[5]),
        .Q(n29[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[6]),
        .Q(n29[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n28[7]),
        .Q(n29[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n29_reg[7]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\NLW_n29_reg[7]_i_1_CO_UNCONNECTED [7],\n29_reg[7]_i_1_n_1 ,\n29_reg[7]_i_1_n_2 ,\n29_reg[7]_i_1_n_3 ,\n29_reg[7]_i_1_n_4 ,\n29_reg[7]_i_1_n_5 ,\n29_reg[7]_i_1_n_6 ,\n29_reg[7]_i_1_n_7 }),
        .DI({1'b0,n24[6:0]}),
        .O(n28),
        .S({\n29[7]_i_2_n_0 ,\n29[7]_i_3_n_0 ,\n29[7]_i_4_n_0 ,\n29[7]_i_5_n_0 ,\n29[7]_i_6_n_0 ,\n29[7]_i_7_n_0 ,\n29[7]_i_8_n_0 ,\n29[7]_i_9_n_0 }));
  LUT2 #(
    .INIT(4'h6)) 
    \n33[0]_i_1 
       (.I0(n29[0]),
        .I1(n10[0]),
        .O(n31[0]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[10]_i_1 
       (.I0(n21[2]),
        .I1(\n8_reg_n_0_[2] ),
        .I2(\n8_reg_n_0_[1] ),
        .I3(n21[1]),
        .I4(\n8_reg_n_0_[0] ),
        .I5(n21[0]),
        .O(\n33[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[11]_i_1 
       (.I0(n21[3]),
        .I1(\n8_reg_n_0_[3] ),
        .I2(\n33[12]_i_2_n_0 ),
        .O(\n33[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[12]_i_1 
       (.I0(n21[4]),
        .I1(\n8_reg_n_0_[4] ),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[3]),
        .I4(\n33[12]_i_2_n_0 ),
        .O(\n33[12]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[12]_i_2 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n33[12]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[13]_i_1 
       (.I0(n21[5]),
        .I1(\n8_reg_n_0_[5] ),
        .I2(\n33[14]_i_2_n_0 ),
        .O(\n33[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[14]_i_1 
       (.I0(n21[6]),
        .I1(\n8_reg_n_0_[6] ),
        .I2(\n8_reg_n_0_[5] ),
        .I3(n21[5]),
        .I4(\n33[14]_i_2_n_0 ),
        .O(\n33[14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[14]_i_2 
       (.I0(\n33[12]_i_2_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n33[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[15]_i_1 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n33[15]_i_2_n_0 ),
        .O(n30));
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[15]_i_2 
       (.I0(\n33[14]_i_2_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n33[15]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[1]_i_1 
       (.I0(n29[1]),
        .I1(n10[1]),
        .I2(n10[0]),
        .I3(n29[0]),
        .O(n31[1]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[2]_i_1 
       (.I0(n29[2]),
        .I1(n10[2]),
        .I2(n10[1]),
        .I3(n29[1]),
        .I4(n10[0]),
        .I5(n29[0]),
        .O(\n33[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[3]_i_1 
       (.I0(n29[3]),
        .I1(n10[3]),
        .I2(\n33[4]_i_2_n_0 ),
        .O(\n33[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[4]_i_1 
       (.I0(n29[4]),
        .I1(n10[4]),
        .I2(n10[3]),
        .I3(n29[3]),
        .I4(\n33[4]_i_2_n_0 ),
        .O(\n33[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[4]_i_2 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n33[4]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[5]_i_1 
       (.I0(n29[5]),
        .I1(n10[5]),
        .I2(\n33[6]_i_2_n_0 ),
        .O(\n33[5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[6]_i_1 
       (.I0(n29[6]),
        .I1(n10[6]),
        .I2(n10[5]),
        .I3(n29[5]),
        .I4(\n33[6]_i_2_n_0 ),
        .O(\n33[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[6]_i_2 
       (.I0(\n33[4]_i_2_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n33[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[7]_i_1 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n33[7]_i_2_n_0 ),
        .O(n31[7]));
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[7]_i_2 
       (.I0(\n33[6]_i_2_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n33[7]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[9]_i_1 
       (.I0(n21[1]),
        .I1(\n8_reg_n_0_[1] ),
        .I2(\n8_reg_n_0_[0] ),
        .I3(n21[0]),
        .O(\n33[9]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[0]),
        .Q(i1[15]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[10]_i_1_n_0 ),
        .Q(i1[24]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[11]_i_1_n_0 ),
        .Q(i1[25]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[12]_i_1_n_0 ),
        .Q(i1[26]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[13]_i_1_n_0 ),
        .Q(i1[27]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[14]_i_1_n_0 ),
        .Q(i1[28]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n30),
        .Q(i1[29]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[1]),
        .Q(i1[16]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[2]_i_1_n_0 ),
        .Q(i1[17]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[3]_i_1_n_0 ),
        .Q(i1[18]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[4]_i_1_n_0 ),
        .Q(i1[19]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[5]_i_1_n_0 ),
        .Q(i1[20]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[6]_i_1_n_0 ),
        .Q(i1[21]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[7]),
        .Q(i1[22]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[9]_i_1_n_0 ),
        .Q(i1[23]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[10]_i_1 
       (.I0(\n8_reg_n_0_[1] ),
        .I1(n21[1]),
        .I2(n21[0]),
        .I3(\n8_reg_n_0_[0] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(n341_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[11]_i_1 
       (.I0(\n37[12]_i_2_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .O(n341_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[12]_i_1 
       (.I0(\n8_reg_n_0_[3] ),
        .I1(n21[3]),
        .I2(\n37[12]_i_2_n_0 ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(n341_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[12]_i_2 
       (.I0(\n8_reg_n_0_[0] ),
        .I1(n21[0]),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n37[12]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[13]_i_1 
       (.I0(\n37[14]_i_2_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(n341_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[14]_i_1 
       (.I0(\n8_reg_n_0_[5] ),
        .I1(n21[5]),
        .I2(\n37[14]_i_2_n_0 ),
        .I3(n21[6]),
        .I4(\n8_reg_n_0_[6] ),
        .O(n341_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[14]_i_2 
       (.I0(\n37[12]_i_2_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n37[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[15]_i_1 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n37[15]_i_2_n_0 ),
        .O(n341_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[15]_i_2 
       (.I0(\n37[14]_i_2_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n37[15]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[1]_i_1 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .O(n350_out[1]));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[2]_i_1 
       (.I0(n10[1]),
        .I1(n29[1]),
        .I2(n29[0]),
        .I3(n10[0]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(n350_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[3]_i_1 
       (.I0(\n37[4]_i_2_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .O(n350_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[4]_i_1 
       (.I0(n10[3]),
        .I1(n29[3]),
        .I2(\n37[4]_i_2_n_0 ),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(n350_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[4]_i_2 
       (.I0(n10[0]),
        .I1(n29[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n37[4]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[5]_i_1 
       (.I0(\n37[6]_i_2_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(n350_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[6]_i_1 
       (.I0(n10[5]),
        .I1(n29[5]),
        .I2(\n37[6]_i_2_n_0 ),
        .I3(n29[6]),
        .I4(n10[6]),
        .O(n350_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[6]_i_2 
       (.I0(\n37[4]_i_2_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n37[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[7]_i_1 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n37[7]_i_2_n_0 ),
        .O(n350_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[7]_i_2 
       (.I0(\n37[6]_i_2_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n37[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n37[8]_i_1 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .O(n341_out[0]));
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[9]_i_1 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .O(n341_out[1]));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[2]),
        .Q(i1[9]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[3]),
        .Q(i1[10]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[4]),
        .Q(i1[11]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[5]),
        .Q(i1[12]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[6]),
        .Q(i1[13]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[7]),
        .Q(i1[14]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[1]),
        .Q(i1[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[2]),
        .Q(i1[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[3]),
        .Q(i1[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[4]),
        .Q(i1[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[5]),
        .Q(i1[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[6]),
        .Q(i1[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[7]),
        .Q(i1[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[0]),
        .Q(i1[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[1]),
        .Q(i1[8]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[0]),
        .Q(n4[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[1]),
        .Q(n4[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[2]),
        .Q(n4[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[3]),
        .Q(n4[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[4]),
        .Q(n4[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[5]),
        .Q(n4[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[6]),
        .Q(n4[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s2_3[7]),
        .Q(n4[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[0]),
        .Q(\n7_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[1]),
        .Q(\n7_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[2]),
        .Q(\n7_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[3]),
        .Q(\n7_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[4]),
        .Q(\n7_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[5]),
        .Q(\n7_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[6]),
        .Q(\n7_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[7]),
        .Q(\n7_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[0] ),
        .Q(\n8_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[1] ),
        .Q(\n8_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[2] ),
        .Q(\n8_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[3] ),
        .Q(\n8_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[4] ),
        .Q(\n8_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[5] ),
        .Q(\n8_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[6] ),
        .Q(\n8_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[7] ),
        .Q(\n8_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[0] ),
        .Q(\n9_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[1] ),
        .Q(\n9_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[2] ),
        .Q(\n9_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[3] ),
        .Q(\n9_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[4] ),
        .Q(\n9_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[5] ),
        .Q(\n9_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[6] ),
        .Q(\n9_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[7] ),
        .Q(\n9_reg_n_0_[7] ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_21" *) 
module switch_elements_cf_fft_512_8_21
   (\n9_reg[0] ,
    D,
    s1_3,
    rst_i,
    enable_i,
    clk_i,
    n22,
    \n1_reg[15] ,
    \n4_reg[7] );
  output \n9_reg[0] ;
  output [15:0]D;
  output [15:0]s1_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [7:0]n22;
  input [15:0]\n1_reg[15] ;
  input [7:0]\n4_reg[7] ;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire [15:0]\n1_reg[15] ;
  wire [7:0]n22;
  wire [15:0]n33;
  wire [15:1]n37;
  wire n4;
  wire [7:0]\n4_reg[7] ;
  wire \n9_reg[0] ;
  wire rst_i;
  wire [15:0]s1_3;

  switch_elements_cf_fft_512_8_37_22 s25
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .\n1_reg[15]_0 (\n1_reg[15] ),
        .n22_0(n22),
        .\n4_reg[7]_0 (\n4_reg[7] ),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_31_23 s26
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i8(i8),
        .n4(n4),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_27_24 s27
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .i8(i8),
        .\n9_reg[0]_0 (\n9_reg[0] ),
        .rst_i(rst_i),
        .s1_3(s1_3));
  switch_elements_cf_fft_512_8_26_25 s28
       (.D(D),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n37[8],n33[7:0],n37[15:9],n37[7:1]}),
        .i8(i8),
        .\n1_reg[15] (\n9_reg[0] ),
        .n4(n4),
        .rst_i(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_26" *) 
module switch_elements_cf_fft_512_8_26
   (D,
    n4,
    \n1_reg[0] ,
    i8,
    rst_i,
    enable_i,
    clk_i,
    i1);
  output [15:0]D;
  output n4;
  input \n1_reg[0] ;
  input [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [29:0]i1;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [6:0]n11a;
  wire [5:0]n11a__0;
  wire n11m_reg_0_63_0_6_n_0;
  wire n11m_reg_0_63_0_6_n_1;
  wire n11m_reg_0_63_0_6_n_2;
  wire n11m_reg_0_63_0_6_n_3;
  wire n11m_reg_0_63_0_6_n_4;
  wire n11m_reg_0_63_0_6_n_5;
  wire n11m_reg_0_63_0_6_n_6;
  wire n11m_reg_0_63_14_20_n_0;
  wire n11m_reg_0_63_14_20_n_1;
  wire n11m_reg_0_63_14_20_n_2;
  wire n11m_reg_0_63_14_20_n_3;
  wire n11m_reg_0_63_14_20_n_4;
  wire n11m_reg_0_63_14_20_n_5;
  wire n11m_reg_0_63_14_20_n_6;
  wire n11m_reg_0_63_21_27_n_0;
  wire n11m_reg_0_63_21_27_n_1;
  wire n11m_reg_0_63_21_27_n_2;
  wire n11m_reg_0_63_21_27_n_3;
  wire n11m_reg_0_63_21_27_n_4;
  wire n11m_reg_0_63_21_27_n_5;
  wire n11m_reg_0_63_21_27_n_6;
  wire n11m_reg_0_63_28_31_n_0;
  wire n11m_reg_0_63_28_31_n_1;
  wire n11m_reg_0_63_28_31_n_2;
  wire n11m_reg_0_63_28_31_n_3;
  wire n11m_reg_0_63_7_13_n_0;
  wire n11m_reg_0_63_7_13_n_1;
  wire n11m_reg_0_63_7_13_n_2;
  wire n11m_reg_0_63_7_13_n_3;
  wire n11m_reg_0_63_7_13_n_4;
  wire n11m_reg_0_63_7_13_n_5;
  wire n11m_reg_0_63_7_13_n_6;
  wire \n1[0]_i_2__5_n_0 ;
  wire \n1[0]_i_3__5_n_0 ;
  wire \n1[10]_i_2__5_n_0 ;
  wire \n1[10]_i_3__5_n_0 ;
  wire \n1[11]_i_2__5_n_0 ;
  wire \n1[11]_i_3__5_n_0 ;
  wire \n1[12]_i_2__5_n_0 ;
  wire \n1[12]_i_3__5_n_0 ;
  wire \n1[13]_i_2__5_n_0 ;
  wire \n1[13]_i_3__5_n_0 ;
  wire \n1[14]_i_2__5_n_0 ;
  wire \n1[14]_i_3__5_n_0 ;
  wire \n1[15]_i_2__5_n_0 ;
  wire \n1[15]_i_3__5_n_0 ;
  wire \n1[1]_i_2__5_n_0 ;
  wire \n1[1]_i_3__5_n_0 ;
  wire \n1[2]_i_2__5_n_0 ;
  wire \n1[2]_i_3__5_n_0 ;
  wire \n1[3]_i_2__5_n_0 ;
  wire \n1[3]_i_3__5_n_0 ;
  wire \n1[4]_i_2__5_n_0 ;
  wire \n1[4]_i_3__5_n_0 ;
  wire \n1[5]_i_2__5_n_0 ;
  wire \n1[5]_i_3__5_n_0 ;
  wire \n1[6]_i_2__5_n_0 ;
  wire \n1[6]_i_3__5_n_0 ;
  wire \n1[7]_i_2__5_n_0 ;
  wire \n1[7]_i_3__5_n_0 ;
  wire \n1[8]_i_2__5_n_0 ;
  wire \n1[8]_i_3__5_n_0 ;
  wire \n1[9]_i_2__5_n_0 ;
  wire \n1[9]_i_3__5_n_0 ;
  wire \n1_reg[0] ;
  wire [6:0]n2__0;
  wire \n3[6]_i_2__6_n_0 ;
  wire [6:0]n3_reg;
  wire n4;
  wire \n5[0]_i_2__6_n_0 ;
  wire n9m_reg_0_63_0_6_n_0;
  wire n9m_reg_0_63_0_6_n_1;
  wire n9m_reg_0_63_0_6_n_2;
  wire n9m_reg_0_63_0_6_n_3;
  wire n9m_reg_0_63_0_6_n_4;
  wire n9m_reg_0_63_0_6_n_5;
  wire n9m_reg_0_63_0_6_n_6;
  wire n9m_reg_0_63_14_20_n_0;
  wire n9m_reg_0_63_14_20_n_1;
  wire n9m_reg_0_63_14_20_n_2;
  wire n9m_reg_0_63_14_20_n_3;
  wire n9m_reg_0_63_14_20_n_4;
  wire n9m_reg_0_63_14_20_n_5;
  wire n9m_reg_0_63_14_20_n_6;
  wire n9m_reg_0_63_21_27_n_0;
  wire n9m_reg_0_63_21_27_n_1;
  wire n9m_reg_0_63_21_27_n_2;
  wire n9m_reg_0_63_21_27_n_3;
  wire n9m_reg_0_63_21_27_n_4;
  wire n9m_reg_0_63_21_27_n_5;
  wire n9m_reg_0_63_21_27_n_6;
  wire n9m_reg_0_63_28_31_n_0;
  wire n9m_reg_0_63_28_31_n_1;
  wire n9m_reg_0_63_28_31_n_2;
  wire n9m_reg_0_63_28_31_n_3;
  wire n9m_reg_0_63_7_13_n_0;
  wire n9m_reg_0_63_7_13_n_1;
  wire n9m_reg_0_63_7_13_n_2;
  wire n9m_reg_0_63_7_13_n_3;
  wire n9m_reg_0_63_7_13_n_4;
  wire n9m_reg_0_63_7_13_n_5;
  wire n9m_reg_0_63_7_13_n_6;
  wire n9m_reg_64_127_0_6_n_0;
  wire n9m_reg_64_127_0_6_n_1;
  wire n9m_reg_64_127_0_6_n_2;
  wire n9m_reg_64_127_0_6_n_3;
  wire n9m_reg_64_127_0_6_n_4;
  wire n9m_reg_64_127_0_6_n_5;
  wire n9m_reg_64_127_0_6_n_6;
  wire n9m_reg_64_127_14_20_n_0;
  wire n9m_reg_64_127_14_20_n_1;
  wire n9m_reg_64_127_14_20_n_2;
  wire n9m_reg_64_127_14_20_n_3;
  wire n9m_reg_64_127_14_20_n_4;
  wire n9m_reg_64_127_14_20_n_5;
  wire n9m_reg_64_127_14_20_n_6;
  wire n9m_reg_64_127_21_27_n_0;
  wire n9m_reg_64_127_21_27_n_1;
  wire n9m_reg_64_127_21_27_n_2;
  wire n9m_reg_64_127_21_27_n_3;
  wire n9m_reg_64_127_21_27_n_4;
  wire n9m_reg_64_127_21_27_n_5;
  wire n9m_reg_64_127_21_27_n_6;
  wire n9m_reg_64_127_28_31_n_0;
  wire n9m_reg_64_127_28_31_n_1;
  wire n9m_reg_64_127_28_31_n_2;
  wire n9m_reg_64_127_28_31_n_3;
  wire n9m_reg_64_127_7_13_n_0;
  wire n9m_reg_64_127_7_13_n_1;
  wire n9m_reg_64_127_7_13_n_2;
  wire n9m_reg_64_127_7_13_n_3;
  wire n9m_reg_64_127_7_13_n_4;
  wire n9m_reg_64_127_7_13_n_5;
  wire n9m_reg_64_127_7_13_n_6;
  wire rst_i;
  wire NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED;

  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39883 n11m_reg_0_63_0_6
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_0_6_n_0),
        .DOB(n11m_reg_0_63_0_6_n_1),
        .DOC(n11m_reg_0_63_0_6_n_2),
        .DOD(n11m_reg_0_63_0_6_n_3),
        .DOE(n11m_reg_0_63_0_6_n_4),
        .DOF(n11m_reg_0_63_0_6_n_5),
        .DOG(n11m_reg_0_63_0_6_n_6),
        .DOH(NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39884 n11m_reg_0_63_14_20
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_14_20_n_0),
        .DOB(n11m_reg_0_63_14_20_n_1),
        .DOC(n11m_reg_0_63_14_20_n_2),
        .DOD(n11m_reg_0_63_14_20_n_3),
        .DOE(n11m_reg_0_63_14_20_n_4),
        .DOF(n11m_reg_0_63_14_20_n_5),
        .DOG(n11m_reg_0_63_14_20_n_6),
        .DOH(NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39885 n11m_reg_0_63_21_27
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_21_27_n_0),
        .DOB(n11m_reg_0_63_21_27_n_1),
        .DOC(n11m_reg_0_63_21_27_n_2),
        .DOD(n11m_reg_0_63_21_27_n_3),
        .DOE(n11m_reg_0_63_21_27_n_4),
        .DOF(n11m_reg_0_63_21_27_n_5),
        .DOG(n11m_reg_0_63_21_27_n_6),
        .DOH(NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39886 n11m_reg_0_63_28_31
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_28_31_n_0),
        .DOB(n11m_reg_0_63_28_31_n_1),
        .DOC(n11m_reg_0_63_28_31_n_2),
        .DOD(n11m_reg_0_63_28_31_n_3),
        .DOE(NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39887 n11m_reg_0_63_7_13
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_7_13_n_0),
        .DOB(n11m_reg_0_63_7_13_n_1),
        .DOC(n11m_reg_0_63_7_13_n_2),
        .DOD(n11m_reg_0_63_7_13_n_3),
        .DOE(n11m_reg_0_63_7_13_n_4),
        .DOF(n11m_reg_0_63_7_13_n_5),
        .DOG(n11m_reg_0_63_7_13_n_6),
        .DOH(NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[0]_i_1__5 
       (.I0(n11m_reg_0_63_0_6_n_0),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[0]_i_2__5_n_0 ),
        .I4(\n1[0]_i_3__5_n_0 ),
        .O(D[0]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[0]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_0),
        .O(\n1[0]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[0]_i_3__5 
       (.I0(n11m_reg_0_63_14_20_n_2),
        .I1(n9m_reg_64_127_14_20_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[0]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[10]_i_1__5 
       (.I0(n11m_reg_0_63_7_13_n_3),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[10]_i_2__5_n_0 ),
        .I4(\n1[10]_i_3__5_n_0 ),
        .O(D[10]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[10]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_3),
        .O(\n1[10]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[10]_i_3__5 
       (.I0(n11m_reg_0_63_21_27_n_5),
        .I1(n9m_reg_64_127_21_27_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[10]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[11]_i_1__5 
       (.I0(n11m_reg_0_63_7_13_n_4),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[11]_i_2__5_n_0 ),
        .I4(\n1[11]_i_3__5_n_0 ),
        .O(D[11]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[11]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_4),
        .O(\n1[11]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[11]_i_3__5 
       (.I0(n11m_reg_0_63_21_27_n_6),
        .I1(n9m_reg_64_127_21_27_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[11]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[12]_i_1__5 
       (.I0(n11m_reg_0_63_7_13_n_5),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[12]_i_2__5_n_0 ),
        .I4(\n1[12]_i_3__5_n_0 ),
        .O(D[12]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[12]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_5),
        .O(\n1[12]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[12]_i_3__5 
       (.I0(n11m_reg_0_63_28_31_n_0),
        .I1(n9m_reg_64_127_28_31_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[12]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[13]_i_1__5 
       (.I0(n11m_reg_0_63_7_13_n_6),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[13]_i_2__5_n_0 ),
        .I4(\n1[13]_i_3__5_n_0 ),
        .O(D[13]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[13]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_6),
        .O(\n1[13]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[13]_i_3__5 
       (.I0(n11m_reg_0_63_28_31_n_1),
        .I1(n9m_reg_64_127_28_31_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[13]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[14]_i_1__5 
       (.I0(n11m_reg_0_63_14_20_n_0),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[14]_i_2__5_n_0 ),
        .I4(\n1[14]_i_3__5_n_0 ),
        .O(D[14]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[14]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_0),
        .O(\n1[14]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[14]_i_3__5 
       (.I0(n11m_reg_0_63_28_31_n_2),
        .I1(n9m_reg_64_127_28_31_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[14]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[15]_i_1__5 
       (.I0(n11m_reg_0_63_14_20_n_1),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[15]_i_2__5_n_0 ),
        .I4(\n1[15]_i_3__5_n_0 ),
        .O(D[15]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[15]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_1),
        .O(\n1[15]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[15]_i_3__5 
       (.I0(n11m_reg_0_63_28_31_n_3),
        .I1(n9m_reg_64_127_28_31_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[15]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[1]_i_1__5 
       (.I0(n11m_reg_0_63_0_6_n_1),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[1]_i_2__5_n_0 ),
        .I4(\n1[1]_i_3__5_n_0 ),
        .O(D[1]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[1]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_1),
        .O(\n1[1]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[1]_i_3__5 
       (.I0(n11m_reg_0_63_14_20_n_3),
        .I1(n9m_reg_64_127_14_20_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[1]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[2]_i_1__5 
       (.I0(n11m_reg_0_63_0_6_n_2),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[2]_i_2__5_n_0 ),
        .I4(\n1[2]_i_3__5_n_0 ),
        .O(D[2]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[2]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_2),
        .O(\n1[2]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[2]_i_3__5 
       (.I0(n11m_reg_0_63_14_20_n_4),
        .I1(n9m_reg_64_127_14_20_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[2]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[3]_i_1__5 
       (.I0(n11m_reg_0_63_0_6_n_3),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[3]_i_2__5_n_0 ),
        .I4(\n1[3]_i_3__5_n_0 ),
        .O(D[3]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[3]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_3),
        .O(\n1[3]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[3]_i_3__5 
       (.I0(n11m_reg_0_63_14_20_n_5),
        .I1(n9m_reg_64_127_14_20_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[3]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[4]_i_1__5 
       (.I0(n11m_reg_0_63_0_6_n_4),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[4]_i_2__5_n_0 ),
        .I4(\n1[4]_i_3__5_n_0 ),
        .O(D[4]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[4]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_4),
        .O(\n1[4]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[4]_i_3__5 
       (.I0(n11m_reg_0_63_14_20_n_6),
        .I1(n9m_reg_64_127_14_20_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[4]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[5]_i_1__5 
       (.I0(n11m_reg_0_63_0_6_n_5),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[5]_i_2__5_n_0 ),
        .I4(\n1[5]_i_3__5_n_0 ),
        .O(D[5]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[5]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_5),
        .O(\n1[5]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[5]_i_3__5 
       (.I0(n11m_reg_0_63_21_27_n_0),
        .I1(n9m_reg_64_127_21_27_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[5]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[6]_i_1__5 
       (.I0(n11m_reg_0_63_0_6_n_6),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[6]_i_2__5_n_0 ),
        .I4(\n1[6]_i_3__5_n_0 ),
        .O(D[6]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[6]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_6),
        .O(\n1[6]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[6]_i_3__5 
       (.I0(n11m_reg_0_63_21_27_n_1),
        .I1(n9m_reg_64_127_21_27_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[6]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[7]_i_1__5 
       (.I0(n11m_reg_0_63_7_13_n_0),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[7]_i_2__5_n_0 ),
        .I4(\n1[7]_i_3__5_n_0 ),
        .O(D[7]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[7]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_0),
        .O(\n1[7]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[7]_i_3__5 
       (.I0(n11m_reg_0_63_21_27_n_2),
        .I1(n9m_reg_64_127_21_27_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[7]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[8]_i_1__5 
       (.I0(n11m_reg_0_63_7_13_n_1),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[8]_i_2__5_n_0 ),
        .I4(\n1[8]_i_3__5_n_0 ),
        .O(D[8]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[8]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_1),
        .O(\n1[8]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[8]_i_3__5 
       (.I0(n11m_reg_0_63_21_27_n_3),
        .I1(n9m_reg_64_127_21_27_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[8]_i_3__5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[9]_i_1__5 
       (.I0(n11m_reg_0_63_7_13_n_2),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[9]_i_2__5_n_0 ),
        .I4(\n1[9]_i_3__5_n_0 ),
        .O(D[9]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[9]_i_2__5 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_2),
        .O(\n1[9]_i_2__5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[9]_i_3__5 
       (.I0(n11m_reg_0_63_21_27_n_4),
        .I1(n9m_reg_64_127_21_27_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[9]_i_3__5_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__13 
       (.I0(n3_reg[0]),
        .O(n2__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__13 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__13 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__13 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__13 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__0[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__13 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__0[5]));
  LUT3 #(
    .INIT(8'hD2)) 
    \n3[6]_i_1__6 
       (.I0(n3_reg[5]),
        .I1(\n3[6]_i_2__6_n_0 ),
        .I2(n3_reg[6]),
        .O(n2__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \n3[6]_i_2__6 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(\n3[6]_i_2__6_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[6]),
        .Q(n3_reg[6]),
        .R(rst_i));
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \n5[0]_i_1__6 
       (.I0(n3_reg[0]),
        .I1(\n5[0]_i_2__6_n_0 ),
        .I2(i8),
        .O(n4));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \n5[0]_i_2__6 
       (.I0(n3_reg[3]),
        .I1(n3_reg[4]),
        .I2(n3_reg[1]),
        .I3(n3_reg[2]),
        .I4(n3_reg[6]),
        .I5(n3_reg[5]),
        .O(\n5[0]_i_2__6_n_0 ));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[6]),
        .Q(n11a[6]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39888 n9m_reg_0_63_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_0_6_n_0),
        .DOB(n9m_reg_0_63_0_6_n_1),
        .DOC(n9m_reg_0_63_0_6_n_2),
        .DOD(n9m_reg_0_63_0_6_n_3),
        .DOE(n9m_reg_0_63_0_6_n_4),
        .DOF(n9m_reg_0_63_0_6_n_5),
        .DOG(n9m_reg_0_63_0_6_n_6),
        .DOH(NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39889 n9m_reg_0_63_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_14_20_n_0),
        .DOB(n9m_reg_0_63_14_20_n_1),
        .DOC(n9m_reg_0_63_14_20_n_2),
        .DOD(n9m_reg_0_63_14_20_n_3),
        .DOE(n9m_reg_0_63_14_20_n_4),
        .DOF(n9m_reg_0_63_14_20_n_5),
        .DOG(n9m_reg_0_63_14_20_n_6),
        .DOH(NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39890 n9m_reg_0_63_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_21_27_n_0),
        .DOB(n9m_reg_0_63_21_27_n_1),
        .DOC(n9m_reg_0_63_21_27_n_2),
        .DOD(n9m_reg_0_63_21_27_n_3),
        .DOE(n9m_reg_0_63_21_27_n_4),
        .DOF(n9m_reg_0_63_21_27_n_5),
        .DOG(n9m_reg_0_63_21_27_n_6),
        .DOH(NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39891 n9m_reg_0_63_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_28_31_n_0),
        .DOB(n9m_reg_0_63_28_31_n_1),
        .DOC(n9m_reg_0_63_28_31_n_2),
        .DOD(n9m_reg_0_63_28_31_n_3),
        .DOE(NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39892 n9m_reg_0_63_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_7_13_n_0),
        .DOB(n9m_reg_0_63_7_13_n_1),
        .DOC(n9m_reg_0_63_7_13_n_2),
        .DOD(n9m_reg_0_63_7_13_n_3),
        .DOE(n9m_reg_0_63_7_13_n_4),
        .DOF(n9m_reg_0_63_7_13_n_5),
        .DOG(n9m_reg_0_63_7_13_n_6),
        .DOH(NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39893 n9m_reg_64_127_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_0_6_n_0),
        .DOB(n9m_reg_64_127_0_6_n_1),
        .DOC(n9m_reg_64_127_0_6_n_2),
        .DOD(n9m_reg_64_127_0_6_n_3),
        .DOE(n9m_reg_64_127_0_6_n_4),
        .DOF(n9m_reg_64_127_0_6_n_5),
        .DOG(n9m_reg_64_127_0_6_n_6),
        .DOH(NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39894 n9m_reg_64_127_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_14_20_n_0),
        .DOB(n9m_reg_64_127_14_20_n_1),
        .DOC(n9m_reg_64_127_14_20_n_2),
        .DOD(n9m_reg_64_127_14_20_n_3),
        .DOE(n9m_reg_64_127_14_20_n_4),
        .DOF(n9m_reg_64_127_14_20_n_5),
        .DOG(n9m_reg_64_127_14_20_n_6),
        .DOH(NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39895 n9m_reg_64_127_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_21_27_n_0),
        .DOB(n9m_reg_64_127_21_27_n_1),
        .DOC(n9m_reg_64_127_21_27_n_2),
        .DOD(n9m_reg_64_127_21_27_n_3),
        .DOE(n9m_reg_64_127_21_27_n_4),
        .DOF(n9m_reg_64_127_21_27_n_5),
        .DOG(n9m_reg_64_127_21_27_n_6),
        .DOH(NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39896 n9m_reg_64_127_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_28_31_n_0),
        .DOB(n9m_reg_64_127_28_31_n_1),
        .DOC(n9m_reg_64_127_28_31_n_2),
        .DOD(n9m_reg_64_127_28_31_n_3),
        .DOE(NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39897 n9m_reg_64_127_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_7_13_n_0),
        .DOB(n9m_reg_64_127_7_13_n_1),
        .DOC(n9m_reg_64_127_7_13_n_2),
        .DOD(n9m_reg_64_127_7_13_n_3),
        .DOE(n9m_reg_64_127_7_13_n_4),
        .DOF(n9m_reg_64_127_7_13_n_5),
        .DOG(n9m_reg_64_127_7_13_n_6),
        .DOH(NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_26" *) 
module switch_elements_cf_fft_512_8_26_11
   (\n9_reg[0] ,
    n4,
    \n1_reg[0] ,
    i8,
    rst_i,
    enable_i,
    clk_i,
    i1);
  output [15:0]\n9_reg[0] ;
  output n4;
  input \n1_reg[0] ;
  input [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [31:0]n11;
  wire [6:0]n11a;
  wire [5:0]n11a__0;
  wire \n1[0]_i_2__1_n_0 ;
  wire \n1[0]_i_3__1_n_0 ;
  wire \n1[10]_i_2__1_n_0 ;
  wire \n1[10]_i_3__1_n_0 ;
  wire \n1[11]_i_2__1_n_0 ;
  wire \n1[11]_i_3__1_n_0 ;
  wire \n1[12]_i_2__1_n_0 ;
  wire \n1[12]_i_3__1_n_0 ;
  wire \n1[13]_i_2__1_n_0 ;
  wire \n1[13]_i_3__1_n_0 ;
  wire \n1[14]_i_2__1_n_0 ;
  wire \n1[14]_i_3__1_n_0 ;
  wire \n1[15]_i_2__1_n_0 ;
  wire \n1[15]_i_3__1_n_0 ;
  wire \n1[1]_i_2__1_n_0 ;
  wire \n1[1]_i_3__1_n_0 ;
  wire \n1[2]_i_2__1_n_0 ;
  wire \n1[2]_i_3__1_n_0 ;
  wire \n1[3]_i_2__1_n_0 ;
  wire \n1[3]_i_3__1_n_0 ;
  wire \n1[4]_i_2__1_n_0 ;
  wire \n1[4]_i_3__1_n_0 ;
  wire \n1[5]_i_2__1_n_0 ;
  wire \n1[5]_i_3__1_n_0 ;
  wire \n1[6]_i_2__1_n_0 ;
  wire \n1[6]_i_3__1_n_0 ;
  wire \n1[7]_i_2__1_n_0 ;
  wire \n1[7]_i_3__1_n_0 ;
  wire \n1[8]_i_2__1_n_0 ;
  wire \n1[8]_i_3__1_n_0 ;
  wire \n1[9]_i_2__1_n_0 ;
  wire \n1[9]_i_3__1_n_0 ;
  wire \n1_reg[0] ;
  wire [6:0]n2__0;
  wire \n3[6]_i_2__2_n_0 ;
  wire [6:0]n3_reg;
  wire n4;
  wire \n5[0]_i_2__2_n_0 ;
  wire [15:0]\n9_reg[0] ;
  wire n9m_reg_0_63_0_6_n_0;
  wire n9m_reg_0_63_0_6_n_1;
  wire n9m_reg_0_63_0_6_n_2;
  wire n9m_reg_0_63_0_6_n_3;
  wire n9m_reg_0_63_0_6_n_4;
  wire n9m_reg_0_63_0_6_n_5;
  wire n9m_reg_0_63_0_6_n_6;
  wire n9m_reg_0_63_14_20_n_0;
  wire n9m_reg_0_63_14_20_n_1;
  wire n9m_reg_0_63_14_20_n_2;
  wire n9m_reg_0_63_14_20_n_3;
  wire n9m_reg_0_63_14_20_n_4;
  wire n9m_reg_0_63_14_20_n_5;
  wire n9m_reg_0_63_14_20_n_6;
  wire n9m_reg_0_63_21_27_n_0;
  wire n9m_reg_0_63_21_27_n_1;
  wire n9m_reg_0_63_21_27_n_2;
  wire n9m_reg_0_63_21_27_n_3;
  wire n9m_reg_0_63_21_27_n_4;
  wire n9m_reg_0_63_21_27_n_5;
  wire n9m_reg_0_63_21_27_n_6;
  wire n9m_reg_0_63_28_31_n_0;
  wire n9m_reg_0_63_28_31_n_1;
  wire n9m_reg_0_63_28_31_n_2;
  wire n9m_reg_0_63_28_31_n_3;
  wire n9m_reg_0_63_7_13_n_0;
  wire n9m_reg_0_63_7_13_n_1;
  wire n9m_reg_0_63_7_13_n_2;
  wire n9m_reg_0_63_7_13_n_3;
  wire n9m_reg_0_63_7_13_n_4;
  wire n9m_reg_0_63_7_13_n_5;
  wire n9m_reg_0_63_7_13_n_6;
  wire n9m_reg_64_127_0_6_n_0;
  wire n9m_reg_64_127_0_6_n_1;
  wire n9m_reg_64_127_0_6_n_2;
  wire n9m_reg_64_127_0_6_n_3;
  wire n9m_reg_64_127_0_6_n_4;
  wire n9m_reg_64_127_0_6_n_5;
  wire n9m_reg_64_127_0_6_n_6;
  wire n9m_reg_64_127_14_20_n_0;
  wire n9m_reg_64_127_14_20_n_1;
  wire n9m_reg_64_127_14_20_n_2;
  wire n9m_reg_64_127_14_20_n_3;
  wire n9m_reg_64_127_14_20_n_4;
  wire n9m_reg_64_127_14_20_n_5;
  wire n9m_reg_64_127_14_20_n_6;
  wire n9m_reg_64_127_21_27_n_0;
  wire n9m_reg_64_127_21_27_n_1;
  wire n9m_reg_64_127_21_27_n_2;
  wire n9m_reg_64_127_21_27_n_3;
  wire n9m_reg_64_127_21_27_n_4;
  wire n9m_reg_64_127_21_27_n_5;
  wire n9m_reg_64_127_21_27_n_6;
  wire n9m_reg_64_127_28_31_n_0;
  wire n9m_reg_64_127_28_31_n_1;
  wire n9m_reg_64_127_28_31_n_2;
  wire n9m_reg_64_127_28_31_n_3;
  wire n9m_reg_64_127_7_13_n_0;
  wire n9m_reg_64_127_7_13_n_1;
  wire n9m_reg_64_127_7_13_n_2;
  wire n9m_reg_64_127_7_13_n_3;
  wire n9m_reg_64_127_7_13_n_4;
  wire n9m_reg_64_127_7_13_n_5;
  wire n9m_reg_64_127_7_13_n_6;
  wire rst_i;
  wire NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED;

  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39783 n11m_reg_0_63_0_6
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[0]),
        .DIB(i1[1]),
        .DIC(i1[2]),
        .DID(i1[3]),
        .DIE(i1[4]),
        .DIF(i1[5]),
        .DIG(i1[6]),
        .DIH(1'b0),
        .DOA(n11[0]),
        .DOB(n11[1]),
        .DOC(n11[2]),
        .DOD(n11[3]),
        .DOE(n11[4]),
        .DOF(n11[5]),
        .DOG(n11[6]),
        .DOH(NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39784 n11m_reg_0_63_14_20
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[0]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n11[14]),
        .DOB(n11[15]),
        .DOC(n11[16]),
        .DOD(n11[17]),
        .DOE(n11[18]),
        .DOF(n11[19]),
        .DOG(n11[20]),
        .DOH(NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39785 n11m_reg_0_63_21_27
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n11[21]),
        .DOB(n11[22]),
        .DOC(n11[23]),
        .DOD(n11[24]),
        .DOE(n11[25]),
        .DOF(n11[26]),
        .DOG(n11[27]),
        .DOH(NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39786 n11m_reg_0_63_28_31
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n11[28]),
        .DOB(n11[29]),
        .DOC(n11[30]),
        .DOD(n11[31]),
        .DOE(NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39787 n11m_reg_0_63_7_13
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[7]),
        .DIB(i1[22]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n11[7]),
        .DOB(n11[8]),
        .DOC(n11[9]),
        .DOD(n11[10]),
        .DOE(n11[11]),
        .DOF(n11[12]),
        .DOG(n11[13]),
        .DOH(NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[0]_i_1__1 
       (.I0(n11[0]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[0]_i_2__1_n_0 ),
        .I4(\n1[0]_i_3__1_n_0 ),
        .O(\n9_reg[0] [0]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[0]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_0),
        .O(\n1[0]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[0]_i_3__1 
       (.I0(n11[16]),
        .I1(n9m_reg_64_127_14_20_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[0]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[10]_i_1__1 
       (.I0(n11[10]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[10]_i_2__1_n_0 ),
        .I4(\n1[10]_i_3__1_n_0 ),
        .O(\n9_reg[0] [10]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[10]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_3),
        .O(\n1[10]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[10]_i_3__1 
       (.I0(n11[26]),
        .I1(n9m_reg_64_127_21_27_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[10]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[11]_i_1__1 
       (.I0(n11[11]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[11]_i_2__1_n_0 ),
        .I4(\n1[11]_i_3__1_n_0 ),
        .O(\n9_reg[0] [11]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[11]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_4),
        .O(\n1[11]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[11]_i_3__1 
       (.I0(n11[27]),
        .I1(n9m_reg_64_127_21_27_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[11]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[12]_i_1__1 
       (.I0(n11[12]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[12]_i_2__1_n_0 ),
        .I4(\n1[12]_i_3__1_n_0 ),
        .O(\n9_reg[0] [12]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[12]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_5),
        .O(\n1[12]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[12]_i_3__1 
       (.I0(n11[28]),
        .I1(n9m_reg_64_127_28_31_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[12]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[13]_i_1__1 
       (.I0(n11[13]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[13]_i_2__1_n_0 ),
        .I4(\n1[13]_i_3__1_n_0 ),
        .O(\n9_reg[0] [13]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[13]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_6),
        .O(\n1[13]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[13]_i_3__1 
       (.I0(n11[29]),
        .I1(n9m_reg_64_127_28_31_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[13]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[14]_i_1__1 
       (.I0(n11[14]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[14]_i_2__1_n_0 ),
        .I4(\n1[14]_i_3__1_n_0 ),
        .O(\n9_reg[0] [14]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[14]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_0),
        .O(\n1[14]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[14]_i_3__1 
       (.I0(n11[30]),
        .I1(n9m_reg_64_127_28_31_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[14]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[15]_i_1__1 
       (.I0(n11[15]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[15]_i_2__1_n_0 ),
        .I4(\n1[15]_i_3__1_n_0 ),
        .O(\n9_reg[0] [15]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[15]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_1),
        .O(\n1[15]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[15]_i_3__1 
       (.I0(n11[31]),
        .I1(n9m_reg_64_127_28_31_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[15]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[1]_i_1__1 
       (.I0(n11[1]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[1]_i_2__1_n_0 ),
        .I4(\n1[1]_i_3__1_n_0 ),
        .O(\n9_reg[0] [1]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[1]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_1),
        .O(\n1[1]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[1]_i_3__1 
       (.I0(n11[17]),
        .I1(n9m_reg_64_127_14_20_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[1]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[2]_i_1__1 
       (.I0(n11[2]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[2]_i_2__1_n_0 ),
        .I4(\n1[2]_i_3__1_n_0 ),
        .O(\n9_reg[0] [2]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[2]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_2),
        .O(\n1[2]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[2]_i_3__1 
       (.I0(n11[18]),
        .I1(n9m_reg_64_127_14_20_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[2]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[3]_i_1__1 
       (.I0(n11[3]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[3]_i_2__1_n_0 ),
        .I4(\n1[3]_i_3__1_n_0 ),
        .O(\n9_reg[0] [3]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[3]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_3),
        .O(\n1[3]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[3]_i_3__1 
       (.I0(n11[19]),
        .I1(n9m_reg_64_127_14_20_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[3]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[4]_i_1__1 
       (.I0(n11[4]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[4]_i_2__1_n_0 ),
        .I4(\n1[4]_i_3__1_n_0 ),
        .O(\n9_reg[0] [4]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[4]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_4),
        .O(\n1[4]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[4]_i_3__1 
       (.I0(n11[20]),
        .I1(n9m_reg_64_127_14_20_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[4]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[5]_i_1__1 
       (.I0(n11[5]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[5]_i_2__1_n_0 ),
        .I4(\n1[5]_i_3__1_n_0 ),
        .O(\n9_reg[0] [5]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[5]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_5),
        .O(\n1[5]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[5]_i_3__1 
       (.I0(n11[21]),
        .I1(n9m_reg_64_127_21_27_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[5]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[6]_i_1__1 
       (.I0(n11[6]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[6]_i_2__1_n_0 ),
        .I4(\n1[6]_i_3__1_n_0 ),
        .O(\n9_reg[0] [6]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[6]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_6),
        .O(\n1[6]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[6]_i_3__1 
       (.I0(n11[22]),
        .I1(n9m_reg_64_127_21_27_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[6]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[7]_i_1__1 
       (.I0(n11[7]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[7]_i_2__1_n_0 ),
        .I4(\n1[7]_i_3__1_n_0 ),
        .O(\n9_reg[0] [7]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[7]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_0),
        .O(\n1[7]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[7]_i_3__1 
       (.I0(n11[23]),
        .I1(n9m_reg_64_127_21_27_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[7]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[8]_i_1__1 
       (.I0(n11[8]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[8]_i_2__1_n_0 ),
        .I4(\n1[8]_i_3__1_n_0 ),
        .O(\n9_reg[0] [8]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[8]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_1),
        .O(\n1[8]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[8]_i_3__1 
       (.I0(n11[24]),
        .I1(n9m_reg_64_127_21_27_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[8]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[9]_i_1__1 
       (.I0(n11[9]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[9]_i_2__1_n_0 ),
        .I4(\n1[9]_i_3__1_n_0 ),
        .O(\n9_reg[0] [9]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[9]_i_2__1 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_2),
        .O(\n1[9]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[9]_i_3__1 
       (.I0(n11[25]),
        .I1(n9m_reg_64_127_21_27_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[9]_i_3__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__5 
       (.I0(n3_reg[0]),
        .O(n2__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__5 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__5 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__5 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__5 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__0[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__5 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__0[5]));
  LUT3 #(
    .INIT(8'hD2)) 
    \n3[6]_i_1__2 
       (.I0(n3_reg[5]),
        .I1(\n3[6]_i_2__2_n_0 ),
        .I2(n3_reg[6]),
        .O(n2__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \n3[6]_i_2__2 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(\n3[6]_i_2__2_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[6]),
        .Q(n3_reg[6]),
        .R(rst_i));
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \n5[0]_i_1__2 
       (.I0(n3_reg[0]),
        .I1(\n5[0]_i_2__2_n_0 ),
        .I2(i8),
        .O(n4));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \n5[0]_i_2__2 
       (.I0(n3_reg[3]),
        .I1(n3_reg[4]),
        .I2(n3_reg[1]),
        .I3(n3_reg[2]),
        .I4(n3_reg[6]),
        .I5(n3_reg[5]),
        .O(\n5[0]_i_2__2_n_0 ));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[6]),
        .Q(n11a[6]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39788 n9m_reg_0_63_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[0]),
        .DIB(i1[1]),
        .DIC(i1[2]),
        .DID(i1[3]),
        .DIE(i1[4]),
        .DIF(i1[5]),
        .DIG(i1[6]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_0_6_n_0),
        .DOB(n9m_reg_0_63_0_6_n_1),
        .DOC(n9m_reg_0_63_0_6_n_2),
        .DOD(n9m_reg_0_63_0_6_n_3),
        .DOE(n9m_reg_0_63_0_6_n_4),
        .DOF(n9m_reg_0_63_0_6_n_5),
        .DOG(n9m_reg_0_63_0_6_n_6),
        .DOH(NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39789 n9m_reg_0_63_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[0]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_14_20_n_0),
        .DOB(n9m_reg_0_63_14_20_n_1),
        .DOC(n9m_reg_0_63_14_20_n_2),
        .DOD(n9m_reg_0_63_14_20_n_3),
        .DOE(n9m_reg_0_63_14_20_n_4),
        .DOF(n9m_reg_0_63_14_20_n_5),
        .DOG(n9m_reg_0_63_14_20_n_6),
        .DOH(NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39790 n9m_reg_0_63_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_21_27_n_0),
        .DOB(n9m_reg_0_63_21_27_n_1),
        .DOC(n9m_reg_0_63_21_27_n_2),
        .DOD(n9m_reg_0_63_21_27_n_3),
        .DOE(n9m_reg_0_63_21_27_n_4),
        .DOF(n9m_reg_0_63_21_27_n_5),
        .DOG(n9m_reg_0_63_21_27_n_6),
        .DOH(NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39791 n9m_reg_0_63_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_28_31_n_0),
        .DOB(n9m_reg_0_63_28_31_n_1),
        .DOC(n9m_reg_0_63_28_31_n_2),
        .DOD(n9m_reg_0_63_28_31_n_3),
        .DOE(NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39792 n9m_reg_0_63_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[7]),
        .DIB(i1[22]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_7_13_n_0),
        .DOB(n9m_reg_0_63_7_13_n_1),
        .DOC(n9m_reg_0_63_7_13_n_2),
        .DOD(n9m_reg_0_63_7_13_n_3),
        .DOE(n9m_reg_0_63_7_13_n_4),
        .DOF(n9m_reg_0_63_7_13_n_5),
        .DOG(n9m_reg_0_63_7_13_n_6),
        .DOH(NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39793 n9m_reg_64_127_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[0]),
        .DIB(i1[1]),
        .DIC(i1[2]),
        .DID(i1[3]),
        .DIE(i1[4]),
        .DIF(i1[5]),
        .DIG(i1[6]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_0_6_n_0),
        .DOB(n9m_reg_64_127_0_6_n_1),
        .DOC(n9m_reg_64_127_0_6_n_2),
        .DOD(n9m_reg_64_127_0_6_n_3),
        .DOE(n9m_reg_64_127_0_6_n_4),
        .DOF(n9m_reg_64_127_0_6_n_5),
        .DOG(n9m_reg_64_127_0_6_n_6),
        .DOH(NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39794 n9m_reg_64_127_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[0]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_14_20_n_0),
        .DOB(n9m_reg_64_127_14_20_n_1),
        .DOC(n9m_reg_64_127_14_20_n_2),
        .DOD(n9m_reg_64_127_14_20_n_3),
        .DOE(n9m_reg_64_127_14_20_n_4),
        .DOF(n9m_reg_64_127_14_20_n_5),
        .DOG(n9m_reg_64_127_14_20_n_6),
        .DOH(NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39795 n9m_reg_64_127_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_21_27_n_0),
        .DOB(n9m_reg_64_127_21_27_n_1),
        .DOC(n9m_reg_64_127_21_27_n_2),
        .DOD(n9m_reg_64_127_21_27_n_3),
        .DOE(n9m_reg_64_127_21_27_n_4),
        .DOF(n9m_reg_64_127_21_27_n_5),
        .DOG(n9m_reg_64_127_21_27_n_6),
        .DOH(NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39796 n9m_reg_64_127_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_28_31_n_0),
        .DOB(n9m_reg_64_127_28_31_n_1),
        .DOC(n9m_reg_64_127_28_31_n_2),
        .DOD(n9m_reg_64_127_28_31_n_3),
        .DOE(NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39797 n9m_reg_64_127_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[7]),
        .DIB(i1[22]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_7_13_n_0),
        .DOB(n9m_reg_64_127_7_13_n_1),
        .DOC(n9m_reg_64_127_7_13_n_2),
        .DOD(n9m_reg_64_127_7_13_n_3),
        .DOE(n9m_reg_64_127_7_13_n_4),
        .DOF(n9m_reg_64_127_7_13_n_5),
        .DOG(n9m_reg_64_127_7_13_n_6),
        .DOH(NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_26" *) 
module switch_elements_cf_fft_512_8_26_14
   (\n9_reg[0] ,
    n4,
    \n1_reg[0] ,
    i8,
    rst_i,
    enable_i,
    clk_i,
    i1);
  output [15:0]\n9_reg[0] ;
  output n4;
  input \n1_reg[0] ;
  input [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [31:0]n11;
  wire [6:0]n11a;
  wire [5:0]n11a__0;
  wire \n1[0]_i_2__0_n_0 ;
  wire \n1[0]_i_3__0_n_0 ;
  wire \n1[10]_i_2__0_n_0 ;
  wire \n1[10]_i_3__0_n_0 ;
  wire \n1[11]_i_2__0_n_0 ;
  wire \n1[11]_i_3__0_n_0 ;
  wire \n1[12]_i_2__0_n_0 ;
  wire \n1[12]_i_3__0_n_0 ;
  wire \n1[13]_i_2__0_n_0 ;
  wire \n1[13]_i_3__0_n_0 ;
  wire \n1[14]_i_2__0_n_0 ;
  wire \n1[14]_i_3__0_n_0 ;
  wire \n1[15]_i_2__0_n_0 ;
  wire \n1[15]_i_3__0_n_0 ;
  wire \n1[1]_i_2__0_n_0 ;
  wire \n1[1]_i_3__0_n_0 ;
  wire \n1[2]_i_2__0_n_0 ;
  wire \n1[2]_i_3__0_n_0 ;
  wire \n1[3]_i_2__0_n_0 ;
  wire \n1[3]_i_3__0_n_0 ;
  wire \n1[4]_i_2__0_n_0 ;
  wire \n1[4]_i_3__0_n_0 ;
  wire \n1[5]_i_2__0_n_0 ;
  wire \n1[5]_i_3__0_n_0 ;
  wire \n1[6]_i_2__0_n_0 ;
  wire \n1[6]_i_3__0_n_0 ;
  wire \n1[7]_i_2__0_n_0 ;
  wire \n1[7]_i_3__0_n_0 ;
  wire \n1[8]_i_2__0_n_0 ;
  wire \n1[8]_i_3__0_n_0 ;
  wire \n1[9]_i_2__0_n_0 ;
  wire \n1[9]_i_3__0_n_0 ;
  wire \n1_reg[0] ;
  wire [6:0]n2__0;
  wire \n3[6]_i_2__1_n_0 ;
  wire [6:0]n3_reg;
  wire n4;
  wire \n5[0]_i_2__1_n_0 ;
  wire [15:0]\n9_reg[0] ;
  wire n9m_reg_0_63_0_6_n_0;
  wire n9m_reg_0_63_0_6_n_1;
  wire n9m_reg_0_63_0_6_n_2;
  wire n9m_reg_0_63_0_6_n_3;
  wire n9m_reg_0_63_0_6_n_4;
  wire n9m_reg_0_63_0_6_n_5;
  wire n9m_reg_0_63_0_6_n_6;
  wire n9m_reg_0_63_14_20_n_0;
  wire n9m_reg_0_63_14_20_n_1;
  wire n9m_reg_0_63_14_20_n_2;
  wire n9m_reg_0_63_14_20_n_3;
  wire n9m_reg_0_63_14_20_n_4;
  wire n9m_reg_0_63_14_20_n_5;
  wire n9m_reg_0_63_14_20_n_6;
  wire n9m_reg_0_63_21_27_n_0;
  wire n9m_reg_0_63_21_27_n_1;
  wire n9m_reg_0_63_21_27_n_2;
  wire n9m_reg_0_63_21_27_n_3;
  wire n9m_reg_0_63_21_27_n_4;
  wire n9m_reg_0_63_21_27_n_5;
  wire n9m_reg_0_63_21_27_n_6;
  wire n9m_reg_0_63_28_31_n_0;
  wire n9m_reg_0_63_28_31_n_1;
  wire n9m_reg_0_63_28_31_n_2;
  wire n9m_reg_0_63_28_31_n_3;
  wire n9m_reg_0_63_7_13_n_0;
  wire n9m_reg_0_63_7_13_n_1;
  wire n9m_reg_0_63_7_13_n_2;
  wire n9m_reg_0_63_7_13_n_3;
  wire n9m_reg_0_63_7_13_n_4;
  wire n9m_reg_0_63_7_13_n_5;
  wire n9m_reg_0_63_7_13_n_6;
  wire n9m_reg_64_127_0_6_n_0;
  wire n9m_reg_64_127_0_6_n_1;
  wire n9m_reg_64_127_0_6_n_2;
  wire n9m_reg_64_127_0_6_n_3;
  wire n9m_reg_64_127_0_6_n_4;
  wire n9m_reg_64_127_0_6_n_5;
  wire n9m_reg_64_127_0_6_n_6;
  wire n9m_reg_64_127_14_20_n_0;
  wire n9m_reg_64_127_14_20_n_1;
  wire n9m_reg_64_127_14_20_n_2;
  wire n9m_reg_64_127_14_20_n_3;
  wire n9m_reg_64_127_14_20_n_4;
  wire n9m_reg_64_127_14_20_n_5;
  wire n9m_reg_64_127_14_20_n_6;
  wire n9m_reg_64_127_21_27_n_0;
  wire n9m_reg_64_127_21_27_n_1;
  wire n9m_reg_64_127_21_27_n_2;
  wire n9m_reg_64_127_21_27_n_3;
  wire n9m_reg_64_127_21_27_n_4;
  wire n9m_reg_64_127_21_27_n_5;
  wire n9m_reg_64_127_21_27_n_6;
  wire n9m_reg_64_127_28_31_n_0;
  wire n9m_reg_64_127_28_31_n_1;
  wire n9m_reg_64_127_28_31_n_2;
  wire n9m_reg_64_127_28_31_n_3;
  wire n9m_reg_64_127_7_13_n_0;
  wire n9m_reg_64_127_7_13_n_1;
  wire n9m_reg_64_127_7_13_n_2;
  wire n9m_reg_64_127_7_13_n_3;
  wire n9m_reg_64_127_7_13_n_4;
  wire n9m_reg_64_127_7_13_n_5;
  wire n9m_reg_64_127_7_13_n_6;
  wire rst_i;
  wire NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED;

  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39758 n11m_reg_0_63_0_6
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[0]),
        .DIB(i1[1]),
        .DIC(i1[2]),
        .DID(i1[3]),
        .DIE(i1[4]),
        .DIF(i1[5]),
        .DIG(i1[6]),
        .DIH(1'b0),
        .DOA(n11[0]),
        .DOB(n11[1]),
        .DOC(n11[2]),
        .DOD(n11[3]),
        .DOE(n11[4]),
        .DOF(n11[5]),
        .DOG(n11[6]),
        .DOH(NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39759 n11m_reg_0_63_14_20
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[0]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n11[14]),
        .DOB(n11[15]),
        .DOC(n11[16]),
        .DOD(n11[17]),
        .DOE(n11[18]),
        .DOF(n11[19]),
        .DOG(n11[20]),
        .DOH(NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39760 n11m_reg_0_63_21_27
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n11[21]),
        .DOB(n11[22]),
        .DOC(n11[23]),
        .DOD(n11[24]),
        .DOE(n11[25]),
        .DOF(n11[26]),
        .DOG(n11[27]),
        .DOH(NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39761 n11m_reg_0_63_28_31
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n11[28]),
        .DOB(n11[29]),
        .DOC(n11[30]),
        .DOD(n11[31]),
        .DOE(NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39762 n11m_reg_0_63_7_13
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[7]),
        .DIB(i1[22]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n11[7]),
        .DOB(n11[8]),
        .DOC(n11[9]),
        .DOD(n11[10]),
        .DOE(n11[11]),
        .DOF(n11[12]),
        .DOG(n11[13]),
        .DOH(NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[0]_i_1__0 
       (.I0(n11[0]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[0]_i_2__0_n_0 ),
        .I4(\n1[0]_i_3__0_n_0 ),
        .O(\n9_reg[0] [0]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[0]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_0),
        .O(\n1[0]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[0]_i_3__0 
       (.I0(n11[16]),
        .I1(n9m_reg_64_127_14_20_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[0]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[10]_i_1__0 
       (.I0(n11[10]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[10]_i_2__0_n_0 ),
        .I4(\n1[10]_i_3__0_n_0 ),
        .O(\n9_reg[0] [10]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[10]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_3),
        .O(\n1[10]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[10]_i_3__0 
       (.I0(n11[26]),
        .I1(n9m_reg_64_127_21_27_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[10]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[11]_i_1__0 
       (.I0(n11[11]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[11]_i_2__0_n_0 ),
        .I4(\n1[11]_i_3__0_n_0 ),
        .O(\n9_reg[0] [11]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[11]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_4),
        .O(\n1[11]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[11]_i_3__0 
       (.I0(n11[27]),
        .I1(n9m_reg_64_127_21_27_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[11]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[12]_i_1__0 
       (.I0(n11[12]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[12]_i_2__0_n_0 ),
        .I4(\n1[12]_i_3__0_n_0 ),
        .O(\n9_reg[0] [12]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[12]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_5),
        .O(\n1[12]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[12]_i_3__0 
       (.I0(n11[28]),
        .I1(n9m_reg_64_127_28_31_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[12]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[13]_i_1__0 
       (.I0(n11[13]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[13]_i_2__0_n_0 ),
        .I4(\n1[13]_i_3__0_n_0 ),
        .O(\n9_reg[0] [13]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[13]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_6),
        .O(\n1[13]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[13]_i_3__0 
       (.I0(n11[29]),
        .I1(n9m_reg_64_127_28_31_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[13]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[14]_i_1__0 
       (.I0(n11[14]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[14]_i_2__0_n_0 ),
        .I4(\n1[14]_i_3__0_n_0 ),
        .O(\n9_reg[0] [14]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[14]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_0),
        .O(\n1[14]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[14]_i_3__0 
       (.I0(n11[30]),
        .I1(n9m_reg_64_127_28_31_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[14]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[15]_i_1__0 
       (.I0(n11[15]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[15]_i_2__0_n_0 ),
        .I4(\n1[15]_i_3__0_n_0 ),
        .O(\n9_reg[0] [15]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[15]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_1),
        .O(\n1[15]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[15]_i_3__0 
       (.I0(n11[31]),
        .I1(n9m_reg_64_127_28_31_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[15]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[1]_i_1__0 
       (.I0(n11[1]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[1]_i_2__0_n_0 ),
        .I4(\n1[1]_i_3__0_n_0 ),
        .O(\n9_reg[0] [1]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[1]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_1),
        .O(\n1[1]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[1]_i_3__0 
       (.I0(n11[17]),
        .I1(n9m_reg_64_127_14_20_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[1]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[2]_i_1__0 
       (.I0(n11[2]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[2]_i_2__0_n_0 ),
        .I4(\n1[2]_i_3__0_n_0 ),
        .O(\n9_reg[0] [2]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[2]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_2),
        .O(\n1[2]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[2]_i_3__0 
       (.I0(n11[18]),
        .I1(n9m_reg_64_127_14_20_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[2]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[3]_i_1__0 
       (.I0(n11[3]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[3]_i_2__0_n_0 ),
        .I4(\n1[3]_i_3__0_n_0 ),
        .O(\n9_reg[0] [3]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[3]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_3),
        .O(\n1[3]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[3]_i_3__0 
       (.I0(n11[19]),
        .I1(n9m_reg_64_127_14_20_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[3]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[4]_i_1__0 
       (.I0(n11[4]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[4]_i_2__0_n_0 ),
        .I4(\n1[4]_i_3__0_n_0 ),
        .O(\n9_reg[0] [4]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[4]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_4),
        .O(\n1[4]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[4]_i_3__0 
       (.I0(n11[20]),
        .I1(n9m_reg_64_127_14_20_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[4]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[5]_i_1__0 
       (.I0(n11[5]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[5]_i_2__0_n_0 ),
        .I4(\n1[5]_i_3__0_n_0 ),
        .O(\n9_reg[0] [5]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[5]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_5),
        .O(\n1[5]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[5]_i_3__0 
       (.I0(n11[21]),
        .I1(n9m_reg_64_127_21_27_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[5]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[6]_i_1__0 
       (.I0(n11[6]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[6]_i_2__0_n_0 ),
        .I4(\n1[6]_i_3__0_n_0 ),
        .O(\n9_reg[0] [6]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[6]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_6),
        .O(\n1[6]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[6]_i_3__0 
       (.I0(n11[22]),
        .I1(n9m_reg_64_127_21_27_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[6]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[7]_i_1__0 
       (.I0(n11[7]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[7]_i_2__0_n_0 ),
        .I4(\n1[7]_i_3__0_n_0 ),
        .O(\n9_reg[0] [7]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[7]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_0),
        .O(\n1[7]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[7]_i_3__0 
       (.I0(n11[23]),
        .I1(n9m_reg_64_127_21_27_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[7]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[8]_i_1__0 
       (.I0(n11[8]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[8]_i_2__0_n_0 ),
        .I4(\n1[8]_i_3__0_n_0 ),
        .O(\n9_reg[0] [8]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[8]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_1),
        .O(\n1[8]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[8]_i_3__0 
       (.I0(n11[24]),
        .I1(n9m_reg_64_127_21_27_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[8]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[9]_i_1__0 
       (.I0(n11[9]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[9]_i_2__0_n_0 ),
        .I4(\n1[9]_i_3__0_n_0 ),
        .O(\n9_reg[0] [9]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[9]_i_2__0 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_2),
        .O(\n1[9]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[9]_i_3__0 
       (.I0(n11[25]),
        .I1(n9m_reg_64_127_21_27_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[9]_i_3__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__3 
       (.I0(n3_reg[0]),
        .O(n2__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__3 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__3 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__3 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__3 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__0[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__3 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__0[5]));
  LUT3 #(
    .INIT(8'hD2)) 
    \n3[6]_i_1__1 
       (.I0(n3_reg[5]),
        .I1(\n3[6]_i_2__1_n_0 ),
        .I2(n3_reg[6]),
        .O(n2__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \n3[6]_i_2__1 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(\n3[6]_i_2__1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[6]),
        .Q(n3_reg[6]),
        .R(rst_i));
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \n5[0]_i_1__1 
       (.I0(n3_reg[0]),
        .I1(\n5[0]_i_2__1_n_0 ),
        .I2(i8),
        .O(n4));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \n5[0]_i_2__1 
       (.I0(n3_reg[3]),
        .I1(n3_reg[4]),
        .I2(n3_reg[1]),
        .I3(n3_reg[2]),
        .I4(n3_reg[6]),
        .I5(n3_reg[5]),
        .O(\n5[0]_i_2__1_n_0 ));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[6]),
        .Q(n11a[6]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39763 n9m_reg_0_63_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[0]),
        .DIB(i1[1]),
        .DIC(i1[2]),
        .DID(i1[3]),
        .DIE(i1[4]),
        .DIF(i1[5]),
        .DIG(i1[6]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_0_6_n_0),
        .DOB(n9m_reg_0_63_0_6_n_1),
        .DOC(n9m_reg_0_63_0_6_n_2),
        .DOD(n9m_reg_0_63_0_6_n_3),
        .DOE(n9m_reg_0_63_0_6_n_4),
        .DOF(n9m_reg_0_63_0_6_n_5),
        .DOG(n9m_reg_0_63_0_6_n_6),
        .DOH(NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39764 n9m_reg_0_63_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[0]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_14_20_n_0),
        .DOB(n9m_reg_0_63_14_20_n_1),
        .DOC(n9m_reg_0_63_14_20_n_2),
        .DOD(n9m_reg_0_63_14_20_n_3),
        .DOE(n9m_reg_0_63_14_20_n_4),
        .DOF(n9m_reg_0_63_14_20_n_5),
        .DOG(n9m_reg_0_63_14_20_n_6),
        .DOH(NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39765 n9m_reg_0_63_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_21_27_n_0),
        .DOB(n9m_reg_0_63_21_27_n_1),
        .DOC(n9m_reg_0_63_21_27_n_2),
        .DOD(n9m_reg_0_63_21_27_n_3),
        .DOE(n9m_reg_0_63_21_27_n_4),
        .DOF(n9m_reg_0_63_21_27_n_5),
        .DOG(n9m_reg_0_63_21_27_n_6),
        .DOH(NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39766 n9m_reg_0_63_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_28_31_n_0),
        .DOB(n9m_reg_0_63_28_31_n_1),
        .DOC(n9m_reg_0_63_28_31_n_2),
        .DOD(n9m_reg_0_63_28_31_n_3),
        .DOE(NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39767 n9m_reg_0_63_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[7]),
        .DIB(i1[22]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_7_13_n_0),
        .DOB(n9m_reg_0_63_7_13_n_1),
        .DOC(n9m_reg_0_63_7_13_n_2),
        .DOD(n9m_reg_0_63_7_13_n_3),
        .DOE(n9m_reg_0_63_7_13_n_4),
        .DOF(n9m_reg_0_63_7_13_n_5),
        .DOG(n9m_reg_0_63_7_13_n_6),
        .DOH(NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39768 n9m_reg_64_127_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[0]),
        .DIB(i1[1]),
        .DIC(i1[2]),
        .DID(i1[3]),
        .DIE(i1[4]),
        .DIF(i1[5]),
        .DIG(i1[6]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_0_6_n_0),
        .DOB(n9m_reg_64_127_0_6_n_1),
        .DOC(n9m_reg_64_127_0_6_n_2),
        .DOD(n9m_reg_64_127_0_6_n_3),
        .DOE(n9m_reg_64_127_0_6_n_4),
        .DOF(n9m_reg_64_127_0_6_n_5),
        .DOG(n9m_reg_64_127_0_6_n_6),
        .DOH(NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39769 n9m_reg_64_127_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[0]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_14_20_n_0),
        .DOB(n9m_reg_64_127_14_20_n_1),
        .DOC(n9m_reg_64_127_14_20_n_2),
        .DOD(n9m_reg_64_127_14_20_n_3),
        .DOE(n9m_reg_64_127_14_20_n_4),
        .DOF(n9m_reg_64_127_14_20_n_5),
        .DOG(n9m_reg_64_127_14_20_n_6),
        .DOH(NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39770 n9m_reg_64_127_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_21_27_n_0),
        .DOB(n9m_reg_64_127_21_27_n_1),
        .DOC(n9m_reg_64_127_21_27_n_2),
        .DOD(n9m_reg_64_127_21_27_n_3),
        .DOE(n9m_reg_64_127_21_27_n_4),
        .DOF(n9m_reg_64_127_21_27_n_5),
        .DOG(n9m_reg_64_127_21_27_n_6),
        .DOH(NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39771 n9m_reg_64_127_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_28_31_n_0),
        .DOB(n9m_reg_64_127_28_31_n_1),
        .DOC(n9m_reg_64_127_28_31_n_2),
        .DOD(n9m_reg_64_127_28_31_n_3),
        .DOE(NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39772 n9m_reg_64_127_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[7]),
        .DIB(i1[22]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_7_13_n_0),
        .DOB(n9m_reg_64_127_7_13_n_1),
        .DOC(n9m_reg_64_127_7_13_n_2),
        .DOD(n9m_reg_64_127_7_13_n_3),
        .DOE(n9m_reg_64_127_7_13_n_4),
        .DOF(n9m_reg_64_127_7_13_n_5),
        .DOG(n9m_reg_64_127_7_13_n_6),
        .DOH(NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_26" *) 
module switch_elements_cf_fft_512_8_26_18
   (\n9_reg[0] ,
    n4,
    \n1_reg[0] ,
    i8,
    rst_i,
    enable_i,
    clk_i,
    i1);
  output [15:0]\n9_reg[0] ;
  output n4;
  input \n1_reg[0] ;
  input [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [31:0]n11;
  wire [6:0]n11a;
  wire [5:0]n11a__0;
  wire \n1[0]_i_2_n_0 ;
  wire \n1[0]_i_3_n_0 ;
  wire \n1[10]_i_2_n_0 ;
  wire \n1[10]_i_3_n_0 ;
  wire \n1[11]_i_2_n_0 ;
  wire \n1[11]_i_3_n_0 ;
  wire \n1[12]_i_2_n_0 ;
  wire \n1[12]_i_3_n_0 ;
  wire \n1[13]_i_2_n_0 ;
  wire \n1[13]_i_3_n_0 ;
  wire \n1[14]_i_2_n_0 ;
  wire \n1[14]_i_3_n_0 ;
  wire \n1[15]_i_2_n_0 ;
  wire \n1[15]_i_3_n_0 ;
  wire \n1[1]_i_2_n_0 ;
  wire \n1[1]_i_3_n_0 ;
  wire \n1[2]_i_2_n_0 ;
  wire \n1[2]_i_3_n_0 ;
  wire \n1[3]_i_2_n_0 ;
  wire \n1[3]_i_3_n_0 ;
  wire \n1[4]_i_2_n_0 ;
  wire \n1[4]_i_3_n_0 ;
  wire \n1[5]_i_2_n_0 ;
  wire \n1[5]_i_3_n_0 ;
  wire \n1[6]_i_2_n_0 ;
  wire \n1[6]_i_3_n_0 ;
  wire \n1[7]_i_2_n_0 ;
  wire \n1[7]_i_3_n_0 ;
  wire \n1[8]_i_2_n_0 ;
  wire \n1[8]_i_3_n_0 ;
  wire \n1[9]_i_2_n_0 ;
  wire \n1[9]_i_3_n_0 ;
  wire \n1_reg[0] ;
  wire [6:0]n2__0;
  wire \n3[6]_i_2__0_n_0 ;
  wire [6:0]n3_reg;
  wire n4;
  wire \n5[0]_i_2__0_n_0 ;
  wire [15:0]\n9_reg[0] ;
  wire n9m_reg_0_63_0_6_n_0;
  wire n9m_reg_0_63_0_6_n_1;
  wire n9m_reg_0_63_0_6_n_2;
  wire n9m_reg_0_63_0_6_n_3;
  wire n9m_reg_0_63_0_6_n_4;
  wire n9m_reg_0_63_0_6_n_5;
  wire n9m_reg_0_63_0_6_n_6;
  wire n9m_reg_0_63_14_20_n_0;
  wire n9m_reg_0_63_14_20_n_1;
  wire n9m_reg_0_63_14_20_n_2;
  wire n9m_reg_0_63_14_20_n_3;
  wire n9m_reg_0_63_14_20_n_4;
  wire n9m_reg_0_63_14_20_n_5;
  wire n9m_reg_0_63_14_20_n_6;
  wire n9m_reg_0_63_21_27_n_0;
  wire n9m_reg_0_63_21_27_n_1;
  wire n9m_reg_0_63_21_27_n_2;
  wire n9m_reg_0_63_21_27_n_3;
  wire n9m_reg_0_63_21_27_n_4;
  wire n9m_reg_0_63_21_27_n_5;
  wire n9m_reg_0_63_21_27_n_6;
  wire n9m_reg_0_63_28_31_n_0;
  wire n9m_reg_0_63_28_31_n_1;
  wire n9m_reg_0_63_28_31_n_2;
  wire n9m_reg_0_63_28_31_n_3;
  wire n9m_reg_0_63_7_13_n_0;
  wire n9m_reg_0_63_7_13_n_1;
  wire n9m_reg_0_63_7_13_n_2;
  wire n9m_reg_0_63_7_13_n_3;
  wire n9m_reg_0_63_7_13_n_4;
  wire n9m_reg_0_63_7_13_n_5;
  wire n9m_reg_0_63_7_13_n_6;
  wire n9m_reg_64_127_0_6_n_0;
  wire n9m_reg_64_127_0_6_n_1;
  wire n9m_reg_64_127_0_6_n_2;
  wire n9m_reg_64_127_0_6_n_3;
  wire n9m_reg_64_127_0_6_n_4;
  wire n9m_reg_64_127_0_6_n_5;
  wire n9m_reg_64_127_0_6_n_6;
  wire n9m_reg_64_127_14_20_n_0;
  wire n9m_reg_64_127_14_20_n_1;
  wire n9m_reg_64_127_14_20_n_2;
  wire n9m_reg_64_127_14_20_n_3;
  wire n9m_reg_64_127_14_20_n_4;
  wire n9m_reg_64_127_14_20_n_5;
  wire n9m_reg_64_127_14_20_n_6;
  wire n9m_reg_64_127_21_27_n_0;
  wire n9m_reg_64_127_21_27_n_1;
  wire n9m_reg_64_127_21_27_n_2;
  wire n9m_reg_64_127_21_27_n_3;
  wire n9m_reg_64_127_21_27_n_4;
  wire n9m_reg_64_127_21_27_n_5;
  wire n9m_reg_64_127_21_27_n_6;
  wire n9m_reg_64_127_28_31_n_0;
  wire n9m_reg_64_127_28_31_n_1;
  wire n9m_reg_64_127_28_31_n_2;
  wire n9m_reg_64_127_28_31_n_3;
  wire n9m_reg_64_127_7_13_n_0;
  wire n9m_reg_64_127_7_13_n_1;
  wire n9m_reg_64_127_7_13_n_2;
  wire n9m_reg_64_127_7_13_n_3;
  wire n9m_reg_64_127_7_13_n_4;
  wire n9m_reg_64_127_7_13_n_5;
  wire n9m_reg_64_127_7_13_n_6;
  wire rst_i;
  wire NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED;

  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39743 n11m_reg_0_63_0_6
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[14]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n11[0]),
        .DOB(n11[1]),
        .DOC(n11[2]),
        .DOD(n11[3]),
        .DOE(n11[4]),
        .DOF(n11[5]),
        .DOG(n11[6]),
        .DOH(NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39744 n11m_reg_0_63_14_20
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[12]),
        .DIB(i1[13]),
        .DIC(i1[14]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n11[14]),
        .DOB(n11[15]),
        .DOC(n11[16]),
        .DOD(n11[17]),
        .DOE(n11[18]),
        .DOF(n11[19]),
        .DOG(n11[20]),
        .DOH(NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39745 n11m_reg_0_63_21_27
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n11[21]),
        .DOB(n11[22]),
        .DOC(n11[23]),
        .DOD(n11[24]),
        .DOE(n11[25]),
        .DOF(n11[26]),
        .DOG(n11[27]),
        .DOH(NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39746 n11m_reg_0_63_28_31
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n11[28]),
        .DOB(n11[29]),
        .DOC(n11[30]),
        .DOD(n11[31]),
        .DOE(NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39747 n11m_reg_0_63_7_13
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[22]),
        .DIC(i1[7]),
        .DID(i1[8]),
        .DIE(i1[9]),
        .DIF(i1[10]),
        .DIG(i1[11]),
        .DIH(1'b0),
        .DOA(n11[7]),
        .DOB(n11[8]),
        .DOC(n11[9]),
        .DOD(n11[10]),
        .DOE(n11[11]),
        .DOF(n11[12]),
        .DOG(n11[13]),
        .DOH(NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[0]_i_1 
       (.I0(n11[0]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[0]_i_2_n_0 ),
        .I4(\n1[0]_i_3_n_0 ),
        .O(\n9_reg[0] [0]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[0]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_0),
        .O(\n1[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[0]_i_3 
       (.I0(n11[16]),
        .I1(n9m_reg_64_127_14_20_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[0]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[10]_i_1 
       (.I0(n11[10]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[10]_i_2_n_0 ),
        .I4(\n1[10]_i_3_n_0 ),
        .O(\n9_reg[0] [10]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[10]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_3),
        .O(\n1[10]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[10]_i_3 
       (.I0(n11[26]),
        .I1(n9m_reg_64_127_21_27_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[10]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[11]_i_1 
       (.I0(n11[11]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[11]_i_2_n_0 ),
        .I4(\n1[11]_i_3_n_0 ),
        .O(\n9_reg[0] [11]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[11]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_4),
        .O(\n1[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[11]_i_3 
       (.I0(n11[27]),
        .I1(n9m_reg_64_127_21_27_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[11]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[12]_i_1 
       (.I0(n11[12]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[12]_i_2_n_0 ),
        .I4(\n1[12]_i_3_n_0 ),
        .O(\n9_reg[0] [12]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[12]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_5),
        .O(\n1[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[12]_i_3 
       (.I0(n11[28]),
        .I1(n9m_reg_64_127_28_31_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[12]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[13]_i_1 
       (.I0(n11[13]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[13]_i_2_n_0 ),
        .I4(\n1[13]_i_3_n_0 ),
        .O(\n9_reg[0] [13]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[13]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_6),
        .O(\n1[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[13]_i_3 
       (.I0(n11[29]),
        .I1(n9m_reg_64_127_28_31_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[13]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[14]_i_1 
       (.I0(n11[14]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[14]_i_2_n_0 ),
        .I4(\n1[14]_i_3_n_0 ),
        .O(\n9_reg[0] [14]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[14]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_0),
        .O(\n1[14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[14]_i_3 
       (.I0(n11[30]),
        .I1(n9m_reg_64_127_28_31_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[14]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[15]_i_1 
       (.I0(n11[15]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[15]_i_2_n_0 ),
        .I4(\n1[15]_i_3_n_0 ),
        .O(\n9_reg[0] [15]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[15]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_1),
        .O(\n1[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[15]_i_3 
       (.I0(n11[31]),
        .I1(n9m_reg_64_127_28_31_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[15]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[1]_i_1 
       (.I0(n11[1]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[1]_i_2_n_0 ),
        .I4(\n1[1]_i_3_n_0 ),
        .O(\n9_reg[0] [1]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[1]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_1),
        .O(\n1[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[1]_i_3 
       (.I0(n11[17]),
        .I1(n9m_reg_64_127_14_20_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[1]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[2]_i_1 
       (.I0(n11[2]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[2]_i_2_n_0 ),
        .I4(\n1[2]_i_3_n_0 ),
        .O(\n9_reg[0] [2]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[2]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_2),
        .O(\n1[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[2]_i_3 
       (.I0(n11[18]),
        .I1(n9m_reg_64_127_14_20_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[2]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[3]_i_1 
       (.I0(n11[3]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[3]_i_2_n_0 ),
        .I4(\n1[3]_i_3_n_0 ),
        .O(\n9_reg[0] [3]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[3]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_3),
        .O(\n1[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[3]_i_3 
       (.I0(n11[19]),
        .I1(n9m_reg_64_127_14_20_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[3]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[4]_i_1 
       (.I0(n11[4]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[4]_i_2_n_0 ),
        .I4(\n1[4]_i_3_n_0 ),
        .O(\n9_reg[0] [4]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[4]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_4),
        .O(\n1[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[4]_i_3 
       (.I0(n11[20]),
        .I1(n9m_reg_64_127_14_20_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[4]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[5]_i_1 
       (.I0(n11[5]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[5]_i_2_n_0 ),
        .I4(\n1[5]_i_3_n_0 ),
        .O(\n9_reg[0] [5]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[5]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_5),
        .O(\n1[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[5]_i_3 
       (.I0(n11[21]),
        .I1(n9m_reg_64_127_21_27_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[5]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[6]_i_1 
       (.I0(n11[6]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[6]_i_2_n_0 ),
        .I4(\n1[6]_i_3_n_0 ),
        .O(\n9_reg[0] [6]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[6]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_6),
        .O(\n1[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[6]_i_3 
       (.I0(n11[22]),
        .I1(n9m_reg_64_127_21_27_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[7]_i_1 
       (.I0(n11[7]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[7]_i_2_n_0 ),
        .I4(\n1[7]_i_3_n_0 ),
        .O(\n9_reg[0] [7]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[7]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_0),
        .O(\n1[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[7]_i_3 
       (.I0(n11[23]),
        .I1(n9m_reg_64_127_21_27_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[7]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[8]_i_1 
       (.I0(n11[8]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[8]_i_2_n_0 ),
        .I4(\n1[8]_i_3_n_0 ),
        .O(\n9_reg[0] [8]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[8]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_1),
        .O(\n1[8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[8]_i_3 
       (.I0(n11[24]),
        .I1(n9m_reg_64_127_21_27_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[8]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[9]_i_1 
       (.I0(n11[9]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[9]_i_2_n_0 ),
        .I4(\n1[9]_i_3_n_0 ),
        .O(\n9_reg[0] [9]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[9]_i_2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_2),
        .O(\n1[9]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[9]_i_3 
       (.I0(n11[25]),
        .I1(n9m_reg_64_127_21_27_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[9]_i_3_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__1 
       (.I0(n3_reg[0]),
        .O(n2__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__1 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__1 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__1 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__1 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__0[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__1 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__0[5]));
  LUT3 #(
    .INIT(8'hD2)) 
    \n3[6]_i_1__0 
       (.I0(n3_reg[5]),
        .I1(\n3[6]_i_2__0_n_0 ),
        .I2(n3_reg[6]),
        .O(n2__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \n3[6]_i_2__0 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(\n3[6]_i_2__0_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[6]),
        .Q(n3_reg[6]),
        .R(rst_i));
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \n5[0]_i_1__0 
       (.I0(n3_reg[0]),
        .I1(\n5[0]_i_2__0_n_0 ),
        .I2(i8),
        .O(n4));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \n5[0]_i_2__0 
       (.I0(n3_reg[3]),
        .I1(n3_reg[4]),
        .I2(n3_reg[1]),
        .I3(n3_reg[2]),
        .I4(n3_reg[6]),
        .I5(n3_reg[5]),
        .O(\n5[0]_i_2__0_n_0 ));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[6]),
        .Q(n11a[6]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39748 n9m_reg_0_63_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[14]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_0_6_n_0),
        .DOB(n9m_reg_0_63_0_6_n_1),
        .DOC(n9m_reg_0_63_0_6_n_2),
        .DOD(n9m_reg_0_63_0_6_n_3),
        .DOE(n9m_reg_0_63_0_6_n_4),
        .DOF(n9m_reg_0_63_0_6_n_5),
        .DOG(n9m_reg_0_63_0_6_n_6),
        .DOH(NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39749 n9m_reg_0_63_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[12]),
        .DIB(i1[13]),
        .DIC(i1[14]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_14_20_n_0),
        .DOB(n9m_reg_0_63_14_20_n_1),
        .DOC(n9m_reg_0_63_14_20_n_2),
        .DOD(n9m_reg_0_63_14_20_n_3),
        .DOE(n9m_reg_0_63_14_20_n_4),
        .DOF(n9m_reg_0_63_14_20_n_5),
        .DOG(n9m_reg_0_63_14_20_n_6),
        .DOH(NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39750 n9m_reg_0_63_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_21_27_n_0),
        .DOB(n9m_reg_0_63_21_27_n_1),
        .DOC(n9m_reg_0_63_21_27_n_2),
        .DOD(n9m_reg_0_63_21_27_n_3),
        .DOE(n9m_reg_0_63_21_27_n_4),
        .DOF(n9m_reg_0_63_21_27_n_5),
        .DOG(n9m_reg_0_63_21_27_n_6),
        .DOH(NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39751 n9m_reg_0_63_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_28_31_n_0),
        .DOB(n9m_reg_0_63_28_31_n_1),
        .DOC(n9m_reg_0_63_28_31_n_2),
        .DOD(n9m_reg_0_63_28_31_n_3),
        .DOE(NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39752 n9m_reg_0_63_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[22]),
        .DIC(i1[7]),
        .DID(i1[8]),
        .DIE(i1[9]),
        .DIF(i1[10]),
        .DIG(i1[11]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_7_13_n_0),
        .DOB(n9m_reg_0_63_7_13_n_1),
        .DOC(n9m_reg_0_63_7_13_n_2),
        .DOD(n9m_reg_0_63_7_13_n_3),
        .DOE(n9m_reg_0_63_7_13_n_4),
        .DOF(n9m_reg_0_63_7_13_n_5),
        .DOG(n9m_reg_0_63_7_13_n_6),
        .DOH(NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39753 n9m_reg_64_127_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[14]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_0_6_n_0),
        .DOB(n9m_reg_64_127_0_6_n_1),
        .DOC(n9m_reg_64_127_0_6_n_2),
        .DOD(n9m_reg_64_127_0_6_n_3),
        .DOE(n9m_reg_64_127_0_6_n_4),
        .DOF(n9m_reg_64_127_0_6_n_5),
        .DOG(n9m_reg_64_127_0_6_n_6),
        .DOH(NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39754 n9m_reg_64_127_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[12]),
        .DIB(i1[13]),
        .DIC(i1[14]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_14_20_n_0),
        .DOB(n9m_reg_64_127_14_20_n_1),
        .DOC(n9m_reg_64_127_14_20_n_2),
        .DOD(n9m_reg_64_127_14_20_n_3),
        .DOE(n9m_reg_64_127_14_20_n_4),
        .DOF(n9m_reg_64_127_14_20_n_5),
        .DOG(n9m_reg_64_127_14_20_n_6),
        .DOH(NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39755 n9m_reg_64_127_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_21_27_n_0),
        .DOB(n9m_reg_64_127_21_27_n_1),
        .DOC(n9m_reg_64_127_21_27_n_2),
        .DOD(n9m_reg_64_127_21_27_n_3),
        .DOE(n9m_reg_64_127_21_27_n_4),
        .DOF(n9m_reg_64_127_21_27_n_5),
        .DOG(n9m_reg_64_127_21_27_n_6),
        .DOH(NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39756 n9m_reg_64_127_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_28_31_n_0),
        .DOB(n9m_reg_64_127_28_31_n_1),
        .DOC(n9m_reg_64_127_28_31_n_2),
        .DOD(n9m_reg_64_127_28_31_n_3),
        .DOE(NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39757 n9m_reg_64_127_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[22]),
        .DIC(i1[7]),
        .DID(i1[8]),
        .DIE(i1[9]),
        .DIF(i1[10]),
        .DIG(i1[11]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_7_13_n_0),
        .DOB(n9m_reg_64_127_7_13_n_1),
        .DOC(n9m_reg_64_127_7_13_n_2),
        .DOD(n9m_reg_64_127_7_13_n_3),
        .DOE(n9m_reg_64_127_7_13_n_4),
        .DOF(n9m_reg_64_127_7_13_n_5),
        .DOG(n9m_reg_64_127_7_13_n_6),
        .DOH(NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_26" *) 
module switch_elements_cf_fft_512_8_26_2
   (\n9_reg[0] ,
    n4,
    \n1_reg[0] ,
    i8,
    rst_i,
    enable_i,
    clk_i,
    i1);
  output [15:0]\n9_reg[0] ;
  output n4;
  input \n1_reg[0] ;
  input [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [31:0]n11;
  wire [6:0]n11a;
  wire [5:0]n11a__0;
  wire \n1[0]_i_2__4_n_0 ;
  wire \n1[0]_i_3__4_n_0 ;
  wire \n1[10]_i_2__4_n_0 ;
  wire \n1[10]_i_3__4_n_0 ;
  wire \n1[11]_i_2__4_n_0 ;
  wire \n1[11]_i_3__4_n_0 ;
  wire \n1[12]_i_2__4_n_0 ;
  wire \n1[12]_i_3__4_n_0 ;
  wire \n1[13]_i_2__4_n_0 ;
  wire \n1[13]_i_3__4_n_0 ;
  wire \n1[14]_i_2__4_n_0 ;
  wire \n1[14]_i_3__4_n_0 ;
  wire \n1[15]_i_2__4_n_0 ;
  wire \n1[15]_i_3__4_n_0 ;
  wire \n1[1]_i_2__4_n_0 ;
  wire \n1[1]_i_3__4_n_0 ;
  wire \n1[2]_i_2__4_n_0 ;
  wire \n1[2]_i_3__4_n_0 ;
  wire \n1[3]_i_2__4_n_0 ;
  wire \n1[3]_i_3__4_n_0 ;
  wire \n1[4]_i_2__4_n_0 ;
  wire \n1[4]_i_3__4_n_0 ;
  wire \n1[5]_i_2__4_n_0 ;
  wire \n1[5]_i_3__4_n_0 ;
  wire \n1[6]_i_2__4_n_0 ;
  wire \n1[6]_i_3__4_n_0 ;
  wire \n1[7]_i_2__4_n_0 ;
  wire \n1[7]_i_3__4_n_0 ;
  wire \n1[8]_i_2__4_n_0 ;
  wire \n1[8]_i_3__4_n_0 ;
  wire \n1[9]_i_2__4_n_0 ;
  wire \n1[9]_i_3__4_n_0 ;
  wire \n1_reg[0] ;
  wire [6:0]n2__0;
  wire \n3[6]_i_2__5_n_0 ;
  wire [6:0]n3_reg;
  wire n4;
  wire \n5[0]_i_2__5_n_0 ;
  wire [15:0]\n9_reg[0] ;
  wire n9m_reg_0_63_0_6_n_0;
  wire n9m_reg_0_63_0_6_n_1;
  wire n9m_reg_0_63_0_6_n_2;
  wire n9m_reg_0_63_0_6_n_3;
  wire n9m_reg_0_63_0_6_n_4;
  wire n9m_reg_0_63_0_6_n_5;
  wire n9m_reg_0_63_0_6_n_6;
  wire n9m_reg_0_63_14_20_n_0;
  wire n9m_reg_0_63_14_20_n_1;
  wire n9m_reg_0_63_14_20_n_2;
  wire n9m_reg_0_63_14_20_n_3;
  wire n9m_reg_0_63_14_20_n_4;
  wire n9m_reg_0_63_14_20_n_5;
  wire n9m_reg_0_63_14_20_n_6;
  wire n9m_reg_0_63_21_27_n_0;
  wire n9m_reg_0_63_21_27_n_1;
  wire n9m_reg_0_63_21_27_n_2;
  wire n9m_reg_0_63_21_27_n_3;
  wire n9m_reg_0_63_21_27_n_4;
  wire n9m_reg_0_63_21_27_n_5;
  wire n9m_reg_0_63_21_27_n_6;
  wire n9m_reg_0_63_28_31_n_0;
  wire n9m_reg_0_63_28_31_n_1;
  wire n9m_reg_0_63_28_31_n_2;
  wire n9m_reg_0_63_28_31_n_3;
  wire n9m_reg_0_63_7_13_n_0;
  wire n9m_reg_0_63_7_13_n_1;
  wire n9m_reg_0_63_7_13_n_2;
  wire n9m_reg_0_63_7_13_n_3;
  wire n9m_reg_0_63_7_13_n_4;
  wire n9m_reg_0_63_7_13_n_5;
  wire n9m_reg_0_63_7_13_n_6;
  wire n9m_reg_64_127_0_6_n_0;
  wire n9m_reg_64_127_0_6_n_1;
  wire n9m_reg_64_127_0_6_n_2;
  wire n9m_reg_64_127_0_6_n_3;
  wire n9m_reg_64_127_0_6_n_4;
  wire n9m_reg_64_127_0_6_n_5;
  wire n9m_reg_64_127_0_6_n_6;
  wire n9m_reg_64_127_14_20_n_0;
  wire n9m_reg_64_127_14_20_n_1;
  wire n9m_reg_64_127_14_20_n_2;
  wire n9m_reg_64_127_14_20_n_3;
  wire n9m_reg_64_127_14_20_n_4;
  wire n9m_reg_64_127_14_20_n_5;
  wire n9m_reg_64_127_14_20_n_6;
  wire n9m_reg_64_127_21_27_n_0;
  wire n9m_reg_64_127_21_27_n_1;
  wire n9m_reg_64_127_21_27_n_2;
  wire n9m_reg_64_127_21_27_n_3;
  wire n9m_reg_64_127_21_27_n_4;
  wire n9m_reg_64_127_21_27_n_5;
  wire n9m_reg_64_127_21_27_n_6;
  wire n9m_reg_64_127_28_31_n_0;
  wire n9m_reg_64_127_28_31_n_1;
  wire n9m_reg_64_127_28_31_n_2;
  wire n9m_reg_64_127_28_31_n_3;
  wire n9m_reg_64_127_7_13_n_0;
  wire n9m_reg_64_127_7_13_n_1;
  wire n9m_reg_64_127_7_13_n_2;
  wire n9m_reg_64_127_7_13_n_3;
  wire n9m_reg_64_127_7_13_n_4;
  wire n9m_reg_64_127_7_13_n_5;
  wire n9m_reg_64_127_7_13_n_6;
  wire rst_i;
  wire NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED;

  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39858 n11m_reg_0_63_0_6
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n11[0]),
        .DOB(n11[1]),
        .DOC(n11[2]),
        .DOD(n11[3]),
        .DOE(n11[4]),
        .DOF(n11[5]),
        .DOG(n11[6]),
        .DOH(NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39859 n11m_reg_0_63_14_20
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n11[14]),
        .DOB(n11[15]),
        .DOC(n11[16]),
        .DOD(n11[17]),
        .DOE(n11[18]),
        .DOF(n11[19]),
        .DOG(n11[20]),
        .DOH(NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39860 n11m_reg_0_63_21_27
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n11[21]),
        .DOB(n11[22]),
        .DOC(n11[23]),
        .DOD(n11[24]),
        .DOE(n11[25]),
        .DOF(n11[26]),
        .DOG(n11[27]),
        .DOH(NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39861 n11m_reg_0_63_28_31
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n11[28]),
        .DOB(n11[29]),
        .DOC(n11[30]),
        .DOD(n11[31]),
        .DOE(NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39862 n11m_reg_0_63_7_13
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n11[7]),
        .DOB(n11[8]),
        .DOC(n11[9]),
        .DOD(n11[10]),
        .DOE(n11[11]),
        .DOF(n11[12]),
        .DOG(n11[13]),
        .DOH(NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[0]_i_1__4 
       (.I0(n11[0]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[0]_i_2__4_n_0 ),
        .I4(\n1[0]_i_3__4_n_0 ),
        .O(\n9_reg[0] [0]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[0]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_0),
        .O(\n1[0]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[0]_i_3__4 
       (.I0(n11[16]),
        .I1(n9m_reg_64_127_14_20_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[0]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[10]_i_1__4 
       (.I0(n11[10]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[10]_i_2__4_n_0 ),
        .I4(\n1[10]_i_3__4_n_0 ),
        .O(\n9_reg[0] [10]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[10]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_3),
        .O(\n1[10]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[10]_i_3__4 
       (.I0(n11[26]),
        .I1(n9m_reg_64_127_21_27_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[10]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[11]_i_1__4 
       (.I0(n11[11]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[11]_i_2__4_n_0 ),
        .I4(\n1[11]_i_3__4_n_0 ),
        .O(\n9_reg[0] [11]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[11]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_4),
        .O(\n1[11]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[11]_i_3__4 
       (.I0(n11[27]),
        .I1(n9m_reg_64_127_21_27_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[11]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[12]_i_1__4 
       (.I0(n11[12]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[12]_i_2__4_n_0 ),
        .I4(\n1[12]_i_3__4_n_0 ),
        .O(\n9_reg[0] [12]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[12]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_5),
        .O(\n1[12]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[12]_i_3__4 
       (.I0(n11[28]),
        .I1(n9m_reg_64_127_28_31_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[12]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[13]_i_1__4 
       (.I0(n11[13]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[13]_i_2__4_n_0 ),
        .I4(\n1[13]_i_3__4_n_0 ),
        .O(\n9_reg[0] [13]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[13]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_6),
        .O(\n1[13]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[13]_i_3__4 
       (.I0(n11[29]),
        .I1(n9m_reg_64_127_28_31_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[13]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[14]_i_1__4 
       (.I0(n11[14]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[14]_i_2__4_n_0 ),
        .I4(\n1[14]_i_3__4_n_0 ),
        .O(\n9_reg[0] [14]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[14]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_0),
        .O(\n1[14]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[14]_i_3__4 
       (.I0(n11[30]),
        .I1(n9m_reg_64_127_28_31_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[14]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[15]_i_1__4 
       (.I0(n11[15]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[15]_i_2__4_n_0 ),
        .I4(\n1[15]_i_3__4_n_0 ),
        .O(\n9_reg[0] [15]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[15]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_1),
        .O(\n1[15]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[15]_i_3__4 
       (.I0(n11[31]),
        .I1(n9m_reg_64_127_28_31_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[15]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[1]_i_1__4 
       (.I0(n11[1]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[1]_i_2__4_n_0 ),
        .I4(\n1[1]_i_3__4_n_0 ),
        .O(\n9_reg[0] [1]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[1]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_1),
        .O(\n1[1]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[1]_i_3__4 
       (.I0(n11[17]),
        .I1(n9m_reg_64_127_14_20_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[1]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[2]_i_1__4 
       (.I0(n11[2]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[2]_i_2__4_n_0 ),
        .I4(\n1[2]_i_3__4_n_0 ),
        .O(\n9_reg[0] [2]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[2]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_2),
        .O(\n1[2]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[2]_i_3__4 
       (.I0(n11[18]),
        .I1(n9m_reg_64_127_14_20_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[2]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[3]_i_1__4 
       (.I0(n11[3]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[3]_i_2__4_n_0 ),
        .I4(\n1[3]_i_3__4_n_0 ),
        .O(\n9_reg[0] [3]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[3]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_3),
        .O(\n1[3]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[3]_i_3__4 
       (.I0(n11[19]),
        .I1(n9m_reg_64_127_14_20_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[3]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[4]_i_1__4 
       (.I0(n11[4]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[4]_i_2__4_n_0 ),
        .I4(\n1[4]_i_3__4_n_0 ),
        .O(\n9_reg[0] [4]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[4]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_4),
        .O(\n1[4]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[4]_i_3__4 
       (.I0(n11[20]),
        .I1(n9m_reg_64_127_14_20_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[4]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[5]_i_1__4 
       (.I0(n11[5]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[5]_i_2__4_n_0 ),
        .I4(\n1[5]_i_3__4_n_0 ),
        .O(\n9_reg[0] [5]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[5]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_5),
        .O(\n1[5]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[5]_i_3__4 
       (.I0(n11[21]),
        .I1(n9m_reg_64_127_21_27_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[5]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[6]_i_1__4 
       (.I0(n11[6]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[6]_i_2__4_n_0 ),
        .I4(\n1[6]_i_3__4_n_0 ),
        .O(\n9_reg[0] [6]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[6]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_6),
        .O(\n1[6]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[6]_i_3__4 
       (.I0(n11[22]),
        .I1(n9m_reg_64_127_21_27_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[6]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[7]_i_1__4 
       (.I0(n11[7]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[7]_i_2__4_n_0 ),
        .I4(\n1[7]_i_3__4_n_0 ),
        .O(\n9_reg[0] [7]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[7]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_0),
        .O(\n1[7]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[7]_i_3__4 
       (.I0(n11[23]),
        .I1(n9m_reg_64_127_21_27_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[7]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[8]_i_1__4 
       (.I0(n11[8]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[8]_i_2__4_n_0 ),
        .I4(\n1[8]_i_3__4_n_0 ),
        .O(\n9_reg[0] [8]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[8]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_1),
        .O(\n1[8]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[8]_i_3__4 
       (.I0(n11[24]),
        .I1(n9m_reg_64_127_21_27_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[8]_i_3__4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[9]_i_1__4 
       (.I0(n11[9]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[9]_i_2__4_n_0 ),
        .I4(\n1[9]_i_3__4_n_0 ),
        .O(\n9_reg[0] [9]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[9]_i_2__4 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_2),
        .O(\n1[9]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[9]_i_3__4 
       (.I0(n11[25]),
        .I1(n9m_reg_64_127_21_27_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[9]_i_3__4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__11 
       (.I0(n3_reg[0]),
        .O(n2__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__11 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__11 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__11 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__11 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__0[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__11 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__0[5]));
  LUT3 #(
    .INIT(8'hD2)) 
    \n3[6]_i_1__5 
       (.I0(n3_reg[5]),
        .I1(\n3[6]_i_2__5_n_0 ),
        .I2(n3_reg[6]),
        .O(n2__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \n3[6]_i_2__5 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(\n3[6]_i_2__5_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[6]),
        .Q(n3_reg[6]),
        .R(rst_i));
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \n5[0]_i_1__5 
       (.I0(n3_reg[0]),
        .I1(\n5[0]_i_2__5_n_0 ),
        .I2(i8),
        .O(n4));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \n5[0]_i_2__5 
       (.I0(n3_reg[3]),
        .I1(n3_reg[4]),
        .I2(n3_reg[1]),
        .I3(n3_reg[2]),
        .I4(n3_reg[6]),
        .I5(n3_reg[5]),
        .O(\n5[0]_i_2__5_n_0 ));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[6]),
        .Q(n11a[6]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39863 n9m_reg_0_63_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_0_6_n_0),
        .DOB(n9m_reg_0_63_0_6_n_1),
        .DOC(n9m_reg_0_63_0_6_n_2),
        .DOD(n9m_reg_0_63_0_6_n_3),
        .DOE(n9m_reg_0_63_0_6_n_4),
        .DOF(n9m_reg_0_63_0_6_n_5),
        .DOG(n9m_reg_0_63_0_6_n_6),
        .DOH(NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39864 n9m_reg_0_63_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_14_20_n_0),
        .DOB(n9m_reg_0_63_14_20_n_1),
        .DOC(n9m_reg_0_63_14_20_n_2),
        .DOD(n9m_reg_0_63_14_20_n_3),
        .DOE(n9m_reg_0_63_14_20_n_4),
        .DOF(n9m_reg_0_63_14_20_n_5),
        .DOG(n9m_reg_0_63_14_20_n_6),
        .DOH(NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39865 n9m_reg_0_63_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_21_27_n_0),
        .DOB(n9m_reg_0_63_21_27_n_1),
        .DOC(n9m_reg_0_63_21_27_n_2),
        .DOD(n9m_reg_0_63_21_27_n_3),
        .DOE(n9m_reg_0_63_21_27_n_4),
        .DOF(n9m_reg_0_63_21_27_n_5),
        .DOG(n9m_reg_0_63_21_27_n_6),
        .DOH(NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39866 n9m_reg_0_63_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_28_31_n_0),
        .DOB(n9m_reg_0_63_28_31_n_1),
        .DOC(n9m_reg_0_63_28_31_n_2),
        .DOD(n9m_reg_0_63_28_31_n_3),
        .DOE(NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39867 n9m_reg_0_63_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_7_13_n_0),
        .DOB(n9m_reg_0_63_7_13_n_1),
        .DOC(n9m_reg_0_63_7_13_n_2),
        .DOD(n9m_reg_0_63_7_13_n_3),
        .DOE(n9m_reg_0_63_7_13_n_4),
        .DOF(n9m_reg_0_63_7_13_n_5),
        .DOG(n9m_reg_0_63_7_13_n_6),
        .DOH(NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39868 n9m_reg_64_127_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_0_6_n_0),
        .DOB(n9m_reg_64_127_0_6_n_1),
        .DOC(n9m_reg_64_127_0_6_n_2),
        .DOD(n9m_reg_64_127_0_6_n_3),
        .DOE(n9m_reg_64_127_0_6_n_4),
        .DOF(n9m_reg_64_127_0_6_n_5),
        .DOG(n9m_reg_64_127_0_6_n_6),
        .DOH(NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39869 n9m_reg_64_127_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_14_20_n_0),
        .DOB(n9m_reg_64_127_14_20_n_1),
        .DOC(n9m_reg_64_127_14_20_n_2),
        .DOD(n9m_reg_64_127_14_20_n_3),
        .DOE(n9m_reg_64_127_14_20_n_4),
        .DOF(n9m_reg_64_127_14_20_n_5),
        .DOG(n9m_reg_64_127_14_20_n_6),
        .DOH(NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39870 n9m_reg_64_127_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_21_27_n_0),
        .DOB(n9m_reg_64_127_21_27_n_1),
        .DOC(n9m_reg_64_127_21_27_n_2),
        .DOD(n9m_reg_64_127_21_27_n_3),
        .DOE(n9m_reg_64_127_21_27_n_4),
        .DOF(n9m_reg_64_127_21_27_n_5),
        .DOG(n9m_reg_64_127_21_27_n_6),
        .DOH(NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39871 n9m_reg_64_127_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_28_31_n_0),
        .DOB(n9m_reg_64_127_28_31_n_1),
        .DOC(n9m_reg_64_127_28_31_n_2),
        .DOD(n9m_reg_64_127_28_31_n_3),
        .DOE(NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39872 n9m_reg_64_127_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_7_13_n_0),
        .DOB(n9m_reg_64_127_7_13_n_1),
        .DOC(n9m_reg_64_127_7_13_n_2),
        .DOD(n9m_reg_64_127_7_13_n_3),
        .DOE(n9m_reg_64_127_7_13_n_4),
        .DOF(n9m_reg_64_127_7_13_n_5),
        .DOG(n9m_reg_64_127_7_13_n_6),
        .DOH(NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_26" *) 
module switch_elements_cf_fft_512_8_26_21
   (n12,
    p_6_out,
    \n12_reg[0]_0 ,
    n4,
    rst_i,
    enable_i,
    clk_i,
    inf4_s,
    enable_s,
    i8,
    i1);
  output n12;
  output [19:0]p_6_out;
  output [15:0]\n12_reg[0]_0 ;
  output n4;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [7:0]inf4_s;
  input [27:0]enable_s;
  input [0:0]i8;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [27:0]enable_s;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [7:0]inf4_s;
  wire [31:0]n11;
  wire [6:0]n11a;
  wire [5:0]n11a__0;
  wire n12;
  wire [15:0]\n12_reg[0]_0 ;
  wire [6:0]n2__0;
  wire \n3[6]_i_2_n_0 ;
  wire [6:0]n3_reg;
  wire n4;
  wire \n5[0]_i_2_n_0 ;
  wire n6m_reg_0_63_14_20_i_10_n_0;
  wire n6m_reg_0_63_14_20_i_11_n_0;
  wire n6m_reg_0_63_14_20_i_12_n_0;
  wire n6m_reg_0_63_14_20_i_13_n_0;
  wire n6m_reg_0_63_14_20_i_14_n_0;
  wire n6m_reg_0_63_14_20_i_15_n_0;
  wire n6m_reg_0_63_14_20_i_16_n_0;
  wire n6m_reg_0_63_14_20_i_17_n_0;
  wire n6m_reg_0_63_14_20_i_8_n_0;
  wire n6m_reg_0_63_14_20_i_9_n_0;
  wire n6m_reg_0_63_21_27_i_10_n_0;
  wire n6m_reg_0_63_21_27_i_11_n_0;
  wire n6m_reg_0_63_21_27_i_12_n_0;
  wire n6m_reg_0_63_21_27_i_13_n_0;
  wire n6m_reg_0_63_21_27_i_14_n_0;
  wire n6m_reg_0_63_21_27_i_15_n_0;
  wire n6m_reg_0_63_21_27_i_16_n_0;
  wire n6m_reg_0_63_21_27_i_17_n_0;
  wire n6m_reg_0_63_21_27_i_18_n_0;
  wire n6m_reg_0_63_21_27_i_19_n_0;
  wire n6m_reg_0_63_21_27_i_20_n_0;
  wire n6m_reg_0_63_21_27_i_21_n_0;
  wire n6m_reg_0_63_21_27_i_8_n_0;
  wire n6m_reg_0_63_21_27_i_9_n_0;
  wire n6m_reg_0_63_28_31_i_10_n_0;
  wire n6m_reg_0_63_28_31_i_11_n_0;
  wire n6m_reg_0_63_28_31_i_12_n_0;
  wire n6m_reg_0_63_28_31_i_5_n_0;
  wire n6m_reg_0_63_28_31_i_6_n_0;
  wire n6m_reg_0_63_28_31_i_7_n_0;
  wire n6m_reg_0_63_28_31_i_8_n_0;
  wire n6m_reg_0_63_28_31_i_9_n_0;
  wire n9m_reg_0_63_0_6_n_0;
  wire n9m_reg_0_63_0_6_n_1;
  wire n9m_reg_0_63_0_6_n_2;
  wire n9m_reg_0_63_0_6_n_3;
  wire n9m_reg_0_63_0_6_n_4;
  wire n9m_reg_0_63_0_6_n_5;
  wire n9m_reg_0_63_0_6_n_6;
  wire n9m_reg_0_63_14_20_n_0;
  wire n9m_reg_0_63_14_20_n_1;
  wire n9m_reg_0_63_14_20_n_2;
  wire n9m_reg_0_63_14_20_n_3;
  wire n9m_reg_0_63_14_20_n_4;
  wire n9m_reg_0_63_14_20_n_5;
  wire n9m_reg_0_63_14_20_n_6;
  wire n9m_reg_0_63_21_27_n_0;
  wire n9m_reg_0_63_21_27_n_1;
  wire n9m_reg_0_63_21_27_n_2;
  wire n9m_reg_0_63_21_27_n_3;
  wire n9m_reg_0_63_21_27_n_4;
  wire n9m_reg_0_63_21_27_n_5;
  wire n9m_reg_0_63_21_27_n_6;
  wire n9m_reg_0_63_28_31_n_0;
  wire n9m_reg_0_63_28_31_n_1;
  wire n9m_reg_0_63_28_31_n_2;
  wire n9m_reg_0_63_28_31_n_3;
  wire n9m_reg_0_63_7_13_n_0;
  wire n9m_reg_0_63_7_13_n_1;
  wire n9m_reg_0_63_7_13_n_2;
  wire n9m_reg_0_63_7_13_n_3;
  wire n9m_reg_0_63_7_13_n_4;
  wire n9m_reg_0_63_7_13_n_5;
  wire n9m_reg_0_63_7_13_n_6;
  wire n9m_reg_64_127_0_6_n_0;
  wire n9m_reg_64_127_0_6_n_1;
  wire n9m_reg_64_127_0_6_n_2;
  wire n9m_reg_64_127_0_6_n_3;
  wire n9m_reg_64_127_0_6_n_4;
  wire n9m_reg_64_127_0_6_n_5;
  wire n9m_reg_64_127_0_6_n_6;
  wire n9m_reg_64_127_14_20_n_0;
  wire n9m_reg_64_127_14_20_n_1;
  wire n9m_reg_64_127_14_20_n_2;
  wire n9m_reg_64_127_14_20_n_3;
  wire n9m_reg_64_127_14_20_n_4;
  wire n9m_reg_64_127_14_20_n_5;
  wire n9m_reg_64_127_14_20_n_6;
  wire n9m_reg_64_127_21_27_n_0;
  wire n9m_reg_64_127_21_27_n_1;
  wire n9m_reg_64_127_21_27_n_2;
  wire n9m_reg_64_127_21_27_n_3;
  wire n9m_reg_64_127_21_27_n_4;
  wire n9m_reg_64_127_21_27_n_5;
  wire n9m_reg_64_127_21_27_n_6;
  wire n9m_reg_64_127_28_31_n_0;
  wire n9m_reg_64_127_28_31_n_1;
  wire n9m_reg_64_127_28_31_n_2;
  wire n9m_reg_64_127_28_31_n_3;
  wire n9m_reg_64_127_7_13_n_0;
  wire n9m_reg_64_127_7_13_n_1;
  wire n9m_reg_64_127_7_13_n_2;
  wire n9m_reg_64_127_7_13_n_3;
  wire n9m_reg_64_127_7_13_n_4;
  wire n9m_reg_64_127_7_13_n_5;
  wire n9m_reg_64_127_7_13_n_6;
  wire [19:0]p_6_out;
  wire rst_i;
  wire NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED;

  LUT2 #(
    .INIT(4'h6)) 
    \info_o[0]_i_1 
       (.I0(\n12_reg[0]_0 [0]),
        .I1(inf4_s[0]),
        .O(p_6_out[0]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[10]_i_1 
       (.I0(\n12_reg[0]_0 [10]),
        .I1(enable_s[6]),
        .I2(enable_s[22]),
        .O(p_6_out[10]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[11]_i_1 
       (.I0(\n12_reg[0]_0 [11]),
        .I1(enable_s[7]),
        .I2(enable_s[23]),
        .O(p_6_out[11]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[12]_i_1 
       (.I0(\n12_reg[0]_0 [12]),
        .I1(enable_s[8]),
        .I2(enable_s[24]),
        .O(p_6_out[12]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[13]_i_1 
       (.I0(\n12_reg[0]_0 [13]),
        .I1(enable_s[9]),
        .I2(enable_s[25]),
        .O(p_6_out[13]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[14]_i_1 
       (.I0(\n12_reg[0]_0 [14]),
        .I1(enable_s[10]),
        .I2(enable_s[26]),
        .O(p_6_out[14]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[15]_i_1 
       (.I0(\n12_reg[0]_0 [15]),
        .I1(enable_s[11]),
        .I2(enable_s[27]),
        .O(p_6_out[15]));
  LUT2 #(
    .INIT(4'h6)) 
    \info_o[1]_i_1 
       (.I0(\n12_reg[0]_0 [1]),
        .I1(inf4_s[1]),
        .O(p_6_out[1]));
  LUT5 #(
    .INIT(32'h69969669)) 
    \info_o[28]_i_1 
       (.I0(inf4_s[4]),
        .I1(enable_s[12]),
        .I2(\n12_reg[0]_0 [12]),
        .I3(enable_s[8]),
        .I4(\n12_reg[0]_0 [8]),
        .O(p_6_out[16]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \info_o[29]_i_1 
       (.I0(inf4_s[5]),
        .I1(enable_s[13]),
        .I2(\n12_reg[0]_0 [13]),
        .I3(enable_s[9]),
        .I4(\n12_reg[0]_0 [9]),
        .O(p_6_out[17]));
  LUT2 #(
    .INIT(4'h6)) 
    \info_o[2]_i_1 
       (.I0(\n12_reg[0]_0 [2]),
        .I1(inf4_s[2]),
        .O(p_6_out[2]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \info_o[30]_i_1 
       (.I0(inf4_s[6]),
        .I1(enable_s[14]),
        .I2(\n12_reg[0]_0 [14]),
        .I3(enable_s[10]),
        .I4(\n12_reg[0]_0 [10]),
        .O(p_6_out[18]));
  LUT5 #(
    .INIT(32'h96696996)) 
    \info_o[31]_i_1 
       (.I0(inf4_s[7]),
        .I1(enable_s[15]),
        .I2(\n12_reg[0]_0 [15]),
        .I3(enable_s[11]),
        .I4(\n12_reg[0]_0 [11]),
        .O(p_6_out[19]));
  LUT2 #(
    .INIT(4'h6)) 
    \info_o[3]_i_1 
       (.I0(\n12_reg[0]_0 [3]),
        .I1(inf4_s[3]),
        .O(p_6_out[3]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[4]_i_1 
       (.I0(\n12_reg[0]_0 [4]),
        .I1(enable_s[0]),
        .I2(enable_s[16]),
        .O(p_6_out[4]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[5]_i_1 
       (.I0(\n12_reg[0]_0 [5]),
        .I1(enable_s[1]),
        .I2(enable_s[17]),
        .O(p_6_out[5]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[6]_i_1 
       (.I0(\n12_reg[0]_0 [6]),
        .I1(enable_s[2]),
        .I2(enable_s[18]),
        .O(p_6_out[6]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[7]_i_1 
       (.I0(\n12_reg[0]_0 [7]),
        .I1(enable_s[3]),
        .I2(enable_s[19]),
        .O(p_6_out[7]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[8]_i_1 
       (.I0(\n12_reg[0]_0 [8]),
        .I1(enable_s[4]),
        .I2(enable_s[20]),
        .O(p_6_out[8]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[9]_i_1 
       (.I0(\n12_reg[0]_0 [9]),
        .I1(enable_s[5]),
        .I2(enable_s[21]),
        .O(p_6_out[9]));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39718 n11m_reg_0_63_0_6
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[14]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n11[0]),
        .DOB(n11[1]),
        .DOC(n11[2]),
        .DOD(n11[3]),
        .DOE(n11[4]),
        .DOF(n11[5]),
        .DOG(n11[6]),
        .DOH(NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39719 n11m_reg_0_63_14_20
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[12]),
        .DIB(i1[13]),
        .DIC(i1[14]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n11[14]),
        .DOB(n11[15]),
        .DOC(n11[16]),
        .DOD(n11[17]),
        .DOE(n11[18]),
        .DOF(n11[19]),
        .DOG(n11[20]),
        .DOH(NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39720 n11m_reg_0_63_21_27
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n11[21]),
        .DOB(n11[22]),
        .DOC(n11[23]),
        .DOD(n11[24]),
        .DOE(n11[25]),
        .DOF(n11[26]),
        .DOG(n11[27]),
        .DOH(NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39721 n11m_reg_0_63_28_31
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n11[28]),
        .DOB(n11[29]),
        .DOC(n11[30]),
        .DOD(n11[31]),
        .DOE(NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39722 n11m_reg_0_63_7_13
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[22]),
        .DIC(i1[7]),
        .DID(i1[8]),
        .DIE(i1[9]),
        .DIF(i1[10]),
        .DIG(i1[11]),
        .DIH(1'b0),
        .DOA(n11[7]),
        .DOB(n11[8]),
        .DOC(n11[9]),
        .DOD(n11[10]),
        .DOE(n11[11]),
        .DOF(n11[12]),
        .DOG(n11[13]),
        .DOH(NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n12_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(1'b1),
        .Q(n12),
        .R(rst_i));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1 
       (.I0(n3_reg[0]),
        .O(n2__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__0[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__0[5]));
  LUT3 #(
    .INIT(8'hD2)) 
    \n3[6]_i_1 
       (.I0(n3_reg[5]),
        .I1(\n3[6]_i_2_n_0 ),
        .I2(n3_reg[6]),
        .O(n2__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \n3[6]_i_2 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(\n3[6]_i_2_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[6]),
        .Q(n3_reg[6]),
        .R(rst_i));
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \n5[0]_i_1 
       (.I0(n3_reg[0]),
        .I1(\n5[0]_i_2_n_0 ),
        .I2(i8),
        .O(n4));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \n5[0]_i_2 
       (.I0(n3_reg[3]),
        .I1(n3_reg[4]),
        .I2(n3_reg[1]),
        .I3(n3_reg[2]),
        .I4(n3_reg[6]),
        .I5(n3_reg[5]),
        .O(\n5[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_14_20_i_10
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_1),
        .O(n6m_reg_0_63_14_20_i_10_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_14_20_i_11
       (.I0(n11[17]),
        .I1(n9m_reg_64_127_14_20_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_3),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_14_20_i_11_n_0));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_14_20_i_12
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_2),
        .O(n6m_reg_0_63_14_20_i_12_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_14_20_i_13
       (.I0(n11[18]),
        .I1(n9m_reg_64_127_14_20_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_4),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_14_20_i_13_n_0));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_14_20_i_14
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_3),
        .O(n6m_reg_0_63_14_20_i_14_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_14_20_i_15
       (.I0(n11[19]),
        .I1(n9m_reg_64_127_14_20_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_5),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_14_20_i_15_n_0));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_14_20_i_16
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_4),
        .O(n6m_reg_0_63_14_20_i_16_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_14_20_i_17
       (.I0(n11[20]),
        .I1(n9m_reg_64_127_14_20_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_6),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_14_20_i_17_n_0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_14_20_i_3
       (.I0(n11[0]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_i_8_n_0),
        .I4(n6m_reg_0_63_14_20_i_9_n_0),
        .O(\n12_reg[0]_0 [0]));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_14_20_i_4
       (.I0(n11[1]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_i_10_n_0),
        .I4(n6m_reg_0_63_14_20_i_11_n_0),
        .O(\n12_reg[0]_0 [1]));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_14_20_i_5
       (.I0(n11[2]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_i_12_n_0),
        .I4(n6m_reg_0_63_14_20_i_13_n_0),
        .O(\n12_reg[0]_0 [2]));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_14_20_i_6
       (.I0(n11[3]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_i_14_n_0),
        .I4(n6m_reg_0_63_14_20_i_15_n_0),
        .O(\n12_reg[0]_0 [3]));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_14_20_i_7
       (.I0(n11[4]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_i_16_n_0),
        .I4(n6m_reg_0_63_14_20_i_17_n_0),
        .O(\n12_reg[0]_0 [4]));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_14_20_i_8
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_0),
        .O(n6m_reg_0_63_14_20_i_8_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_14_20_i_9
       (.I0(n11[16]),
        .I1(n9m_reg_64_127_14_20_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_2),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_14_20_i_9_n_0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_21_27_i_1
       (.I0(n11[5]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_21_27_i_8_n_0),
        .I4(n6m_reg_0_63_21_27_i_9_n_0),
        .O(\n12_reg[0]_0 [5]));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_21_27_i_10
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_6),
        .O(n6m_reg_0_63_21_27_i_10_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_21_27_i_11
       (.I0(n11[22]),
        .I1(n9m_reg_64_127_21_27_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_1),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_21_27_i_11_n_0));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_21_27_i_12
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_0),
        .O(n6m_reg_0_63_21_27_i_12_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_21_27_i_13
       (.I0(n11[23]),
        .I1(n9m_reg_64_127_21_27_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_2),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_21_27_i_13_n_0));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_21_27_i_14
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_1),
        .O(n6m_reg_0_63_21_27_i_14_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_21_27_i_15
       (.I0(n11[24]),
        .I1(n9m_reg_64_127_21_27_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_3),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_21_27_i_15_n_0));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_21_27_i_16
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_2),
        .O(n6m_reg_0_63_21_27_i_16_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_21_27_i_17
       (.I0(n11[25]),
        .I1(n9m_reg_64_127_21_27_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_4),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_21_27_i_17_n_0));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_21_27_i_18
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_3),
        .O(n6m_reg_0_63_21_27_i_18_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_21_27_i_19
       (.I0(n11[26]),
        .I1(n9m_reg_64_127_21_27_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_5),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_21_27_i_19_n_0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_21_27_i_2
       (.I0(n11[6]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_21_27_i_10_n_0),
        .I4(n6m_reg_0_63_21_27_i_11_n_0),
        .O(\n12_reg[0]_0 [6]));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_21_27_i_20
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_4),
        .O(n6m_reg_0_63_21_27_i_20_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_21_27_i_21
       (.I0(n11[27]),
        .I1(n9m_reg_64_127_21_27_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_6),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_21_27_i_21_n_0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_21_27_i_3
       (.I0(n11[7]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_21_27_i_12_n_0),
        .I4(n6m_reg_0_63_21_27_i_13_n_0),
        .O(\n12_reg[0]_0 [7]));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_21_27_i_4
       (.I0(n11[8]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_21_27_i_14_n_0),
        .I4(n6m_reg_0_63_21_27_i_15_n_0),
        .O(\n12_reg[0]_0 [8]));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_21_27_i_5
       (.I0(n11[9]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_21_27_i_16_n_0),
        .I4(n6m_reg_0_63_21_27_i_17_n_0),
        .O(\n12_reg[0]_0 [9]));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_21_27_i_6
       (.I0(n11[10]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_21_27_i_18_n_0),
        .I4(n6m_reg_0_63_21_27_i_19_n_0),
        .O(\n12_reg[0]_0 [10]));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_21_27_i_7
       (.I0(n11[11]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_21_27_i_20_n_0),
        .I4(n6m_reg_0_63_21_27_i_21_n_0),
        .O(\n12_reg[0]_0 [11]));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_21_27_i_8
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_5),
        .O(n6m_reg_0_63_21_27_i_8_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_21_27_i_9
       (.I0(n11[21]),
        .I1(n9m_reg_64_127_21_27_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_0),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_21_27_i_9_n_0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_28_31_i_1
       (.I0(n11[12]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_28_31_i_5_n_0),
        .I4(n6m_reg_0_63_28_31_i_6_n_0),
        .O(\n12_reg[0]_0 [12]));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_28_31_i_10
       (.I0(n11[30]),
        .I1(n9m_reg_64_127_28_31_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_2),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_28_31_i_10_n_0));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_28_31_i_11
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_1),
        .O(n6m_reg_0_63_28_31_i_11_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_28_31_i_12
       (.I0(n11[31]),
        .I1(n9m_reg_64_127_28_31_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_3),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_28_31_i_12_n_0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_28_31_i_2
       (.I0(n11[13]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_28_31_i_7_n_0),
        .I4(n6m_reg_0_63_28_31_i_8_n_0),
        .O(\n12_reg[0]_0 [13]));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_28_31_i_3
       (.I0(n11[14]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_28_31_i_9_n_0),
        .I4(n6m_reg_0_63_28_31_i_10_n_0),
        .O(\n12_reg[0]_0 [14]));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    n6m_reg_0_63_28_31_i_4
       (.I0(n11[15]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_28_31_i_11_n_0),
        .I4(n6m_reg_0_63_28_31_i_12_n_0),
        .O(\n12_reg[0]_0 [15]));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_28_31_i_5
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_5),
        .O(n6m_reg_0_63_28_31_i_5_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_28_31_i_6
       (.I0(n11[28]),
        .I1(n9m_reg_64_127_28_31_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_0),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_28_31_i_6_n_0));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_28_31_i_7
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_6),
        .O(n6m_reg_0_63_28_31_i_7_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    n6m_reg_0_63_28_31_i_8
       (.I0(n11[29]),
        .I1(n9m_reg_64_127_28_31_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_1),
        .I4(n12),
        .I5(i8),
        .O(n6m_reg_0_63_28_31_i_8_n_0));
  LUT5 #(
    .INIT(32'h44400040)) 
    n6m_reg_0_63_28_31_i_9
       (.I0(n12),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_0),
        .O(n6m_reg_0_63_28_31_i_9_n_0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[6]),
        .Q(n11a[6]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39723 n9m_reg_0_63_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[14]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_0_6_n_0),
        .DOB(n9m_reg_0_63_0_6_n_1),
        .DOC(n9m_reg_0_63_0_6_n_2),
        .DOD(n9m_reg_0_63_0_6_n_3),
        .DOE(n9m_reg_0_63_0_6_n_4),
        .DOF(n9m_reg_0_63_0_6_n_5),
        .DOG(n9m_reg_0_63_0_6_n_6),
        .DOH(NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39724 n9m_reg_0_63_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[12]),
        .DIB(i1[13]),
        .DIC(i1[14]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_14_20_n_0),
        .DOB(n9m_reg_0_63_14_20_n_1),
        .DOC(n9m_reg_0_63_14_20_n_2),
        .DOD(n9m_reg_0_63_14_20_n_3),
        .DOE(n9m_reg_0_63_14_20_n_4),
        .DOF(n9m_reg_0_63_14_20_n_5),
        .DOG(n9m_reg_0_63_14_20_n_6),
        .DOH(NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39725 n9m_reg_0_63_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_21_27_n_0),
        .DOB(n9m_reg_0_63_21_27_n_1),
        .DOC(n9m_reg_0_63_21_27_n_2),
        .DOD(n9m_reg_0_63_21_27_n_3),
        .DOE(n9m_reg_0_63_21_27_n_4),
        .DOF(n9m_reg_0_63_21_27_n_5),
        .DOG(n9m_reg_0_63_21_27_n_6),
        .DOH(NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39726 n9m_reg_0_63_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_28_31_n_0),
        .DOB(n9m_reg_0_63_28_31_n_1),
        .DOC(n9m_reg_0_63_28_31_n_2),
        .DOD(n9m_reg_0_63_28_31_n_3),
        .DOE(NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39727 n9m_reg_0_63_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[22]),
        .DIC(i1[7]),
        .DID(i1[8]),
        .DIE(i1[9]),
        .DIF(i1[10]),
        .DIG(i1[11]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_7_13_n_0),
        .DOB(n9m_reg_0_63_7_13_n_1),
        .DOC(n9m_reg_0_63_7_13_n_2),
        .DOD(n9m_reg_0_63_7_13_n_3),
        .DOE(n9m_reg_0_63_7_13_n_4),
        .DOF(n9m_reg_0_63_7_13_n_5),
        .DOG(n9m_reg_0_63_7_13_n_6),
        .DOH(NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39728 n9m_reg_64_127_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[14]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_0_6_n_0),
        .DOB(n9m_reg_64_127_0_6_n_1),
        .DOC(n9m_reg_64_127_0_6_n_2),
        .DOD(n9m_reg_64_127_0_6_n_3),
        .DOE(n9m_reg_64_127_0_6_n_4),
        .DOF(n9m_reg_64_127_0_6_n_5),
        .DOG(n9m_reg_64_127_0_6_n_6),
        .DOH(NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39729 n9m_reg_64_127_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[12]),
        .DIB(i1[13]),
        .DIC(i1[14]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_14_20_n_0),
        .DOB(n9m_reg_64_127_14_20_n_1),
        .DOC(n9m_reg_64_127_14_20_n_2),
        .DOD(n9m_reg_64_127_14_20_n_3),
        .DOE(n9m_reg_64_127_14_20_n_4),
        .DOF(n9m_reg_64_127_14_20_n_5),
        .DOG(n9m_reg_64_127_14_20_n_6),
        .DOH(NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39730 n9m_reg_64_127_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_21_27_n_0),
        .DOB(n9m_reg_64_127_21_27_n_1),
        .DOC(n9m_reg_64_127_21_27_n_2),
        .DOD(n9m_reg_64_127_21_27_n_3),
        .DOE(n9m_reg_64_127_21_27_n_4),
        .DOF(n9m_reg_64_127_21_27_n_5),
        .DOG(n9m_reg_64_127_21_27_n_6),
        .DOH(NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39731 n9m_reg_64_127_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_28_31_n_0),
        .DOB(n9m_reg_64_127_28_31_n_1),
        .DOC(n9m_reg_64_127_28_31_n_2),
        .DOD(n9m_reg_64_127_28_31_n_3),
        .DOE(NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39732 n9m_reg_64_127_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[22]),
        .DIC(i1[7]),
        .DID(i1[8]),
        .DIE(i1[9]),
        .DIF(i1[10]),
        .DIG(i1[11]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_7_13_n_0),
        .DOB(n9m_reg_64_127_7_13_n_1),
        .DOC(n9m_reg_64_127_7_13_n_2),
        .DOD(n9m_reg_64_127_7_13_n_3),
        .DOE(n9m_reg_64_127_7_13_n_4),
        .DOF(n9m_reg_64_127_7_13_n_5),
        .DOG(n9m_reg_64_127_7_13_n_6),
        .DOH(NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_26" *) 
module switch_elements_cf_fft_512_8_26_25
   (D,
    n4,
    \n1_reg[15] ,
    i8,
    rst_i,
    enable_i,
    clk_i,
    i1);
  output [15:0]D;
  output n4;
  input \n1_reg[15] ;
  input [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [29:0]i1;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [6:0]n11a;
  wire [5:0]n11a__0;
  wire n11m_reg_0_63_0_6_n_0;
  wire n11m_reg_0_63_0_6_n_1;
  wire n11m_reg_0_63_0_6_n_2;
  wire n11m_reg_0_63_0_6_n_3;
  wire n11m_reg_0_63_0_6_n_4;
  wire n11m_reg_0_63_0_6_n_5;
  wire n11m_reg_0_63_0_6_n_6;
  wire n11m_reg_0_63_14_20_n_0;
  wire n11m_reg_0_63_14_20_n_1;
  wire n11m_reg_0_63_14_20_n_2;
  wire n11m_reg_0_63_14_20_n_3;
  wire n11m_reg_0_63_14_20_n_4;
  wire n11m_reg_0_63_14_20_n_5;
  wire n11m_reg_0_63_14_20_n_6;
  wire n11m_reg_0_63_21_27_n_0;
  wire n11m_reg_0_63_21_27_n_1;
  wire n11m_reg_0_63_21_27_n_2;
  wire n11m_reg_0_63_21_27_n_3;
  wire n11m_reg_0_63_21_27_n_4;
  wire n11m_reg_0_63_21_27_n_5;
  wire n11m_reg_0_63_21_27_n_6;
  wire n11m_reg_0_63_28_31_n_0;
  wire n11m_reg_0_63_28_31_n_1;
  wire n11m_reg_0_63_28_31_n_2;
  wire n11m_reg_0_63_28_31_n_3;
  wire n11m_reg_0_63_7_13_n_0;
  wire n11m_reg_0_63_7_13_n_1;
  wire n11m_reg_0_63_7_13_n_2;
  wire n11m_reg_0_63_7_13_n_3;
  wire n11m_reg_0_63_7_13_n_4;
  wire n11m_reg_0_63_7_13_n_5;
  wire n11m_reg_0_63_7_13_n_6;
  wire \n1[0]_i_2__7_n_0 ;
  wire \n1[0]_i_3__7_n_0 ;
  wire \n1[10]_i_2__7_n_0 ;
  wire \n1[10]_i_3__7_n_0 ;
  wire \n1[11]_i_2__7_n_0 ;
  wire \n1[11]_i_3__7_n_0 ;
  wire \n1[12]_i_2__7_n_0 ;
  wire \n1[12]_i_3__7_n_0 ;
  wire \n1[13]_i_2__7_n_0 ;
  wire \n1[13]_i_3__7_n_0 ;
  wire \n1[14]_i_2__7_n_0 ;
  wire \n1[14]_i_3__7_n_0 ;
  wire \n1[15]_i_2__7_n_0 ;
  wire \n1[15]_i_3__7_n_0 ;
  wire \n1[1]_i_2__7_n_0 ;
  wire \n1[1]_i_3__7_n_0 ;
  wire \n1[2]_i_2__7_n_0 ;
  wire \n1[2]_i_3__7_n_0 ;
  wire \n1[3]_i_2__7_n_0 ;
  wire \n1[3]_i_3__7_n_0 ;
  wire \n1[4]_i_2__7_n_0 ;
  wire \n1[4]_i_3__7_n_0 ;
  wire \n1[5]_i_2__7_n_0 ;
  wire \n1[5]_i_3__7_n_0 ;
  wire \n1[6]_i_2__7_n_0 ;
  wire \n1[6]_i_3__7_n_0 ;
  wire \n1[7]_i_2__7_n_0 ;
  wire \n1[7]_i_3__7_n_0 ;
  wire \n1[8]_i_2__7_n_0 ;
  wire \n1[8]_i_3__7_n_0 ;
  wire \n1[9]_i_2__7_n_0 ;
  wire \n1[9]_i_3__7_n_0 ;
  wire \n1_reg[15] ;
  wire [6:0]n2;
  wire \n3[6]_i_2__7_n_0 ;
  wire [6:0]n3_reg;
  wire n4;
  wire \n5[0]_i_2__7_n_0 ;
  wire n9m_reg_0_63_0_6_n_0;
  wire n9m_reg_0_63_0_6_n_1;
  wire n9m_reg_0_63_0_6_n_2;
  wire n9m_reg_0_63_0_6_n_3;
  wire n9m_reg_0_63_0_6_n_4;
  wire n9m_reg_0_63_0_6_n_5;
  wire n9m_reg_0_63_0_6_n_6;
  wire n9m_reg_0_63_14_20_n_0;
  wire n9m_reg_0_63_14_20_n_1;
  wire n9m_reg_0_63_14_20_n_2;
  wire n9m_reg_0_63_14_20_n_3;
  wire n9m_reg_0_63_14_20_n_4;
  wire n9m_reg_0_63_14_20_n_5;
  wire n9m_reg_0_63_14_20_n_6;
  wire n9m_reg_0_63_21_27_n_0;
  wire n9m_reg_0_63_21_27_n_1;
  wire n9m_reg_0_63_21_27_n_2;
  wire n9m_reg_0_63_21_27_n_3;
  wire n9m_reg_0_63_21_27_n_4;
  wire n9m_reg_0_63_21_27_n_5;
  wire n9m_reg_0_63_21_27_n_6;
  wire n9m_reg_0_63_28_31_n_0;
  wire n9m_reg_0_63_28_31_n_1;
  wire n9m_reg_0_63_28_31_n_2;
  wire n9m_reg_0_63_28_31_n_3;
  wire n9m_reg_0_63_7_13_n_0;
  wire n9m_reg_0_63_7_13_n_1;
  wire n9m_reg_0_63_7_13_n_2;
  wire n9m_reg_0_63_7_13_n_3;
  wire n9m_reg_0_63_7_13_n_4;
  wire n9m_reg_0_63_7_13_n_5;
  wire n9m_reg_0_63_7_13_n_6;
  wire n9m_reg_64_127_0_6_n_0;
  wire n9m_reg_64_127_0_6_n_1;
  wire n9m_reg_64_127_0_6_n_2;
  wire n9m_reg_64_127_0_6_n_3;
  wire n9m_reg_64_127_0_6_n_4;
  wire n9m_reg_64_127_0_6_n_5;
  wire n9m_reg_64_127_0_6_n_6;
  wire n9m_reg_64_127_14_20_n_0;
  wire n9m_reg_64_127_14_20_n_1;
  wire n9m_reg_64_127_14_20_n_2;
  wire n9m_reg_64_127_14_20_n_3;
  wire n9m_reg_64_127_14_20_n_4;
  wire n9m_reg_64_127_14_20_n_5;
  wire n9m_reg_64_127_14_20_n_6;
  wire n9m_reg_64_127_21_27_n_0;
  wire n9m_reg_64_127_21_27_n_1;
  wire n9m_reg_64_127_21_27_n_2;
  wire n9m_reg_64_127_21_27_n_3;
  wire n9m_reg_64_127_21_27_n_4;
  wire n9m_reg_64_127_21_27_n_5;
  wire n9m_reg_64_127_21_27_n_6;
  wire n9m_reg_64_127_28_31_n_0;
  wire n9m_reg_64_127_28_31_n_1;
  wire n9m_reg_64_127_28_31_n_2;
  wire n9m_reg_64_127_28_31_n_3;
  wire n9m_reg_64_127_7_13_n_0;
  wire n9m_reg_64_127_7_13_n_1;
  wire n9m_reg_64_127_7_13_n_2;
  wire n9m_reg_64_127_7_13_n_3;
  wire n9m_reg_64_127_7_13_n_4;
  wire n9m_reg_64_127_7_13_n_5;
  wire n9m_reg_64_127_7_13_n_6;
  wire rst_i;
  wire NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED;

  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39693 n11m_reg_0_63_0_6
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[14]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_0_6_n_0),
        .DOB(n11m_reg_0_63_0_6_n_1),
        .DOC(n11m_reg_0_63_0_6_n_2),
        .DOD(n11m_reg_0_63_0_6_n_3),
        .DOE(n11m_reg_0_63_0_6_n_4),
        .DOF(n11m_reg_0_63_0_6_n_5),
        .DOG(n11m_reg_0_63_0_6_n_6),
        .DOH(NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39694 n11m_reg_0_63_14_20
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[12]),
        .DIB(i1[13]),
        .DIC(i1[14]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_14_20_n_0),
        .DOB(n11m_reg_0_63_14_20_n_1),
        .DOC(n11m_reg_0_63_14_20_n_2),
        .DOD(n11m_reg_0_63_14_20_n_3),
        .DOE(n11m_reg_0_63_14_20_n_4),
        .DOF(n11m_reg_0_63_14_20_n_5),
        .DOG(n11m_reg_0_63_14_20_n_6),
        .DOH(NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39695 n11m_reg_0_63_21_27
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_21_27_n_0),
        .DOB(n11m_reg_0_63_21_27_n_1),
        .DOC(n11m_reg_0_63_21_27_n_2),
        .DOD(n11m_reg_0_63_21_27_n_3),
        .DOE(n11m_reg_0_63_21_27_n_4),
        .DOF(n11m_reg_0_63_21_27_n_5),
        .DOG(n11m_reg_0_63_21_27_n_6),
        .DOH(NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39696 n11m_reg_0_63_28_31
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_28_31_n_0),
        .DOB(n11m_reg_0_63_28_31_n_1),
        .DOC(n11m_reg_0_63_28_31_n_2),
        .DOD(n11m_reg_0_63_28_31_n_3),
        .DOE(NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39697 n11m_reg_0_63_7_13
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[22]),
        .DIC(i1[7]),
        .DID(i1[8]),
        .DIE(i1[9]),
        .DIF(i1[10]),
        .DIG(i1[11]),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_7_13_n_0),
        .DOB(n11m_reg_0_63_7_13_n_1),
        .DOC(n11m_reg_0_63_7_13_n_2),
        .DOD(n11m_reg_0_63_7_13_n_3),
        .DOE(n11m_reg_0_63_7_13_n_4),
        .DOF(n11m_reg_0_63_7_13_n_5),
        .DOG(n11m_reg_0_63_7_13_n_6),
        .DOH(NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[0]_i_1__6 
       (.I0(n11m_reg_0_63_0_6_n_0),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[0]_i_2__7_n_0 ),
        .I4(\n1[0]_i_3__7_n_0 ),
        .O(D[0]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[0]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_0),
        .O(\n1[0]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[0]_i_3__7 
       (.I0(n11m_reg_0_63_14_20_n_2),
        .I1(n9m_reg_64_127_14_20_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_2),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[0]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[10]_i_1__6 
       (.I0(n11m_reg_0_63_7_13_n_3),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[10]_i_2__7_n_0 ),
        .I4(\n1[10]_i_3__7_n_0 ),
        .O(D[10]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[10]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_3),
        .O(\n1[10]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[10]_i_3__7 
       (.I0(n11m_reg_0_63_21_27_n_5),
        .I1(n9m_reg_64_127_21_27_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_5),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[10]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[11]_i_1__6 
       (.I0(n11m_reg_0_63_7_13_n_4),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[11]_i_2__7_n_0 ),
        .I4(\n1[11]_i_3__7_n_0 ),
        .O(D[11]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[11]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_4),
        .O(\n1[11]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[11]_i_3__7 
       (.I0(n11m_reg_0_63_21_27_n_6),
        .I1(n9m_reg_64_127_21_27_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_6),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[11]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[12]_i_1__6 
       (.I0(n11m_reg_0_63_7_13_n_5),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[12]_i_2__7_n_0 ),
        .I4(\n1[12]_i_3__7_n_0 ),
        .O(D[12]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[12]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_5),
        .O(\n1[12]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[12]_i_3__7 
       (.I0(n11m_reg_0_63_28_31_n_0),
        .I1(n9m_reg_64_127_28_31_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_0),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[12]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[13]_i_1__6 
       (.I0(n11m_reg_0_63_7_13_n_6),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[13]_i_2__7_n_0 ),
        .I4(\n1[13]_i_3__7_n_0 ),
        .O(D[13]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[13]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_6),
        .O(\n1[13]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[13]_i_3__7 
       (.I0(n11m_reg_0_63_28_31_n_1),
        .I1(n9m_reg_64_127_28_31_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_1),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[13]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[14]_i_1__6 
       (.I0(n11m_reg_0_63_14_20_n_0),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[14]_i_2__7_n_0 ),
        .I4(\n1[14]_i_3__7_n_0 ),
        .O(D[14]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[14]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_0),
        .O(\n1[14]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[14]_i_3__7 
       (.I0(n11m_reg_0_63_28_31_n_2),
        .I1(n9m_reg_64_127_28_31_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_2),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[14]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[15]_i_1__6 
       (.I0(n11m_reg_0_63_14_20_n_1),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[15]_i_2__7_n_0 ),
        .I4(\n1[15]_i_3__7_n_0 ),
        .O(D[15]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[15]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_1),
        .O(\n1[15]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[15]_i_3__7 
       (.I0(n11m_reg_0_63_28_31_n_3),
        .I1(n9m_reg_64_127_28_31_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_3),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[15]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[1]_i_1__6 
       (.I0(n11m_reg_0_63_0_6_n_1),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[1]_i_2__7_n_0 ),
        .I4(\n1[1]_i_3__7_n_0 ),
        .O(D[1]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[1]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_1),
        .O(\n1[1]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[1]_i_3__7 
       (.I0(n11m_reg_0_63_14_20_n_3),
        .I1(n9m_reg_64_127_14_20_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_3),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[1]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[2]_i_1__6 
       (.I0(n11m_reg_0_63_0_6_n_2),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[2]_i_2__7_n_0 ),
        .I4(\n1[2]_i_3__7_n_0 ),
        .O(D[2]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[2]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_2),
        .O(\n1[2]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[2]_i_3__7 
       (.I0(n11m_reg_0_63_14_20_n_4),
        .I1(n9m_reg_64_127_14_20_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_4),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[2]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[3]_i_1__6 
       (.I0(n11m_reg_0_63_0_6_n_3),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[3]_i_2__7_n_0 ),
        .I4(\n1[3]_i_3__7_n_0 ),
        .O(D[3]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[3]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_3),
        .O(\n1[3]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[3]_i_3__7 
       (.I0(n11m_reg_0_63_14_20_n_5),
        .I1(n9m_reg_64_127_14_20_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_5),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[3]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[4]_i_1__6 
       (.I0(n11m_reg_0_63_0_6_n_4),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[4]_i_2__7_n_0 ),
        .I4(\n1[4]_i_3__7_n_0 ),
        .O(D[4]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[4]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_4),
        .O(\n1[4]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[4]_i_3__7 
       (.I0(n11m_reg_0_63_14_20_n_6),
        .I1(n9m_reg_64_127_14_20_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_6),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[4]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[5]_i_1__6 
       (.I0(n11m_reg_0_63_0_6_n_5),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[5]_i_2__7_n_0 ),
        .I4(\n1[5]_i_3__7_n_0 ),
        .O(D[5]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[5]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_5),
        .O(\n1[5]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[5]_i_3__7 
       (.I0(n11m_reg_0_63_21_27_n_0),
        .I1(n9m_reg_64_127_21_27_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_0),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[5]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[6]_i_1__6 
       (.I0(n11m_reg_0_63_0_6_n_6),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[6]_i_2__7_n_0 ),
        .I4(\n1[6]_i_3__7_n_0 ),
        .O(D[6]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[6]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_6),
        .O(\n1[6]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[6]_i_3__7 
       (.I0(n11m_reg_0_63_21_27_n_1),
        .I1(n9m_reg_64_127_21_27_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_1),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[6]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[7]_i_1__6 
       (.I0(n11m_reg_0_63_7_13_n_0),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[7]_i_2__7_n_0 ),
        .I4(\n1[7]_i_3__7_n_0 ),
        .O(D[7]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[7]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_0),
        .O(\n1[7]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[7]_i_3__7 
       (.I0(n11m_reg_0_63_21_27_n_2),
        .I1(n9m_reg_64_127_21_27_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_2),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[7]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[8]_i_1__6 
       (.I0(n11m_reg_0_63_7_13_n_1),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[8]_i_2__7_n_0 ),
        .I4(\n1[8]_i_3__7_n_0 ),
        .O(D[8]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[8]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_1),
        .O(\n1[8]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[8]_i_3__7 
       (.I0(n11m_reg_0_63_21_27_n_3),
        .I1(n9m_reg_64_127_21_27_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_3),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[8]_i_3__7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[9]_i_1__6 
       (.I0(n11m_reg_0_63_7_13_n_2),
        .I1(\n1_reg[15] ),
        .I2(i8),
        .I3(\n1[9]_i_2__7_n_0 ),
        .I4(\n1[9]_i_3__7_n_0 ),
        .O(D[9]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[9]_i_2__7 
       (.I0(\n1_reg[15] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_2),
        .O(\n1[9]_i_2__7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[9]_i_3__7 
       (.I0(n11m_reg_0_63_21_27_n_4),
        .I1(n9m_reg_64_127_21_27_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_4),
        .I4(\n1_reg[15] ),
        .I5(i8),
        .O(\n1[9]_i_3__7_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__15 
       (.I0(n3_reg[0]),
        .O(n2[0]));
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__15 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2[1]));
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__15 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2[2]));
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__15 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2[3]));
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__15 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__15 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2[5]));
  LUT3 #(
    .INIT(8'hD2)) 
    \n3[6]_i_1__7 
       (.I0(n3_reg[5]),
        .I1(\n3[6]_i_2__7_n_0 ),
        .I2(n3_reg[6]),
        .O(n2[6]));
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \n3[6]_i_2__7 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(\n3[6]_i_2__7_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[6]),
        .Q(n3_reg[6]),
        .R(rst_i));
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \n5[0]_i_1__7 
       (.I0(n3_reg[0]),
        .I1(\n5[0]_i_2__7_n_0 ),
        .I2(i8),
        .O(n4));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \n5[0]_i_2__7 
       (.I0(n3_reg[3]),
        .I1(n3_reg[4]),
        .I2(n3_reg[1]),
        .I3(n3_reg[2]),
        .I4(n3_reg[6]),
        .I5(n3_reg[5]),
        .O(\n5[0]_i_2__7_n_0 ));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[6]),
        .Q(n11a[6]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39698 n9m_reg_0_63_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[14]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_0_6_n_0),
        .DOB(n9m_reg_0_63_0_6_n_1),
        .DOC(n9m_reg_0_63_0_6_n_2),
        .DOD(n9m_reg_0_63_0_6_n_3),
        .DOE(n9m_reg_0_63_0_6_n_4),
        .DOF(n9m_reg_0_63_0_6_n_5),
        .DOG(n9m_reg_0_63_0_6_n_6),
        .DOH(NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39699 n9m_reg_0_63_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[12]),
        .DIB(i1[13]),
        .DIC(i1[14]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_14_20_n_0),
        .DOB(n9m_reg_0_63_14_20_n_1),
        .DOC(n9m_reg_0_63_14_20_n_2),
        .DOD(n9m_reg_0_63_14_20_n_3),
        .DOE(n9m_reg_0_63_14_20_n_4),
        .DOF(n9m_reg_0_63_14_20_n_5),
        .DOG(n9m_reg_0_63_14_20_n_6),
        .DOH(NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39700 n9m_reg_0_63_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_21_27_n_0),
        .DOB(n9m_reg_0_63_21_27_n_1),
        .DOC(n9m_reg_0_63_21_27_n_2),
        .DOD(n9m_reg_0_63_21_27_n_3),
        .DOE(n9m_reg_0_63_21_27_n_4),
        .DOF(n9m_reg_0_63_21_27_n_5),
        .DOG(n9m_reg_0_63_21_27_n_6),
        .DOH(NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39701 n9m_reg_0_63_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_28_31_n_0),
        .DOB(n9m_reg_0_63_28_31_n_1),
        .DOC(n9m_reg_0_63_28_31_n_2),
        .DOD(n9m_reg_0_63_28_31_n_3),
        .DOE(NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39702 n9m_reg_0_63_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[22]),
        .DIC(i1[7]),
        .DID(i1[8]),
        .DIE(i1[9]),
        .DIF(i1[10]),
        .DIG(i1[11]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_7_13_n_0),
        .DOB(n9m_reg_0_63_7_13_n_1),
        .DOC(n9m_reg_0_63_7_13_n_2),
        .DOD(n9m_reg_0_63_7_13_n_3),
        .DOE(n9m_reg_0_63_7_13_n_4),
        .DOF(n9m_reg_0_63_7_13_n_5),
        .DOG(n9m_reg_0_63_7_13_n_6),
        .DOH(NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39703 n9m_reg_64_127_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[14]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_0_6_n_0),
        .DOB(n9m_reg_64_127_0_6_n_1),
        .DOC(n9m_reg_64_127_0_6_n_2),
        .DOD(n9m_reg_64_127_0_6_n_3),
        .DOE(n9m_reg_64_127_0_6_n_4),
        .DOF(n9m_reg_64_127_0_6_n_5),
        .DOG(n9m_reg_64_127_0_6_n_6),
        .DOH(NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39704 n9m_reg_64_127_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[12]),
        .DIB(i1[13]),
        .DIC(i1[14]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_14_20_n_0),
        .DOB(n9m_reg_64_127_14_20_n_1),
        .DOC(n9m_reg_64_127_14_20_n_2),
        .DOD(n9m_reg_64_127_14_20_n_3),
        .DOE(n9m_reg_64_127_14_20_n_4),
        .DOF(n9m_reg_64_127_14_20_n_5),
        .DOG(n9m_reg_64_127_14_20_n_6),
        .DOH(NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39705 n9m_reg_64_127_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_21_27_n_0),
        .DOB(n9m_reg_64_127_21_27_n_1),
        .DOC(n9m_reg_64_127_21_27_n_2),
        .DOD(n9m_reg_64_127_21_27_n_3),
        .DOE(n9m_reg_64_127_21_27_n_4),
        .DOF(n9m_reg_64_127_21_27_n_5),
        .DOG(n9m_reg_64_127_21_27_n_6),
        .DOH(NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39706 n9m_reg_64_127_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_28_31_n_0),
        .DOB(n9m_reg_64_127_28_31_n_1),
        .DOC(n9m_reg_64_127_28_31_n_2),
        .DOD(n9m_reg_64_127_28_31_n_3),
        .DOE(NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39707 n9m_reg_64_127_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[22]),
        .DIC(i1[7]),
        .DID(i1[8]),
        .DIE(i1[9]),
        .DIF(i1[10]),
        .DIG(i1[11]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_7_13_n_0),
        .DOB(n9m_reg_64_127_7_13_n_1),
        .DOC(n9m_reg_64_127_7_13_n_2),
        .DOD(n9m_reg_64_127_7_13_n_3),
        .DOE(n9m_reg_64_127_7_13_n_4),
        .DOF(n9m_reg_64_127_7_13_n_5),
        .DOG(n9m_reg_64_127_7_13_n_6),
        .DOH(NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_26" *) 
module switch_elements_cf_fft_512_8_26_5
   (\n9_reg[0] ,
    n4,
    \n1_reg[0] ,
    i8,
    rst_i,
    enable_i,
    clk_i,
    i1);
  output [15:0]\n9_reg[0] ;
  output n4;
  input \n1_reg[0] ;
  input [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [6:0]n11a;
  wire [5:0]n11a__0;
  wire n11m_reg_0_63_0_6_n_0;
  wire n11m_reg_0_63_0_6_n_1;
  wire n11m_reg_0_63_0_6_n_2;
  wire n11m_reg_0_63_0_6_n_3;
  wire n11m_reg_0_63_0_6_n_4;
  wire n11m_reg_0_63_0_6_n_5;
  wire n11m_reg_0_63_0_6_n_6;
  wire n11m_reg_0_63_14_20_n_0;
  wire n11m_reg_0_63_14_20_n_1;
  wire n11m_reg_0_63_14_20_n_2;
  wire n11m_reg_0_63_14_20_n_3;
  wire n11m_reg_0_63_14_20_n_4;
  wire n11m_reg_0_63_14_20_n_5;
  wire n11m_reg_0_63_14_20_n_6;
  wire n11m_reg_0_63_21_27_n_0;
  wire n11m_reg_0_63_21_27_n_1;
  wire n11m_reg_0_63_21_27_n_2;
  wire n11m_reg_0_63_21_27_n_3;
  wire n11m_reg_0_63_21_27_n_4;
  wire n11m_reg_0_63_21_27_n_5;
  wire n11m_reg_0_63_21_27_n_6;
  wire n11m_reg_0_63_28_31_n_0;
  wire n11m_reg_0_63_28_31_n_1;
  wire n11m_reg_0_63_28_31_n_2;
  wire n11m_reg_0_63_28_31_n_3;
  wire n11m_reg_0_63_7_13_n_0;
  wire n11m_reg_0_63_7_13_n_1;
  wire n11m_reg_0_63_7_13_n_2;
  wire n11m_reg_0_63_7_13_n_3;
  wire n11m_reg_0_63_7_13_n_4;
  wire n11m_reg_0_63_7_13_n_5;
  wire n11m_reg_0_63_7_13_n_6;
  wire \n1[0]_i_2__3_n_0 ;
  wire \n1[0]_i_3__3_n_0 ;
  wire \n1[10]_i_2__3_n_0 ;
  wire \n1[10]_i_3__3_n_0 ;
  wire \n1[11]_i_2__3_n_0 ;
  wire \n1[11]_i_3__3_n_0 ;
  wire \n1[12]_i_2__3_n_0 ;
  wire \n1[12]_i_3__3_n_0 ;
  wire \n1[13]_i_2__3_n_0 ;
  wire \n1[13]_i_3__3_n_0 ;
  wire \n1[14]_i_2__3_n_0 ;
  wire \n1[14]_i_3__3_n_0 ;
  wire \n1[15]_i_2__3_n_0 ;
  wire \n1[15]_i_3__3_n_0 ;
  wire \n1[1]_i_2__3_n_0 ;
  wire \n1[1]_i_3__3_n_0 ;
  wire \n1[2]_i_2__3_n_0 ;
  wire \n1[2]_i_3__3_n_0 ;
  wire \n1[3]_i_2__3_n_0 ;
  wire \n1[3]_i_3__3_n_0 ;
  wire \n1[4]_i_2__3_n_0 ;
  wire \n1[4]_i_3__3_n_0 ;
  wire \n1[5]_i_2__3_n_0 ;
  wire \n1[5]_i_3__3_n_0 ;
  wire \n1[6]_i_2__3_n_0 ;
  wire \n1[6]_i_3__3_n_0 ;
  wire \n1[7]_i_2__3_n_0 ;
  wire \n1[7]_i_3__3_n_0 ;
  wire \n1[8]_i_2__3_n_0 ;
  wire \n1[8]_i_3__3_n_0 ;
  wire \n1[9]_i_2__3_n_0 ;
  wire \n1[9]_i_3__3_n_0 ;
  wire \n1_reg[0] ;
  wire [6:0]n2__0;
  wire \n3[6]_i_2__4_n_0 ;
  wire [6:0]n3_reg;
  wire n4;
  wire \n5[0]_i_2__4_n_0 ;
  wire [15:0]\n9_reg[0] ;
  wire n9m_reg_0_63_0_6_n_0;
  wire n9m_reg_0_63_0_6_n_1;
  wire n9m_reg_0_63_0_6_n_2;
  wire n9m_reg_0_63_0_6_n_3;
  wire n9m_reg_0_63_0_6_n_4;
  wire n9m_reg_0_63_0_6_n_5;
  wire n9m_reg_0_63_0_6_n_6;
  wire n9m_reg_0_63_14_20_n_0;
  wire n9m_reg_0_63_14_20_n_1;
  wire n9m_reg_0_63_14_20_n_2;
  wire n9m_reg_0_63_14_20_n_3;
  wire n9m_reg_0_63_14_20_n_4;
  wire n9m_reg_0_63_14_20_n_5;
  wire n9m_reg_0_63_14_20_n_6;
  wire n9m_reg_0_63_21_27_n_0;
  wire n9m_reg_0_63_21_27_n_1;
  wire n9m_reg_0_63_21_27_n_2;
  wire n9m_reg_0_63_21_27_n_3;
  wire n9m_reg_0_63_21_27_n_4;
  wire n9m_reg_0_63_21_27_n_5;
  wire n9m_reg_0_63_21_27_n_6;
  wire n9m_reg_0_63_28_31_n_0;
  wire n9m_reg_0_63_28_31_n_1;
  wire n9m_reg_0_63_28_31_n_2;
  wire n9m_reg_0_63_28_31_n_3;
  wire n9m_reg_0_63_7_13_n_0;
  wire n9m_reg_0_63_7_13_n_1;
  wire n9m_reg_0_63_7_13_n_2;
  wire n9m_reg_0_63_7_13_n_3;
  wire n9m_reg_0_63_7_13_n_4;
  wire n9m_reg_0_63_7_13_n_5;
  wire n9m_reg_0_63_7_13_n_6;
  wire n9m_reg_64_127_0_6_n_0;
  wire n9m_reg_64_127_0_6_n_1;
  wire n9m_reg_64_127_0_6_n_2;
  wire n9m_reg_64_127_0_6_n_3;
  wire n9m_reg_64_127_0_6_n_4;
  wire n9m_reg_64_127_0_6_n_5;
  wire n9m_reg_64_127_0_6_n_6;
  wire n9m_reg_64_127_14_20_n_0;
  wire n9m_reg_64_127_14_20_n_1;
  wire n9m_reg_64_127_14_20_n_2;
  wire n9m_reg_64_127_14_20_n_3;
  wire n9m_reg_64_127_14_20_n_4;
  wire n9m_reg_64_127_14_20_n_5;
  wire n9m_reg_64_127_14_20_n_6;
  wire n9m_reg_64_127_21_27_n_0;
  wire n9m_reg_64_127_21_27_n_1;
  wire n9m_reg_64_127_21_27_n_2;
  wire n9m_reg_64_127_21_27_n_3;
  wire n9m_reg_64_127_21_27_n_4;
  wire n9m_reg_64_127_21_27_n_5;
  wire n9m_reg_64_127_21_27_n_6;
  wire n9m_reg_64_127_28_31_n_0;
  wire n9m_reg_64_127_28_31_n_1;
  wire n9m_reg_64_127_28_31_n_2;
  wire n9m_reg_64_127_28_31_n_3;
  wire n9m_reg_64_127_7_13_n_0;
  wire n9m_reg_64_127_7_13_n_1;
  wire n9m_reg_64_127_7_13_n_2;
  wire n9m_reg_64_127_7_13_n_3;
  wire n9m_reg_64_127_7_13_n_4;
  wire n9m_reg_64_127_7_13_n_5;
  wire n9m_reg_64_127_7_13_n_6;
  wire rst_i;
  wire NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED;

  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39833 n11m_reg_0_63_0_6
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_0_6_n_0),
        .DOB(n11m_reg_0_63_0_6_n_1),
        .DOC(n11m_reg_0_63_0_6_n_2),
        .DOD(n11m_reg_0_63_0_6_n_3),
        .DOE(n11m_reg_0_63_0_6_n_4),
        .DOF(n11m_reg_0_63_0_6_n_5),
        .DOG(n11m_reg_0_63_0_6_n_6),
        .DOH(NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39834 n11m_reg_0_63_14_20
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_14_20_n_0),
        .DOB(n11m_reg_0_63_14_20_n_1),
        .DOC(n11m_reg_0_63_14_20_n_2),
        .DOD(n11m_reg_0_63_14_20_n_3),
        .DOE(n11m_reg_0_63_14_20_n_4),
        .DOF(n11m_reg_0_63_14_20_n_5),
        .DOG(n11m_reg_0_63_14_20_n_6),
        .DOH(NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39835 n11m_reg_0_63_21_27
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_21_27_n_0),
        .DOB(n11m_reg_0_63_21_27_n_1),
        .DOC(n11m_reg_0_63_21_27_n_2),
        .DOD(n11m_reg_0_63_21_27_n_3),
        .DOE(n11m_reg_0_63_21_27_n_4),
        .DOF(n11m_reg_0_63_21_27_n_5),
        .DOG(n11m_reg_0_63_21_27_n_6),
        .DOH(NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39836 n11m_reg_0_63_28_31
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_28_31_n_0),
        .DOB(n11m_reg_0_63_28_31_n_1),
        .DOC(n11m_reg_0_63_28_31_n_2),
        .DOD(n11m_reg_0_63_28_31_n_3),
        .DOE(NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39837 n11m_reg_0_63_7_13
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n11m_reg_0_63_7_13_n_0),
        .DOB(n11m_reg_0_63_7_13_n_1),
        .DOC(n11m_reg_0_63_7_13_n_2),
        .DOD(n11m_reg_0_63_7_13_n_3),
        .DOE(n11m_reg_0_63_7_13_n_4),
        .DOF(n11m_reg_0_63_7_13_n_5),
        .DOG(n11m_reg_0_63_7_13_n_6),
        .DOH(NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[0]_i_1__3 
       (.I0(n11m_reg_0_63_0_6_n_0),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[0]_i_2__3_n_0 ),
        .I4(\n1[0]_i_3__3_n_0 ),
        .O(\n9_reg[0] [0]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[0]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_0),
        .O(\n1[0]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[0]_i_3__3 
       (.I0(n11m_reg_0_63_14_20_n_2),
        .I1(n9m_reg_64_127_14_20_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[0]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[10]_i_1__3 
       (.I0(n11m_reg_0_63_7_13_n_3),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[10]_i_2__3_n_0 ),
        .I4(\n1[10]_i_3__3_n_0 ),
        .O(\n9_reg[0] [10]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[10]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_3),
        .O(\n1[10]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[10]_i_3__3 
       (.I0(n11m_reg_0_63_21_27_n_5),
        .I1(n9m_reg_64_127_21_27_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[10]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[11]_i_1__3 
       (.I0(n11m_reg_0_63_7_13_n_4),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[11]_i_2__3_n_0 ),
        .I4(\n1[11]_i_3__3_n_0 ),
        .O(\n9_reg[0] [11]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[11]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_4),
        .O(\n1[11]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[11]_i_3__3 
       (.I0(n11m_reg_0_63_21_27_n_6),
        .I1(n9m_reg_64_127_21_27_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[11]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[12]_i_1__3 
       (.I0(n11m_reg_0_63_7_13_n_5),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[12]_i_2__3_n_0 ),
        .I4(\n1[12]_i_3__3_n_0 ),
        .O(\n9_reg[0] [12]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[12]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_5),
        .O(\n1[12]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[12]_i_3__3 
       (.I0(n11m_reg_0_63_28_31_n_0),
        .I1(n9m_reg_64_127_28_31_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[12]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[13]_i_1__3 
       (.I0(n11m_reg_0_63_7_13_n_6),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[13]_i_2__3_n_0 ),
        .I4(\n1[13]_i_3__3_n_0 ),
        .O(\n9_reg[0] [13]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[13]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_6),
        .O(\n1[13]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[13]_i_3__3 
       (.I0(n11m_reg_0_63_28_31_n_1),
        .I1(n9m_reg_64_127_28_31_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[13]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[14]_i_1__3 
       (.I0(n11m_reg_0_63_14_20_n_0),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[14]_i_2__3_n_0 ),
        .I4(\n1[14]_i_3__3_n_0 ),
        .O(\n9_reg[0] [14]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[14]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_0),
        .O(\n1[14]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[14]_i_3__3 
       (.I0(n11m_reg_0_63_28_31_n_2),
        .I1(n9m_reg_64_127_28_31_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[14]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[15]_i_1__3 
       (.I0(n11m_reg_0_63_14_20_n_1),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[15]_i_2__3_n_0 ),
        .I4(\n1[15]_i_3__3_n_0 ),
        .O(\n9_reg[0] [15]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[15]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_1),
        .O(\n1[15]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[15]_i_3__3 
       (.I0(n11m_reg_0_63_28_31_n_3),
        .I1(n9m_reg_64_127_28_31_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[15]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[1]_i_1__3 
       (.I0(n11m_reg_0_63_0_6_n_1),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[1]_i_2__3_n_0 ),
        .I4(\n1[1]_i_3__3_n_0 ),
        .O(\n9_reg[0] [1]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[1]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_1),
        .O(\n1[1]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[1]_i_3__3 
       (.I0(n11m_reg_0_63_14_20_n_3),
        .I1(n9m_reg_64_127_14_20_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[1]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[2]_i_1__3 
       (.I0(n11m_reg_0_63_0_6_n_2),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[2]_i_2__3_n_0 ),
        .I4(\n1[2]_i_3__3_n_0 ),
        .O(\n9_reg[0] [2]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[2]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_2),
        .O(\n1[2]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[2]_i_3__3 
       (.I0(n11m_reg_0_63_14_20_n_4),
        .I1(n9m_reg_64_127_14_20_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[2]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[3]_i_1__3 
       (.I0(n11m_reg_0_63_0_6_n_3),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[3]_i_2__3_n_0 ),
        .I4(\n1[3]_i_3__3_n_0 ),
        .O(\n9_reg[0] [3]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[3]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_3),
        .O(\n1[3]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[3]_i_3__3 
       (.I0(n11m_reg_0_63_14_20_n_5),
        .I1(n9m_reg_64_127_14_20_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[3]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[4]_i_1__3 
       (.I0(n11m_reg_0_63_0_6_n_4),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[4]_i_2__3_n_0 ),
        .I4(\n1[4]_i_3__3_n_0 ),
        .O(\n9_reg[0] [4]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[4]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_4),
        .O(\n1[4]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[4]_i_3__3 
       (.I0(n11m_reg_0_63_14_20_n_6),
        .I1(n9m_reg_64_127_14_20_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[4]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[5]_i_1__3 
       (.I0(n11m_reg_0_63_0_6_n_5),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[5]_i_2__3_n_0 ),
        .I4(\n1[5]_i_3__3_n_0 ),
        .O(\n9_reg[0] [5]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[5]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_5),
        .O(\n1[5]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[5]_i_3__3 
       (.I0(n11m_reg_0_63_21_27_n_0),
        .I1(n9m_reg_64_127_21_27_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[5]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[6]_i_1__3 
       (.I0(n11m_reg_0_63_0_6_n_6),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[6]_i_2__3_n_0 ),
        .I4(\n1[6]_i_3__3_n_0 ),
        .O(\n9_reg[0] [6]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[6]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_6),
        .O(\n1[6]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[6]_i_3__3 
       (.I0(n11m_reg_0_63_21_27_n_1),
        .I1(n9m_reg_64_127_21_27_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[6]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[7]_i_1__3 
       (.I0(n11m_reg_0_63_7_13_n_0),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[7]_i_2__3_n_0 ),
        .I4(\n1[7]_i_3__3_n_0 ),
        .O(\n9_reg[0] [7]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[7]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_0),
        .O(\n1[7]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[7]_i_3__3 
       (.I0(n11m_reg_0_63_21_27_n_2),
        .I1(n9m_reg_64_127_21_27_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[7]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[8]_i_1__3 
       (.I0(n11m_reg_0_63_7_13_n_1),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[8]_i_2__3_n_0 ),
        .I4(\n1[8]_i_3__3_n_0 ),
        .O(\n9_reg[0] [8]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[8]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_1),
        .O(\n1[8]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[8]_i_3__3 
       (.I0(n11m_reg_0_63_21_27_n_3),
        .I1(n9m_reg_64_127_21_27_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[8]_i_3__3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[9]_i_1__3 
       (.I0(n11m_reg_0_63_7_13_n_2),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[9]_i_2__3_n_0 ),
        .I4(\n1[9]_i_3__3_n_0 ),
        .O(\n9_reg[0] [9]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[9]_i_2__3 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_2),
        .O(\n1[9]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[9]_i_3__3 
       (.I0(n11m_reg_0_63_21_27_n_4),
        .I1(n9m_reg_64_127_21_27_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[9]_i_3__3_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__9 
       (.I0(n3_reg[0]),
        .O(n2__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__9 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__9 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__9 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__9 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__0[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__9 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__0[5]));
  LUT3 #(
    .INIT(8'hD2)) 
    \n3[6]_i_1__4 
       (.I0(n3_reg[5]),
        .I1(\n3[6]_i_2__4_n_0 ),
        .I2(n3_reg[6]),
        .O(n2__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \n3[6]_i_2__4 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(\n3[6]_i_2__4_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[6]),
        .Q(n3_reg[6]),
        .R(rst_i));
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \n5[0]_i_1__4 
       (.I0(n3_reg[0]),
        .I1(\n5[0]_i_2__4_n_0 ),
        .I2(i8),
        .O(n4));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \n5[0]_i_2__4 
       (.I0(n3_reg[3]),
        .I1(n3_reg[4]),
        .I2(n3_reg[1]),
        .I3(n3_reg[2]),
        .I4(n3_reg[6]),
        .I5(n3_reg[5]),
        .O(\n5[0]_i_2__4_n_0 ));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[6]),
        .Q(n11a[6]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39838 n9m_reg_0_63_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_0_6_n_0),
        .DOB(n9m_reg_0_63_0_6_n_1),
        .DOC(n9m_reg_0_63_0_6_n_2),
        .DOD(n9m_reg_0_63_0_6_n_3),
        .DOE(n9m_reg_0_63_0_6_n_4),
        .DOF(n9m_reg_0_63_0_6_n_5),
        .DOG(n9m_reg_0_63_0_6_n_6),
        .DOH(NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39839 n9m_reg_0_63_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_14_20_n_0),
        .DOB(n9m_reg_0_63_14_20_n_1),
        .DOC(n9m_reg_0_63_14_20_n_2),
        .DOD(n9m_reg_0_63_14_20_n_3),
        .DOE(n9m_reg_0_63_14_20_n_4),
        .DOF(n9m_reg_0_63_14_20_n_5),
        .DOG(n9m_reg_0_63_14_20_n_6),
        .DOH(NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39840 n9m_reg_0_63_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_21_27_n_0),
        .DOB(n9m_reg_0_63_21_27_n_1),
        .DOC(n9m_reg_0_63_21_27_n_2),
        .DOD(n9m_reg_0_63_21_27_n_3),
        .DOE(n9m_reg_0_63_21_27_n_4),
        .DOF(n9m_reg_0_63_21_27_n_5),
        .DOG(n9m_reg_0_63_21_27_n_6),
        .DOH(NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39841 n9m_reg_0_63_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_28_31_n_0),
        .DOB(n9m_reg_0_63_28_31_n_1),
        .DOC(n9m_reg_0_63_28_31_n_2),
        .DOD(n9m_reg_0_63_28_31_n_3),
        .DOE(NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39842 n9m_reg_0_63_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_7_13_n_0),
        .DOB(n9m_reg_0_63_7_13_n_1),
        .DOC(n9m_reg_0_63_7_13_n_2),
        .DOD(n9m_reg_0_63_7_13_n_3),
        .DOE(n9m_reg_0_63_7_13_n_4),
        .DOF(n9m_reg_0_63_7_13_n_5),
        .DOG(n9m_reg_0_63_7_13_n_6),
        .DOH(NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39843 n9m_reg_64_127_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_0_6_n_0),
        .DOB(n9m_reg_64_127_0_6_n_1),
        .DOC(n9m_reg_64_127_0_6_n_2),
        .DOD(n9m_reg_64_127_0_6_n_3),
        .DOE(n9m_reg_64_127_0_6_n_4),
        .DOF(n9m_reg_64_127_0_6_n_5),
        .DOG(n9m_reg_64_127_0_6_n_6),
        .DOH(NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39844 n9m_reg_64_127_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_14_20_n_0),
        .DOB(n9m_reg_64_127_14_20_n_1),
        .DOC(n9m_reg_64_127_14_20_n_2),
        .DOD(n9m_reg_64_127_14_20_n_3),
        .DOE(n9m_reg_64_127_14_20_n_4),
        .DOF(n9m_reg_64_127_14_20_n_5),
        .DOG(n9m_reg_64_127_14_20_n_6),
        .DOH(NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39845 n9m_reg_64_127_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_21_27_n_0),
        .DOB(n9m_reg_64_127_21_27_n_1),
        .DOC(n9m_reg_64_127_21_27_n_2),
        .DOD(n9m_reg_64_127_21_27_n_3),
        .DOE(n9m_reg_64_127_21_27_n_4),
        .DOF(n9m_reg_64_127_21_27_n_5),
        .DOG(n9m_reg_64_127_21_27_n_6),
        .DOH(NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39846 n9m_reg_64_127_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_28_31_n_0),
        .DOB(n9m_reg_64_127_28_31_n_1),
        .DOC(n9m_reg_64_127_28_31_n_2),
        .DOD(n9m_reg_64_127_28_31_n_3),
        .DOE(NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39847 n9m_reg_64_127_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_7_13_n_0),
        .DOB(n9m_reg_64_127_7_13_n_1),
        .DOC(n9m_reg_64_127_7_13_n_2),
        .DOD(n9m_reg_64_127_7_13_n_3),
        .DOE(n9m_reg_64_127_7_13_n_4),
        .DOF(n9m_reg_64_127_7_13_n_5),
        .DOG(n9m_reg_64_127_7_13_n_6),
        .DOH(NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_26" *) 
module switch_elements_cf_fft_512_8_26_8
   (\n9_reg[0] ,
    n4,
    \n1_reg[0] ,
    i8,
    rst_i,
    enable_i,
    clk_i,
    i1);
  output [15:0]\n9_reg[0] ;
  output n4;
  input \n1_reg[0] ;
  input [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [31:0]n11;
  wire [6:0]n11a;
  wire [5:0]n11a__0;
  wire \n1[0]_i_2__2_n_0 ;
  wire \n1[0]_i_3__2_n_0 ;
  wire \n1[10]_i_2__2_n_0 ;
  wire \n1[10]_i_3__2_n_0 ;
  wire \n1[11]_i_2__2_n_0 ;
  wire \n1[11]_i_3__2_n_0 ;
  wire \n1[12]_i_2__2_n_0 ;
  wire \n1[12]_i_3__2_n_0 ;
  wire \n1[13]_i_2__2_n_0 ;
  wire \n1[13]_i_3__2_n_0 ;
  wire \n1[14]_i_2__2_n_0 ;
  wire \n1[14]_i_3__2_n_0 ;
  wire \n1[15]_i_2__2_n_0 ;
  wire \n1[15]_i_3__2_n_0 ;
  wire \n1[1]_i_2__2_n_0 ;
  wire \n1[1]_i_3__2_n_0 ;
  wire \n1[2]_i_2__2_n_0 ;
  wire \n1[2]_i_3__2_n_0 ;
  wire \n1[3]_i_2__2_n_0 ;
  wire \n1[3]_i_3__2_n_0 ;
  wire \n1[4]_i_2__2_n_0 ;
  wire \n1[4]_i_3__2_n_0 ;
  wire \n1[5]_i_2__2_n_0 ;
  wire \n1[5]_i_3__2_n_0 ;
  wire \n1[6]_i_2__2_n_0 ;
  wire \n1[6]_i_3__2_n_0 ;
  wire \n1[7]_i_2__2_n_0 ;
  wire \n1[7]_i_3__2_n_0 ;
  wire \n1[8]_i_2__2_n_0 ;
  wire \n1[8]_i_3__2_n_0 ;
  wire \n1[9]_i_2__2_n_0 ;
  wire \n1[9]_i_3__2_n_0 ;
  wire \n1_reg[0] ;
  wire [6:0]n2__0;
  wire \n3[6]_i_2__3_n_0 ;
  wire [6:0]n3_reg;
  wire n4;
  wire \n5[0]_i_2__3_n_0 ;
  wire [15:0]\n9_reg[0] ;
  wire n9m_reg_0_63_0_6_n_0;
  wire n9m_reg_0_63_0_6_n_1;
  wire n9m_reg_0_63_0_6_n_2;
  wire n9m_reg_0_63_0_6_n_3;
  wire n9m_reg_0_63_0_6_n_4;
  wire n9m_reg_0_63_0_6_n_5;
  wire n9m_reg_0_63_0_6_n_6;
  wire n9m_reg_0_63_14_20_n_0;
  wire n9m_reg_0_63_14_20_n_1;
  wire n9m_reg_0_63_14_20_n_2;
  wire n9m_reg_0_63_14_20_n_3;
  wire n9m_reg_0_63_14_20_n_4;
  wire n9m_reg_0_63_14_20_n_5;
  wire n9m_reg_0_63_14_20_n_6;
  wire n9m_reg_0_63_21_27_n_0;
  wire n9m_reg_0_63_21_27_n_1;
  wire n9m_reg_0_63_21_27_n_2;
  wire n9m_reg_0_63_21_27_n_3;
  wire n9m_reg_0_63_21_27_n_4;
  wire n9m_reg_0_63_21_27_n_5;
  wire n9m_reg_0_63_21_27_n_6;
  wire n9m_reg_0_63_28_31_n_0;
  wire n9m_reg_0_63_28_31_n_1;
  wire n9m_reg_0_63_28_31_n_2;
  wire n9m_reg_0_63_28_31_n_3;
  wire n9m_reg_0_63_7_13_n_0;
  wire n9m_reg_0_63_7_13_n_1;
  wire n9m_reg_0_63_7_13_n_2;
  wire n9m_reg_0_63_7_13_n_3;
  wire n9m_reg_0_63_7_13_n_4;
  wire n9m_reg_0_63_7_13_n_5;
  wire n9m_reg_0_63_7_13_n_6;
  wire n9m_reg_64_127_0_6_n_0;
  wire n9m_reg_64_127_0_6_n_1;
  wire n9m_reg_64_127_0_6_n_2;
  wire n9m_reg_64_127_0_6_n_3;
  wire n9m_reg_64_127_0_6_n_4;
  wire n9m_reg_64_127_0_6_n_5;
  wire n9m_reg_64_127_0_6_n_6;
  wire n9m_reg_64_127_14_20_n_0;
  wire n9m_reg_64_127_14_20_n_1;
  wire n9m_reg_64_127_14_20_n_2;
  wire n9m_reg_64_127_14_20_n_3;
  wire n9m_reg_64_127_14_20_n_4;
  wire n9m_reg_64_127_14_20_n_5;
  wire n9m_reg_64_127_14_20_n_6;
  wire n9m_reg_64_127_21_27_n_0;
  wire n9m_reg_64_127_21_27_n_1;
  wire n9m_reg_64_127_21_27_n_2;
  wire n9m_reg_64_127_21_27_n_3;
  wire n9m_reg_64_127_21_27_n_4;
  wire n9m_reg_64_127_21_27_n_5;
  wire n9m_reg_64_127_21_27_n_6;
  wire n9m_reg_64_127_28_31_n_0;
  wire n9m_reg_64_127_28_31_n_1;
  wire n9m_reg_64_127_28_31_n_2;
  wire n9m_reg_64_127_28_31_n_3;
  wire n9m_reg_64_127_7_13_n_0;
  wire n9m_reg_64_127_7_13_n_1;
  wire n9m_reg_64_127_7_13_n_2;
  wire n9m_reg_64_127_7_13_n_3;
  wire n9m_reg_64_127_7_13_n_4;
  wire n9m_reg_64_127_7_13_n_5;
  wire n9m_reg_64_127_7_13_n_6;
  wire rst_i;
  wire NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED;

  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39808 n11m_reg_0_63_0_6
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n11[0]),
        .DOB(n11[1]),
        .DOC(n11[2]),
        .DOD(n11[3]),
        .DOE(n11[4]),
        .DOF(n11[5]),
        .DOG(n11[6]),
        .DOH(NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39809 n11m_reg_0_63_14_20
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n11[14]),
        .DOB(n11[15]),
        .DOC(n11[16]),
        .DOD(n11[17]),
        .DOE(n11[18]),
        .DOF(n11[19]),
        .DOG(n11[20]),
        .DOH(NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39810 n11m_reg_0_63_21_27
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n11[21]),
        .DOB(n11[22]),
        .DOC(n11[23]),
        .DOD(n11[24]),
        .DOE(n11[25]),
        .DOF(n11[26]),
        .DOG(n11[27]),
        .DOH(NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39811 n11m_reg_0_63_28_31
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n11[28]),
        .DOB(n11[29]),
        .DOC(n11[30]),
        .DOD(n11[31]),
        .DOE(NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39812 n11m_reg_0_63_7_13
       (.ADDRA(n11a__0),
        .ADDRB(n11a__0),
        .ADDRC(n11a__0),
        .ADDRD(n11a__0),
        .ADDRE(n11a__0),
        .ADDRF(n11a__0),
        .ADDRG(n11a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n11[7]),
        .DOB(n11[8]),
        .DOC(n11[9]),
        .DOD(n11[10]),
        .DOE(n11[11]),
        .DOF(n11[12]),
        .DOG(n11[13]),
        .DOH(NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[0]_i_1__2 
       (.I0(n11[0]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[0]_i_2__2_n_0 ),
        .I4(\n1[0]_i_3__2_n_0 ),
        .O(\n9_reg[0] [0]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[0]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_0),
        .O(\n1[0]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[0]_i_3__2 
       (.I0(n11[16]),
        .I1(n9m_reg_64_127_14_20_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[0]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[10]_i_1__2 
       (.I0(n11[10]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[10]_i_2__2_n_0 ),
        .I4(\n1[10]_i_3__2_n_0 ),
        .O(\n9_reg[0] [10]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[10]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_3),
        .O(\n1[10]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[10]_i_3__2 
       (.I0(n11[26]),
        .I1(n9m_reg_64_127_21_27_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[10]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[11]_i_1__2 
       (.I0(n11[11]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[11]_i_2__2_n_0 ),
        .I4(\n1[11]_i_3__2_n_0 ),
        .O(\n9_reg[0] [11]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[11]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_4),
        .O(\n1[11]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[11]_i_3__2 
       (.I0(n11[27]),
        .I1(n9m_reg_64_127_21_27_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[11]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[12]_i_1__2 
       (.I0(n11[12]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[12]_i_2__2_n_0 ),
        .I4(\n1[12]_i_3__2_n_0 ),
        .O(\n9_reg[0] [12]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[12]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_5),
        .O(\n1[12]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[12]_i_3__2 
       (.I0(n11[28]),
        .I1(n9m_reg_64_127_28_31_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[12]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[13]_i_1__2 
       (.I0(n11[13]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[13]_i_2__2_n_0 ),
        .I4(\n1[13]_i_3__2_n_0 ),
        .O(\n9_reg[0] [13]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[13]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_6),
        .O(\n1[13]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[13]_i_3__2 
       (.I0(n11[29]),
        .I1(n9m_reg_64_127_28_31_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[13]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[14]_i_1__2 
       (.I0(n11[14]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[14]_i_2__2_n_0 ),
        .I4(\n1[14]_i_3__2_n_0 ),
        .O(\n9_reg[0] [14]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[14]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_0),
        .O(\n1[14]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[14]_i_3__2 
       (.I0(n11[30]),
        .I1(n9m_reg_64_127_28_31_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[14]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[15]_i_1__2 
       (.I0(n11[15]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[15]_i_2__2_n_0 ),
        .I4(\n1[15]_i_3__2_n_0 ),
        .O(\n9_reg[0] [15]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[15]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_14_20_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_14_20_n_1),
        .O(\n1[15]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[15]_i_3__2 
       (.I0(n11[31]),
        .I1(n9m_reg_64_127_28_31_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_28_31_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[15]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[1]_i_1__2 
       (.I0(n11[1]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[1]_i_2__2_n_0 ),
        .I4(\n1[1]_i_3__2_n_0 ),
        .O(\n9_reg[0] [1]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[1]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_1),
        .O(\n1[1]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[1]_i_3__2 
       (.I0(n11[17]),
        .I1(n9m_reg_64_127_14_20_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[1]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[2]_i_1__2 
       (.I0(n11[2]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[2]_i_2__2_n_0 ),
        .I4(\n1[2]_i_3__2_n_0 ),
        .O(\n9_reg[0] [2]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[2]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_2),
        .O(\n1[2]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[2]_i_3__2 
       (.I0(n11[18]),
        .I1(n9m_reg_64_127_14_20_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[2]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[3]_i_1__2 
       (.I0(n11[3]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[3]_i_2__2_n_0 ),
        .I4(\n1[3]_i_3__2_n_0 ),
        .O(\n9_reg[0] [3]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[3]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_3),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_3),
        .O(\n1[3]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[3]_i_3__2 
       (.I0(n11[19]),
        .I1(n9m_reg_64_127_14_20_n_5),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_5),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[3]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[4]_i_1__2 
       (.I0(n11[4]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[4]_i_2__2_n_0 ),
        .I4(\n1[4]_i_3__2_n_0 ),
        .O(\n9_reg[0] [4]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[4]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_4),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_4),
        .O(\n1[4]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[4]_i_3__2 
       (.I0(n11[20]),
        .I1(n9m_reg_64_127_14_20_n_6),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_14_20_n_6),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[4]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[5]_i_1__2 
       (.I0(n11[5]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[5]_i_2__2_n_0 ),
        .I4(\n1[5]_i_3__2_n_0 ),
        .O(\n9_reg[0] [5]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[5]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_5),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_5),
        .O(\n1[5]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[5]_i_3__2 
       (.I0(n11[21]),
        .I1(n9m_reg_64_127_21_27_n_0),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_0),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[5]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[6]_i_1__2 
       (.I0(n11[6]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[6]_i_2__2_n_0 ),
        .I4(\n1[6]_i_3__2_n_0 ),
        .O(\n9_reg[0] [6]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[6]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_0_6_n_6),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_0_6_n_6),
        .O(\n1[6]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[6]_i_3__2 
       (.I0(n11[22]),
        .I1(n9m_reg_64_127_21_27_n_1),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_1),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[6]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[7]_i_1__2 
       (.I0(n11[7]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[7]_i_2__2_n_0 ),
        .I4(\n1[7]_i_3__2_n_0 ),
        .O(\n9_reg[0] [7]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[7]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_0),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_0),
        .O(\n1[7]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[7]_i_3__2 
       (.I0(n11[23]),
        .I1(n9m_reg_64_127_21_27_n_2),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_2),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[7]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[8]_i_1__2 
       (.I0(n11[8]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[8]_i_2__2_n_0 ),
        .I4(\n1[8]_i_3__2_n_0 ),
        .O(\n9_reg[0] [8]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[8]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_1),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_1),
        .O(\n1[8]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[8]_i_3__2 
       (.I0(n11[24]),
        .I1(n9m_reg_64_127_21_27_n_3),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_3),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[8]_i_3__2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF80)) 
    \n1[9]_i_1__2 
       (.I0(n11[9]),
        .I1(\n1_reg[0] ),
        .I2(i8),
        .I3(\n1[9]_i_2__2_n_0 ),
        .I4(\n1[9]_i_3__2_n_0 ),
        .O(\n9_reg[0] [9]));
  LUT5 #(
    .INIT(32'h44400040)) 
    \n1[9]_i_2__2 
       (.I0(\n1_reg[0] ),
        .I1(i8),
        .I2(n9m_reg_0_63_7_13_n_2),
        .I3(n11a[6]),
        .I4(n9m_reg_64_127_7_13_n_2),
        .O(\n1[9]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAACFC0)) 
    \n1[9]_i_3__2 
       (.I0(n11[25]),
        .I1(n9m_reg_64_127_21_27_n_4),
        .I2(n11a[6]),
        .I3(n9m_reg_0_63_21_27_n_4),
        .I4(\n1_reg[0] ),
        .I5(i8),
        .O(\n1[9]_i_3__2_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__7 
       (.I0(n3_reg[0]),
        .O(n2__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__7 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__7 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__7 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__7 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__0[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__7 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__0[5]));
  LUT3 #(
    .INIT(8'hD2)) 
    \n3[6]_i_1__3 
       (.I0(n3_reg[5]),
        .I1(\n3[6]_i_2__3_n_0 ),
        .I2(n3_reg[6]),
        .O(n2__0[6]));
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \n3[6]_i_2__3 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(\n3[6]_i_2__3_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[6]),
        .Q(n3_reg[6]),
        .R(rst_i));
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \n5[0]_i_1__3 
       (.I0(n3_reg[0]),
        .I1(\n5[0]_i_2__3_n_0 ),
        .I2(i8),
        .O(n4));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \n5[0]_i_2__3 
       (.I0(n3_reg[3]),
        .I1(n3_reg[4]),
        .I2(n3_reg[1]),
        .I3(n3_reg[2]),
        .I4(n3_reg[6]),
        .I5(n3_reg[5]),
        .O(\n5[0]_i_2__3_n_0 ));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[6]),
        .Q(n11a[6]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39813 n9m_reg_0_63_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_0_6_n_0),
        .DOB(n9m_reg_0_63_0_6_n_1),
        .DOC(n9m_reg_0_63_0_6_n_2),
        .DOD(n9m_reg_0_63_0_6_n_3),
        .DOE(n9m_reg_0_63_0_6_n_4),
        .DOF(n9m_reg_0_63_0_6_n_5),
        .DOG(n9m_reg_0_63_0_6_n_6),
        .DOH(NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39814 n9m_reg_0_63_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_14_20_n_0),
        .DOB(n9m_reg_0_63_14_20_n_1),
        .DOC(n9m_reg_0_63_14_20_n_2),
        .DOD(n9m_reg_0_63_14_20_n_3),
        .DOE(n9m_reg_0_63_14_20_n_4),
        .DOF(n9m_reg_0_63_14_20_n_5),
        .DOG(n9m_reg_0_63_14_20_n_6),
        .DOH(NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39815 n9m_reg_0_63_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_21_27_n_0),
        .DOB(n9m_reg_0_63_21_27_n_1),
        .DOC(n9m_reg_0_63_21_27_n_2),
        .DOD(n9m_reg_0_63_21_27_n_3),
        .DOE(n9m_reg_0_63_21_27_n_4),
        .DOF(n9m_reg_0_63_21_27_n_5),
        .DOG(n9m_reg_0_63_21_27_n_6),
        .DOH(NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39816 n9m_reg_0_63_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_28_31_n_0),
        .DOB(n9m_reg_0_63_28_31_n_1),
        .DOC(n9m_reg_0_63_28_31_n_2),
        .DOD(n9m_reg_0_63_28_31_n_3),
        .DOE(NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39817 n9m_reg_0_63_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_7_13_n_0),
        .DOB(n9m_reg_0_63_7_13_n_1),
        .DOC(n9m_reg_0_63_7_13_n_2),
        .DOD(n9m_reg_0_63_7_13_n_3),
        .DOE(n9m_reg_0_63_7_13_n_4),
        .DOF(n9m_reg_0_63_7_13_n_5),
        .DOG(n9m_reg_0_63_7_13_n_6),
        .DOH(NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39818 n9m_reg_64_127_0_6
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_0_6_n_0),
        .DOB(n9m_reg_64_127_0_6_n_1),
        .DOC(n9m_reg_64_127_0_6_n_2),
        .DOD(n9m_reg_64_127_0_6_n_3),
        .DOE(n9m_reg_64_127_0_6_n_4),
        .DOF(n9m_reg_64_127_0_6_n_5),
        .DOG(n9m_reg_64_127_0_6_n_6),
        .DOH(NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39819 n9m_reg_64_127_14_20
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_14_20_n_0),
        .DOB(n9m_reg_64_127_14_20_n_1),
        .DOC(n9m_reg_64_127_14_20_n_2),
        .DOD(n9m_reg_64_127_14_20_n_3),
        .DOE(n9m_reg_64_127_14_20_n_4),
        .DOF(n9m_reg_64_127_14_20_n_5),
        .DOG(n9m_reg_64_127_14_20_n_6),
        .DOH(NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39820 n9m_reg_64_127_21_27
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_21_27_n_0),
        .DOB(n9m_reg_64_127_21_27_n_1),
        .DOC(n9m_reg_64_127_21_27_n_2),
        .DOD(n9m_reg_64_127_21_27_n_3),
        .DOE(n9m_reg_64_127_21_27_n_4),
        .DOF(n9m_reg_64_127_21_27_n_5),
        .DOG(n9m_reg_64_127_21_27_n_6),
        .DOH(NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39821 n9m_reg_64_127_28_31
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_28_31_n_0),
        .DOB(n9m_reg_64_127_28_31_n_1),
        .DOC(n9m_reg_64_127_28_31_n_2),
        .DOD(n9m_reg_64_127_28_31_n_3),
        .DOE(NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39822 n9m_reg_64_127_7_13
       (.ADDRA(n11a[5:0]),
        .ADDRB(n11a[5:0]),
        .ADDRC(n11a[5:0]),
        .ADDRD(n11a[5:0]),
        .ADDRE(n11a[5:0]),
        .ADDRF(n11a[5:0]),
        .ADDRG(n11a[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_7_13_n_0),
        .DOB(n9m_reg_64_127_7_13_n_1),
        .DOC(n9m_reg_64_127_7_13_n_2),
        .DOD(n9m_reg_64_127_7_13_n_3),
        .DOE(n9m_reg_64_127_7_13_n_4),
        .DOF(n9m_reg_64_127_7_13_n_5),
        .DOG(n9m_reg_64_127_7_13_n_6),
        .DOH(NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_27" *) 
module switch_elements_cf_fft_512_8_27
   (\n9_reg[0]_0 ,
    s8_3,
    rst_i,
    enable_i,
    clk_i,
    i8,
    i1);
  output \n9_reg[0]_0 ;
  output [15:0]s8_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [0:0]i8;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [5:0]n2__1;
  wire [5:0]n3_reg;
  wire n6m_reg_0_63_0_6_n_0;
  wire n6m_reg_0_63_0_6_n_1;
  wire n6m_reg_0_63_0_6_n_2;
  wire n6m_reg_0_63_0_6_n_3;
  wire n6m_reg_0_63_0_6_n_4;
  wire n6m_reg_0_63_0_6_n_5;
  wire n6m_reg_0_63_0_6_n_6;
  wire n6m_reg_0_63_14_20_n_0;
  wire n6m_reg_0_63_14_20_n_1;
  wire n6m_reg_0_63_14_20_n_2;
  wire n6m_reg_0_63_14_20_n_3;
  wire n6m_reg_0_63_14_20_n_4;
  wire n6m_reg_0_63_14_20_n_5;
  wire n6m_reg_0_63_14_20_n_6;
  wire n6m_reg_0_63_21_27_n_0;
  wire n6m_reg_0_63_21_27_n_1;
  wire n6m_reg_0_63_21_27_n_2;
  wire n6m_reg_0_63_21_27_n_3;
  wire n6m_reg_0_63_21_27_n_4;
  wire n6m_reg_0_63_21_27_n_5;
  wire n6m_reg_0_63_21_27_n_6;
  wire n6m_reg_0_63_28_31_n_0;
  wire n6m_reg_0_63_28_31_n_1;
  wire n6m_reg_0_63_28_31_n_2;
  wire n6m_reg_0_63_28_31_n_3;
  wire n6m_reg_0_63_7_13_n_0;
  wire n6m_reg_0_63_7_13_n_1;
  wire n6m_reg_0_63_7_13_n_2;
  wire n6m_reg_0_63_7_13_n_3;
  wire n6m_reg_0_63_7_13_n_4;
  wire n6m_reg_0_63_7_13_n_5;
  wire n6m_reg_0_63_7_13_n_6;
  wire [31:0]n8;
  wire [5:0]n8a;
  wire [5:0]n8a__0;
  wire \n9_reg[0]_0 ;
  wire rst_i;
  wire [15:0]s8_3;
  wire NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED;

  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__0_i_1__5
       (.I0(n8[14]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_0),
        .I4(n8[30]),
        .I5(n6m_reg_0_63_28_31_n_2),
        .O(s8_3[14]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__1_i_1__5
       (.I0(n8[13]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_6),
        .I4(n8[29]),
        .I5(n6m_reg_0_63_28_31_n_1),
        .O(s8_3[13]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__2_i_1__5
       (.I0(n8[12]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_5),
        .I4(n8[28]),
        .I5(n6m_reg_0_63_28_31_n_0),
        .O(s8_3[12]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__3_i_1__5
       (.I0(n8[11]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_4),
        .I4(n8[27]),
        .I5(n6m_reg_0_63_21_27_n_6),
        .O(s8_3[11]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__4_i_1__5
       (.I0(n8[10]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_3),
        .I4(n8[26]),
        .I5(n6m_reg_0_63_21_27_n_5),
        .O(s8_3[10]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__5_i_1__5
       (.I0(n8[9]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_2),
        .I4(n8[25]),
        .I5(n6m_reg_0_63_21_27_n_4),
        .O(s8_3[9]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__6_i_1__5
       (.I0(n8[8]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_1),
        .I4(n8[24]),
        .I5(n6m_reg_0_63_21_27_n_3),
        .O(s8_3[8]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22_i_1__5
       (.I0(n8[15]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_1),
        .I4(n8[31]),
        .I5(n6m_reg_0_63_28_31_n_3),
        .O(s8_3[15]));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__14 
       (.I0(n3_reg[0]),
        .O(n2__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__14 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__1[1]));
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__14 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__1[2]));
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__14 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__1[3]));
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__14 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__1[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__14 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__1[5]));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[0]_i_1__5 
       (.I0(n8[0]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_0),
        .I4(n8[16]),
        .I5(n6m_reg_0_63_14_20_n_2),
        .O(s8_3[0]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[1]_i_1__5 
       (.I0(n8[1]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_1),
        .I4(n8[17]),
        .I5(n6m_reg_0_63_14_20_n_3),
        .O(s8_3[1]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[2]_i_1__5 
       (.I0(n8[2]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_2),
        .I4(n8[18]),
        .I5(n6m_reg_0_63_14_20_n_4),
        .O(s8_3[2]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[3]_i_1__5 
       (.I0(n8[3]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_3),
        .I4(n8[19]),
        .I5(n6m_reg_0_63_14_20_n_5),
        .O(s8_3[3]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[4]_i_1__5 
       (.I0(n8[4]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_4),
        .I4(n8[20]),
        .I5(n6m_reg_0_63_14_20_n_6),
        .O(s8_3[4]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[5]_i_1__5 
       (.I0(n8[5]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_5),
        .I4(n8[21]),
        .I5(n6m_reg_0_63_21_27_n_0),
        .O(s8_3[5]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[6]_i_1__5 
       (.I0(n8[6]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_6),
        .I4(n8[22]),
        .I5(n6m_reg_0_63_21_27_n_1),
        .O(s8_3[6]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[7]_i_1__5 
       (.I0(n8[7]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_0),
        .I4(n8[23]),
        .I5(n6m_reg_0_63_21_27_n_2),
        .O(s8_3[7]));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a[5]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39898 n6m_reg_0_63_0_6
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_0_6_n_0),
        .DOB(n6m_reg_0_63_0_6_n_1),
        .DOC(n6m_reg_0_63_0_6_n_2),
        .DOD(n6m_reg_0_63_0_6_n_3),
        .DOE(n6m_reg_0_63_0_6_n_4),
        .DOF(n6m_reg_0_63_0_6_n_5),
        .DOG(n6m_reg_0_63_0_6_n_6),
        .DOH(NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39899 n6m_reg_0_63_14_20
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_14_20_n_0),
        .DOB(n6m_reg_0_63_14_20_n_1),
        .DOC(n6m_reg_0_63_14_20_n_2),
        .DOD(n6m_reg_0_63_14_20_n_3),
        .DOE(n6m_reg_0_63_14_20_n_4),
        .DOF(n6m_reg_0_63_14_20_n_5),
        .DOG(n6m_reg_0_63_14_20_n_6),
        .DOH(NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39900 n6m_reg_0_63_21_27
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_21_27_n_0),
        .DOB(n6m_reg_0_63_21_27_n_1),
        .DOC(n6m_reg_0_63_21_27_n_2),
        .DOD(n6m_reg_0_63_21_27_n_3),
        .DOE(n6m_reg_0_63_21_27_n_4),
        .DOF(n6m_reg_0_63_21_27_n_5),
        .DOG(n6m_reg_0_63_21_27_n_6),
        .DOH(NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39901 n6m_reg_0_63_28_31
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_28_31_n_0),
        .DOB(n6m_reg_0_63_28_31_n_1),
        .DOC(n6m_reg_0_63_28_31_n_2),
        .DOD(n6m_reg_0_63_28_31_n_3),
        .DOE(NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39902 n6m_reg_0_63_7_13
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_7_13_n_0),
        .DOB(n6m_reg_0_63_7_13_n_1),
        .DOC(n6m_reg_0_63_7_13_n_2),
        .DOD(n6m_reg_0_63_7_13_n_3),
        .DOE(n6m_reg_0_63_7_13_n_4),
        .DOF(n6m_reg_0_63_7_13_n_5),
        .DOG(n6m_reg_0_63_7_13_n_6),
        .DOH(NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39903 n8m_reg_0_63_0_6
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n8[0]),
        .DOB(n8[1]),
        .DOC(n8[2]),
        .DOD(n8[3]),
        .DOE(n8[4]),
        .DOF(n8[5]),
        .DOG(n8[6]),
        .DOH(NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39904 n8m_reg_0_63_14_20
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n8[14]),
        .DOB(n8[15]),
        .DOC(n8[16]),
        .DOD(n8[17]),
        .DOE(n8[18]),
        .DOF(n8[19]),
        .DOG(n8[20]),
        .DOH(NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39905 n8m_reg_0_63_21_27
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n8[21]),
        .DOB(n8[22]),
        .DOC(n8[23]),
        .DOD(n8[24]),
        .DOE(n8[25]),
        .DOF(n8[26]),
        .DOG(n8[27]),
        .DOH(NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39906 n8m_reg_0_63_28_31
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n8[28]),
        .DOB(n8[29]),
        .DOC(n8[30]),
        .DOD(n8[31]),
        .DOE(NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39907 n8m_reg_0_63_7_13
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n8[7]),
        .DOB(n8[8]),
        .DOC(n8[9]),
        .DOD(n8[10]),
        .DOE(n8[11]),
        .DOF(n8[12]),
        .DOG(n8[13]),
        .DOH(NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(1'b1),
        .Q(\n9_reg[0]_0 ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_27" *) 
module switch_elements_cf_fft_512_8_27_12
   (\n9_reg[0]_0 ,
    s4_3,
    rst_i,
    enable_i,
    clk_i,
    i8,
    i1);
  output \n9_reg[0]_0 ;
  output [15:0]s4_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [0:0]i8;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [5:0]n2__1;
  wire [5:0]n3_reg;
  wire n6m_reg_0_63_0_6_n_0;
  wire n6m_reg_0_63_0_6_n_1;
  wire n6m_reg_0_63_0_6_n_2;
  wire n6m_reg_0_63_0_6_n_3;
  wire n6m_reg_0_63_0_6_n_4;
  wire n6m_reg_0_63_0_6_n_5;
  wire n6m_reg_0_63_0_6_n_6;
  wire n6m_reg_0_63_14_20_n_0;
  wire n6m_reg_0_63_14_20_n_1;
  wire n6m_reg_0_63_14_20_n_2;
  wire n6m_reg_0_63_14_20_n_3;
  wire n6m_reg_0_63_14_20_n_4;
  wire n6m_reg_0_63_14_20_n_5;
  wire n6m_reg_0_63_14_20_n_6;
  wire n6m_reg_0_63_21_27_n_0;
  wire n6m_reg_0_63_21_27_n_1;
  wire n6m_reg_0_63_21_27_n_2;
  wire n6m_reg_0_63_21_27_n_3;
  wire n6m_reg_0_63_21_27_n_4;
  wire n6m_reg_0_63_21_27_n_5;
  wire n6m_reg_0_63_21_27_n_6;
  wire n6m_reg_0_63_28_31_n_0;
  wire n6m_reg_0_63_28_31_n_1;
  wire n6m_reg_0_63_28_31_n_2;
  wire n6m_reg_0_63_28_31_n_3;
  wire n6m_reg_0_63_7_13_n_0;
  wire n6m_reg_0_63_7_13_n_1;
  wire n6m_reg_0_63_7_13_n_2;
  wire n6m_reg_0_63_7_13_n_3;
  wire n6m_reg_0_63_7_13_n_4;
  wire n6m_reg_0_63_7_13_n_5;
  wire n6m_reg_0_63_7_13_n_6;
  wire [31:0]n8;
  wire [5:0]n8a;
  wire [5:0]n8a__0;
  wire \n9_reg[0]_0 ;
  wire rst_i;
  wire [15:0]s4_3;
  wire NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED;

  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__0_i_1__1
       (.I0(n8[14]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_0),
        .I4(n8[30]),
        .I5(n6m_reg_0_63_28_31_n_2),
        .O(s4_3[14]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__1_i_1__1
       (.I0(n8[13]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_6),
        .I4(n8[29]),
        .I5(n6m_reg_0_63_28_31_n_1),
        .O(s4_3[13]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__2_i_1__1
       (.I0(n8[12]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_5),
        .I4(n8[28]),
        .I5(n6m_reg_0_63_28_31_n_0),
        .O(s4_3[12]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__3_i_1__1
       (.I0(n8[11]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_4),
        .I4(n8[27]),
        .I5(n6m_reg_0_63_21_27_n_6),
        .O(s4_3[11]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__4_i_1__1
       (.I0(n8[10]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_3),
        .I4(n8[26]),
        .I5(n6m_reg_0_63_21_27_n_5),
        .O(s4_3[10]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__5_i_1__1
       (.I0(n8[9]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_2),
        .I4(n8[25]),
        .I5(n6m_reg_0_63_21_27_n_4),
        .O(s4_3[9]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__6_i_1__1
       (.I0(n8[8]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_1),
        .I4(n8[24]),
        .I5(n6m_reg_0_63_21_27_n_3),
        .O(s4_3[8]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22_i_1__1
       (.I0(n8[15]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_1),
        .I4(n8[31]),
        .I5(n6m_reg_0_63_28_31_n_3),
        .O(s4_3[15]));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__6 
       (.I0(n3_reg[0]),
        .O(n2__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__6 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__1[1]));
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__6 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__1[2]));
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__6 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__1[3]));
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__6 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__1[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__6 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__1[5]));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[0]_i_1__1 
       (.I0(n8[0]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_0),
        .I4(n8[16]),
        .I5(n6m_reg_0_63_14_20_n_2),
        .O(s4_3[0]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[1]_i_1__1 
       (.I0(n8[1]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_1),
        .I4(n8[17]),
        .I5(n6m_reg_0_63_14_20_n_3),
        .O(s4_3[1]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[2]_i_1__1 
       (.I0(n8[2]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_2),
        .I4(n8[18]),
        .I5(n6m_reg_0_63_14_20_n_4),
        .O(s4_3[2]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[3]_i_1__1 
       (.I0(n8[3]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_3),
        .I4(n8[19]),
        .I5(n6m_reg_0_63_14_20_n_5),
        .O(s4_3[3]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[4]_i_1__1 
       (.I0(n8[4]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_4),
        .I4(n8[20]),
        .I5(n6m_reg_0_63_14_20_n_6),
        .O(s4_3[4]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[5]_i_1__1 
       (.I0(n8[5]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_5),
        .I4(n8[21]),
        .I5(n6m_reg_0_63_21_27_n_0),
        .O(s4_3[5]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[6]_i_1__1 
       (.I0(n8[6]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_6),
        .I4(n8[22]),
        .I5(n6m_reg_0_63_21_27_n_1),
        .O(s4_3[6]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[7]_i_1__1 
       (.I0(n8[7]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_0),
        .I4(n8[23]),
        .I5(n6m_reg_0_63_21_27_n_2),
        .O(s4_3[7]));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a[5]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39798 n6m_reg_0_63_0_6
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[0]),
        .DIB(i1[1]),
        .DIC(i1[2]),
        .DID(i1[3]),
        .DIE(i1[4]),
        .DIF(i1[5]),
        .DIG(i1[6]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_0_6_n_0),
        .DOB(n6m_reg_0_63_0_6_n_1),
        .DOC(n6m_reg_0_63_0_6_n_2),
        .DOD(n6m_reg_0_63_0_6_n_3),
        .DOE(n6m_reg_0_63_0_6_n_4),
        .DOF(n6m_reg_0_63_0_6_n_5),
        .DOG(n6m_reg_0_63_0_6_n_6),
        .DOH(NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39799 n6m_reg_0_63_14_20
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[0]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_14_20_n_0),
        .DOB(n6m_reg_0_63_14_20_n_1),
        .DOC(n6m_reg_0_63_14_20_n_2),
        .DOD(n6m_reg_0_63_14_20_n_3),
        .DOE(n6m_reg_0_63_14_20_n_4),
        .DOF(n6m_reg_0_63_14_20_n_5),
        .DOG(n6m_reg_0_63_14_20_n_6),
        .DOH(NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39800 n6m_reg_0_63_21_27
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_21_27_n_0),
        .DOB(n6m_reg_0_63_21_27_n_1),
        .DOC(n6m_reg_0_63_21_27_n_2),
        .DOD(n6m_reg_0_63_21_27_n_3),
        .DOE(n6m_reg_0_63_21_27_n_4),
        .DOF(n6m_reg_0_63_21_27_n_5),
        .DOG(n6m_reg_0_63_21_27_n_6),
        .DOH(NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39801 n6m_reg_0_63_28_31
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_28_31_n_0),
        .DOB(n6m_reg_0_63_28_31_n_1),
        .DOC(n6m_reg_0_63_28_31_n_2),
        .DOD(n6m_reg_0_63_28_31_n_3),
        .DOE(NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39802 n6m_reg_0_63_7_13
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[7]),
        .DIB(i1[22]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_7_13_n_0),
        .DOB(n6m_reg_0_63_7_13_n_1),
        .DOC(n6m_reg_0_63_7_13_n_2),
        .DOD(n6m_reg_0_63_7_13_n_3),
        .DOE(n6m_reg_0_63_7_13_n_4),
        .DOF(n6m_reg_0_63_7_13_n_5),
        .DOG(n6m_reg_0_63_7_13_n_6),
        .DOH(NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39803 n8m_reg_0_63_0_6
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[0]),
        .DIB(i1[1]),
        .DIC(i1[2]),
        .DID(i1[3]),
        .DIE(i1[4]),
        .DIF(i1[5]),
        .DIG(i1[6]),
        .DIH(1'b0),
        .DOA(n8[0]),
        .DOB(n8[1]),
        .DOC(n8[2]),
        .DOD(n8[3]),
        .DOE(n8[4]),
        .DOF(n8[5]),
        .DOG(n8[6]),
        .DOH(NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39804 n8m_reg_0_63_14_20
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[0]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n8[14]),
        .DOB(n8[15]),
        .DOC(n8[16]),
        .DOD(n8[17]),
        .DOE(n8[18]),
        .DOF(n8[19]),
        .DOG(n8[20]),
        .DOH(NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39805 n8m_reg_0_63_21_27
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n8[21]),
        .DOB(n8[22]),
        .DOC(n8[23]),
        .DOD(n8[24]),
        .DOE(n8[25]),
        .DOF(n8[26]),
        .DOG(n8[27]),
        .DOH(NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39806 n8m_reg_0_63_28_31
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n8[28]),
        .DOB(n8[29]),
        .DOC(n8[30]),
        .DOD(n8[31]),
        .DOE(NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39807 n8m_reg_0_63_7_13
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[7]),
        .DIB(i1[22]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n8[7]),
        .DOB(n8[8]),
        .DOC(n8[9]),
        .DOD(n8[10]),
        .DOE(n8[11]),
        .DOF(n8[12]),
        .DOG(n8[13]),
        .DOH(NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(1'b1),
        .Q(\n9_reg[0]_0 ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_27" *) 
module switch_elements_cf_fft_512_8_27_15
   (\n9_reg[0]_0 ,
    s3_3,
    rst_i,
    enable_i,
    clk_i,
    i8,
    i1);
  output \n9_reg[0]_0 ;
  output [15:0]s3_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [0:0]i8;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [5:0]n2__1;
  wire [5:0]n3_reg;
  wire n6m_reg_0_63_0_6_n_0;
  wire n6m_reg_0_63_0_6_n_1;
  wire n6m_reg_0_63_0_6_n_2;
  wire n6m_reg_0_63_0_6_n_3;
  wire n6m_reg_0_63_0_6_n_4;
  wire n6m_reg_0_63_0_6_n_5;
  wire n6m_reg_0_63_0_6_n_6;
  wire n6m_reg_0_63_14_20_n_0;
  wire n6m_reg_0_63_14_20_n_1;
  wire n6m_reg_0_63_14_20_n_2;
  wire n6m_reg_0_63_14_20_n_3;
  wire n6m_reg_0_63_14_20_n_4;
  wire n6m_reg_0_63_14_20_n_5;
  wire n6m_reg_0_63_14_20_n_6;
  wire n6m_reg_0_63_21_27_n_0;
  wire n6m_reg_0_63_21_27_n_1;
  wire n6m_reg_0_63_21_27_n_2;
  wire n6m_reg_0_63_21_27_n_3;
  wire n6m_reg_0_63_21_27_n_4;
  wire n6m_reg_0_63_21_27_n_5;
  wire n6m_reg_0_63_21_27_n_6;
  wire n6m_reg_0_63_28_31_n_0;
  wire n6m_reg_0_63_28_31_n_1;
  wire n6m_reg_0_63_28_31_n_2;
  wire n6m_reg_0_63_28_31_n_3;
  wire n6m_reg_0_63_7_13_n_0;
  wire n6m_reg_0_63_7_13_n_1;
  wire n6m_reg_0_63_7_13_n_2;
  wire n6m_reg_0_63_7_13_n_3;
  wire n6m_reg_0_63_7_13_n_4;
  wire n6m_reg_0_63_7_13_n_5;
  wire n6m_reg_0_63_7_13_n_6;
  wire [31:0]n8;
  wire [5:0]n8a;
  wire [5:0]n8a__0;
  wire \n9_reg[0]_0 ;
  wire rst_i;
  wire [15:0]s3_3;
  wire NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED;

  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__0_i_1__0
       (.I0(n8[14]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_0),
        .I4(n8[30]),
        .I5(n6m_reg_0_63_28_31_n_2),
        .O(s3_3[14]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__1_i_1__0
       (.I0(n8[13]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_6),
        .I4(n8[29]),
        .I5(n6m_reg_0_63_28_31_n_1),
        .O(s3_3[13]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__2_i_1__0
       (.I0(n8[12]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_5),
        .I4(n8[28]),
        .I5(n6m_reg_0_63_28_31_n_0),
        .O(s3_3[12]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__3_i_1__0
       (.I0(n8[11]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_4),
        .I4(n8[27]),
        .I5(n6m_reg_0_63_21_27_n_6),
        .O(s3_3[11]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__4_i_1__0
       (.I0(n8[10]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_3),
        .I4(n8[26]),
        .I5(n6m_reg_0_63_21_27_n_5),
        .O(s3_3[10]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__5_i_1__0
       (.I0(n8[9]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_2),
        .I4(n8[25]),
        .I5(n6m_reg_0_63_21_27_n_4),
        .O(s3_3[9]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__6_i_1__0
       (.I0(n8[8]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_1),
        .I4(n8[24]),
        .I5(n6m_reg_0_63_21_27_n_3),
        .O(s3_3[8]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22_i_1__0
       (.I0(n8[15]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_1),
        .I4(n8[31]),
        .I5(n6m_reg_0_63_28_31_n_3),
        .O(s3_3[15]));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__4 
       (.I0(n3_reg[0]),
        .O(n2__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__4 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__1[1]));
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__4 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__1[2]));
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__4 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__1[3]));
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__4 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__1[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__4 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__1[5]));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[0]_i_1__0 
       (.I0(n8[0]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_0),
        .I4(n8[16]),
        .I5(n6m_reg_0_63_14_20_n_2),
        .O(s3_3[0]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[1]_i_1__0 
       (.I0(n8[1]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_1),
        .I4(n8[17]),
        .I5(n6m_reg_0_63_14_20_n_3),
        .O(s3_3[1]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[2]_i_1__0 
       (.I0(n8[2]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_2),
        .I4(n8[18]),
        .I5(n6m_reg_0_63_14_20_n_4),
        .O(s3_3[2]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[3]_i_1__0 
       (.I0(n8[3]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_3),
        .I4(n8[19]),
        .I5(n6m_reg_0_63_14_20_n_5),
        .O(s3_3[3]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[4]_i_1__0 
       (.I0(n8[4]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_4),
        .I4(n8[20]),
        .I5(n6m_reg_0_63_14_20_n_6),
        .O(s3_3[4]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[5]_i_1__0 
       (.I0(n8[5]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_5),
        .I4(n8[21]),
        .I5(n6m_reg_0_63_21_27_n_0),
        .O(s3_3[5]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[6]_i_1__0 
       (.I0(n8[6]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_6),
        .I4(n8[22]),
        .I5(n6m_reg_0_63_21_27_n_1),
        .O(s3_3[6]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[7]_i_1__0 
       (.I0(n8[7]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_0),
        .I4(n8[23]),
        .I5(n6m_reg_0_63_21_27_n_2),
        .O(s3_3[7]));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a[5]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39773 n6m_reg_0_63_0_6
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[0]),
        .DIB(i1[1]),
        .DIC(i1[2]),
        .DID(i1[3]),
        .DIE(i1[4]),
        .DIF(i1[5]),
        .DIG(i1[6]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_0_6_n_0),
        .DOB(n6m_reg_0_63_0_6_n_1),
        .DOC(n6m_reg_0_63_0_6_n_2),
        .DOD(n6m_reg_0_63_0_6_n_3),
        .DOE(n6m_reg_0_63_0_6_n_4),
        .DOF(n6m_reg_0_63_0_6_n_5),
        .DOG(n6m_reg_0_63_0_6_n_6),
        .DOH(NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39774 n6m_reg_0_63_14_20
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[0]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_14_20_n_0),
        .DOB(n6m_reg_0_63_14_20_n_1),
        .DOC(n6m_reg_0_63_14_20_n_2),
        .DOD(n6m_reg_0_63_14_20_n_3),
        .DOE(n6m_reg_0_63_14_20_n_4),
        .DOF(n6m_reg_0_63_14_20_n_5),
        .DOG(n6m_reg_0_63_14_20_n_6),
        .DOH(NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39775 n6m_reg_0_63_21_27
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_21_27_n_0),
        .DOB(n6m_reg_0_63_21_27_n_1),
        .DOC(n6m_reg_0_63_21_27_n_2),
        .DOD(n6m_reg_0_63_21_27_n_3),
        .DOE(n6m_reg_0_63_21_27_n_4),
        .DOF(n6m_reg_0_63_21_27_n_5),
        .DOG(n6m_reg_0_63_21_27_n_6),
        .DOH(NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39776 n6m_reg_0_63_28_31
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_28_31_n_0),
        .DOB(n6m_reg_0_63_28_31_n_1),
        .DOC(n6m_reg_0_63_28_31_n_2),
        .DOD(n6m_reg_0_63_28_31_n_3),
        .DOE(NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39777 n6m_reg_0_63_7_13
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[7]),
        .DIB(i1[22]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_7_13_n_0),
        .DOB(n6m_reg_0_63_7_13_n_1),
        .DOC(n6m_reg_0_63_7_13_n_2),
        .DOD(n6m_reg_0_63_7_13_n_3),
        .DOE(n6m_reg_0_63_7_13_n_4),
        .DOF(n6m_reg_0_63_7_13_n_5),
        .DOG(n6m_reg_0_63_7_13_n_6),
        .DOH(NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39778 n8m_reg_0_63_0_6
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[0]),
        .DIB(i1[1]),
        .DIC(i1[2]),
        .DID(i1[3]),
        .DIE(i1[4]),
        .DIF(i1[5]),
        .DIG(i1[6]),
        .DIH(1'b0),
        .DOA(n8[0]),
        .DOB(n8[1]),
        .DOC(n8[2]),
        .DOD(n8[3]),
        .DOE(n8[4]),
        .DOF(n8[5]),
        .DOG(n8[6]),
        .DOH(NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39779 n8m_reg_0_63_14_20
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[0]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n8[14]),
        .DOB(n8[15]),
        .DOC(n8[16]),
        .DOD(n8[17]),
        .DOE(n8[18]),
        .DOF(n8[19]),
        .DOG(n8[20]),
        .DOH(NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39780 n8m_reg_0_63_21_27
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n8[21]),
        .DOB(n8[22]),
        .DOC(n8[23]),
        .DOD(n8[24]),
        .DOE(n8[25]),
        .DOF(n8[26]),
        .DOG(n8[27]),
        .DOH(NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39781 n8m_reg_0_63_28_31
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n8[28]),
        .DOB(n8[29]),
        .DOC(n8[30]),
        .DOD(n8[31]),
        .DOE(NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39782 n8m_reg_0_63_7_13
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[7]),
        .DIB(i1[22]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n8[7]),
        .DOB(n8[8]),
        .DOC(n8[9]),
        .DOD(n8[10]),
        .DOE(n8[11]),
        .DOF(n8[12]),
        .DOG(n8[13]),
        .DOH(NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(1'b1),
        .Q(\n9_reg[0]_0 ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_27" *) 
module switch_elements_cf_fft_512_8_27_17
   (\n9_reg[0]_0 ,
    s2_3,
    rst_i,
    enable_i,
    clk_i,
    i8,
    i1);
  output \n9_reg[0]_0 ;
  output [15:0]s2_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [0:0]i8;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [5:0]n2__1;
  wire [5:0]n3_reg;
  wire n6m_reg_0_63_0_6_n_0;
  wire n6m_reg_0_63_0_6_n_1;
  wire n6m_reg_0_63_0_6_n_2;
  wire n6m_reg_0_63_0_6_n_3;
  wire n6m_reg_0_63_0_6_n_4;
  wire n6m_reg_0_63_0_6_n_5;
  wire n6m_reg_0_63_0_6_n_6;
  wire n6m_reg_0_63_14_20_n_0;
  wire n6m_reg_0_63_14_20_n_1;
  wire n6m_reg_0_63_14_20_n_2;
  wire n6m_reg_0_63_14_20_n_3;
  wire n6m_reg_0_63_14_20_n_4;
  wire n6m_reg_0_63_14_20_n_5;
  wire n6m_reg_0_63_14_20_n_6;
  wire n6m_reg_0_63_21_27_n_0;
  wire n6m_reg_0_63_21_27_n_1;
  wire n6m_reg_0_63_21_27_n_2;
  wire n6m_reg_0_63_21_27_n_3;
  wire n6m_reg_0_63_21_27_n_4;
  wire n6m_reg_0_63_21_27_n_5;
  wire n6m_reg_0_63_21_27_n_6;
  wire n6m_reg_0_63_28_31_n_0;
  wire n6m_reg_0_63_28_31_n_1;
  wire n6m_reg_0_63_28_31_n_2;
  wire n6m_reg_0_63_28_31_n_3;
  wire n6m_reg_0_63_7_13_n_0;
  wire n6m_reg_0_63_7_13_n_1;
  wire n6m_reg_0_63_7_13_n_2;
  wire n6m_reg_0_63_7_13_n_3;
  wire n6m_reg_0_63_7_13_n_4;
  wire n6m_reg_0_63_7_13_n_5;
  wire n6m_reg_0_63_7_13_n_6;
  wire [31:0]n8;
  wire [5:0]n8a;
  wire [5:0]n8a__0;
  wire \n9_reg[0]_0 ;
  wire rst_i;
  wire [15:0]s2_3;
  wire NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED;

  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__0_i_1
       (.I0(n8[14]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_0),
        .I4(n8[30]),
        .I5(n6m_reg_0_63_28_31_n_2),
        .O(s2_3[14]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__1_i_1
       (.I0(n8[13]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_6),
        .I4(n8[29]),
        .I5(n6m_reg_0_63_28_31_n_1),
        .O(s2_3[13]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__2_i_1
       (.I0(n8[12]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_5),
        .I4(n8[28]),
        .I5(n6m_reg_0_63_28_31_n_0),
        .O(s2_3[12]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__3_i_1
       (.I0(n8[11]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_4),
        .I4(n8[27]),
        .I5(n6m_reg_0_63_21_27_n_6),
        .O(s2_3[11]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__4_i_1
       (.I0(n8[10]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_3),
        .I4(n8[26]),
        .I5(n6m_reg_0_63_21_27_n_5),
        .O(s2_3[10]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__5_i_1
       (.I0(n8[9]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_2),
        .I4(n8[25]),
        .I5(n6m_reg_0_63_21_27_n_4),
        .O(s2_3[9]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__6_i_1
       (.I0(n8[8]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_1),
        .I4(n8[24]),
        .I5(n6m_reg_0_63_21_27_n_3),
        .O(s2_3[8]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22_i_1
       (.I0(n8[15]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_1),
        .I4(n8[31]),
        .I5(n6m_reg_0_63_28_31_n_3),
        .O(s2_3[15]));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__2 
       (.I0(n3_reg[0]),
        .O(n2__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__2 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__1[1]));
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__2 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__1[2]));
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__2 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__1[3]));
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__2 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__1[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__2 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__1[5]));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[0]_i_1 
       (.I0(n8[0]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_0),
        .I4(n8[16]),
        .I5(n6m_reg_0_63_14_20_n_2),
        .O(s2_3[0]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[1]_i_1 
       (.I0(n8[1]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_1),
        .I4(n8[17]),
        .I5(n6m_reg_0_63_14_20_n_3),
        .O(s2_3[1]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[2]_i_1 
       (.I0(n8[2]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_2),
        .I4(n8[18]),
        .I5(n6m_reg_0_63_14_20_n_4),
        .O(s2_3[2]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[3]_i_1 
       (.I0(n8[3]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_3),
        .I4(n8[19]),
        .I5(n6m_reg_0_63_14_20_n_5),
        .O(s2_3[3]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[4]_i_1 
       (.I0(n8[4]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_4),
        .I4(n8[20]),
        .I5(n6m_reg_0_63_14_20_n_6),
        .O(s2_3[4]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[5]_i_1 
       (.I0(n8[5]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_5),
        .I4(n8[21]),
        .I5(n6m_reg_0_63_21_27_n_0),
        .O(s2_3[5]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[6]_i_1 
       (.I0(n8[6]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_6),
        .I4(n8[22]),
        .I5(n6m_reg_0_63_21_27_n_1),
        .O(s2_3[6]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[7]_i_1 
       (.I0(n8[7]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_0),
        .I4(n8[23]),
        .I5(n6m_reg_0_63_21_27_n_2),
        .O(s2_3[7]));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a[5]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39733 n6m_reg_0_63_0_6
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[0]),
        .DIB(i1[1]),
        .DIC(i1[2]),
        .DID(i1[3]),
        .DIE(i1[4]),
        .DIF(i1[5]),
        .DIG(i1[6]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_0_6_n_0),
        .DOB(n6m_reg_0_63_0_6_n_1),
        .DOC(n6m_reg_0_63_0_6_n_2),
        .DOD(n6m_reg_0_63_0_6_n_3),
        .DOE(n6m_reg_0_63_0_6_n_4),
        .DOF(n6m_reg_0_63_0_6_n_5),
        .DOG(n6m_reg_0_63_0_6_n_6),
        .DOH(NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39734 n6m_reg_0_63_14_20
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[0]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_14_20_n_0),
        .DOB(n6m_reg_0_63_14_20_n_1),
        .DOC(n6m_reg_0_63_14_20_n_2),
        .DOD(n6m_reg_0_63_14_20_n_3),
        .DOE(n6m_reg_0_63_14_20_n_4),
        .DOF(n6m_reg_0_63_14_20_n_5),
        .DOG(n6m_reg_0_63_14_20_n_6),
        .DOH(NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39735 n6m_reg_0_63_21_27
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_21_27_n_0),
        .DOB(n6m_reg_0_63_21_27_n_1),
        .DOC(n6m_reg_0_63_21_27_n_2),
        .DOD(n6m_reg_0_63_21_27_n_3),
        .DOE(n6m_reg_0_63_21_27_n_4),
        .DOF(n6m_reg_0_63_21_27_n_5),
        .DOG(n6m_reg_0_63_21_27_n_6),
        .DOH(NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39736 n6m_reg_0_63_28_31
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_28_31_n_0),
        .DOB(n6m_reg_0_63_28_31_n_1),
        .DOC(n6m_reg_0_63_28_31_n_2),
        .DOD(n6m_reg_0_63_28_31_n_3),
        .DOE(NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39737 n6m_reg_0_63_7_13
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[7]),
        .DIB(i1[22]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_7_13_n_0),
        .DOB(n6m_reg_0_63_7_13_n_1),
        .DOC(n6m_reg_0_63_7_13_n_2),
        .DOD(n6m_reg_0_63_7_13_n_3),
        .DOE(n6m_reg_0_63_7_13_n_4),
        .DOF(n6m_reg_0_63_7_13_n_5),
        .DOG(n6m_reg_0_63_7_13_n_6),
        .DOH(NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39738 n8m_reg_0_63_0_6
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[0]),
        .DIB(i1[1]),
        .DIC(i1[2]),
        .DID(i1[3]),
        .DIE(i1[4]),
        .DIF(i1[5]),
        .DIG(i1[6]),
        .DIH(1'b0),
        .DOA(n8[0]),
        .DOB(n8[1]),
        .DOC(n8[2]),
        .DOD(n8[3]),
        .DOE(n8[4]),
        .DOF(n8[5]),
        .DOG(n8[6]),
        .DOH(NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39739 n8m_reg_0_63_14_20
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[0]),
        .DID(i1[15]),
        .DIE(i1[16]),
        .DIF(i1[17]),
        .DIG(i1[18]),
        .DIH(1'b0),
        .DOA(n8[14]),
        .DOB(n8[15]),
        .DOC(n8[16]),
        .DOD(n8[17]),
        .DOE(n8[18]),
        .DOF(n8[19]),
        .DOG(n8[20]),
        .DOH(NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39740 n8m_reg_0_63_21_27
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[19]),
        .DIB(i1[20]),
        .DIC(i1[21]),
        .DID(i1[22]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n8[21]),
        .DOB(n8[22]),
        .DOC(n8[23]),
        .DOD(n8[24]),
        .DOE(n8[25]),
        .DOF(n8[26]),
        .DOG(n8[27]),
        .DOH(NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39741 n8m_reg_0_63_28_31
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n8[28]),
        .DOB(n8[29]),
        .DOC(n8[30]),
        .DOD(n8[31]),
        .DOE(NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s28/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39742 n8m_reg_0_63_7_13
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[7]),
        .DIB(i1[22]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n8[7]),
        .DOB(n8[8]),
        .DOC(n8[9]),
        .DOD(n8[10]),
        .DOE(n8[11]),
        .DOF(n8[12]),
        .DOG(n8[13]),
        .DOH(NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(1'b1),
        .Q(\n9_reg[0]_0 ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_27" *) 
module switch_elements_cf_fft_512_8_27_20
   (p_6_out,
    inf4_s,
    \info_o_reg[27] ,
    enable_s,
    n12,
    i8,
    rst_i,
    enable_i,
    clk_i,
    i1);
  output [11:0]p_6_out;
  output [15:0]inf4_s;
  input [7:0]\info_o_reg[27] ;
  input [15:0]enable_s;
  input n12;
  input [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [15:0]enable_s;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [15:0]inf4_s;
  wire [7:0]\info_o_reg[27] ;
  wire n12;
  wire [5:0]n2__1;
  wire [5:0]n3_reg;
  wire n6m_reg_0_63_0_6_n_0;
  wire n6m_reg_0_63_0_6_n_1;
  wire n6m_reg_0_63_0_6_n_2;
  wire n6m_reg_0_63_0_6_n_3;
  wire n6m_reg_0_63_0_6_n_4;
  wire n6m_reg_0_63_0_6_n_5;
  wire n6m_reg_0_63_0_6_n_6;
  wire n6m_reg_0_63_14_20_n_0;
  wire n6m_reg_0_63_14_20_n_1;
  wire n6m_reg_0_63_14_20_n_2;
  wire n6m_reg_0_63_14_20_n_3;
  wire n6m_reg_0_63_14_20_n_4;
  wire n6m_reg_0_63_14_20_n_5;
  wire n6m_reg_0_63_14_20_n_6;
  wire n6m_reg_0_63_21_27_n_0;
  wire n6m_reg_0_63_21_27_n_1;
  wire n6m_reg_0_63_21_27_n_2;
  wire n6m_reg_0_63_21_27_n_3;
  wire n6m_reg_0_63_21_27_n_4;
  wire n6m_reg_0_63_21_27_n_5;
  wire n6m_reg_0_63_21_27_n_6;
  wire n6m_reg_0_63_28_31_n_0;
  wire n6m_reg_0_63_28_31_n_1;
  wire n6m_reg_0_63_28_31_n_2;
  wire n6m_reg_0_63_28_31_n_3;
  wire n6m_reg_0_63_7_13_n_0;
  wire n6m_reg_0_63_7_13_n_1;
  wire n6m_reg_0_63_7_13_n_2;
  wire n6m_reg_0_63_7_13_n_3;
  wire n6m_reg_0_63_7_13_n_4;
  wire n6m_reg_0_63_7_13_n_5;
  wire n6m_reg_0_63_7_13_n_6;
  wire [31:0]n8;
  wire [5:0]n8a;
  wire [5:0]n8a__0;
  wire [11:0]p_6_out;
  wire rst_i;
  wire NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED;

  LUT3 #(
    .INIT(8'h96)) 
    \info_o[16]_i_1 
       (.I0(inf4_s[0]),
        .I1(enable_s[8]),
        .I2(enable_s[12]),
        .O(p_6_out[0]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[17]_i_1 
       (.I0(inf4_s[1]),
        .I1(enable_s[9]),
        .I2(enable_s[13]),
        .O(p_6_out[1]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[18]_i_1 
       (.I0(inf4_s[2]),
        .I1(enable_s[10]),
        .I2(enable_s[14]),
        .O(p_6_out[2]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[19]_i_1 
       (.I0(inf4_s[3]),
        .I1(enable_s[11]),
        .I2(enable_s[15]),
        .O(p_6_out[3]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[20]_i_1 
       (.I0(inf4_s[4]),
        .I1(\info_o_reg[27] [0]),
        .I2(enable_s[0]),
        .O(p_6_out[4]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[21]_i_1 
       (.I0(inf4_s[5]),
        .I1(\info_o_reg[27] [1]),
        .I2(enable_s[1]),
        .O(p_6_out[5]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[22]_i_1 
       (.I0(inf4_s[6]),
        .I1(\info_o_reg[27] [2]),
        .I2(enable_s[2]),
        .O(p_6_out[6]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[23]_i_1 
       (.I0(inf4_s[7]),
        .I1(\info_o_reg[27] [3]),
        .I2(enable_s[3]),
        .O(p_6_out[7]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[24]_i_1 
       (.I0(inf4_s[8]),
        .I1(\info_o_reg[27] [4]),
        .I2(enable_s[4]),
        .O(p_6_out[8]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[25]_i_1 
       (.I0(inf4_s[9]),
        .I1(\info_o_reg[27] [5]),
        .I2(enable_s[5]),
        .O(p_6_out[9]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[26]_i_1 
       (.I0(inf4_s[10]),
        .I1(\info_o_reg[27] [6]),
        .I2(enable_s[6]),
        .O(p_6_out[10]));
  LUT3 #(
    .INIT(8'h96)) 
    \info_o[27]_i_1 
       (.I0(inf4_s[11]),
        .I1(\info_o_reg[27] [7]),
        .I2(enable_s[7]),
        .O(p_6_out[11]));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__0 
       (.I0(n3_reg[0]),
        .O(n2__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__0 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__1[1]));
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__0 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__1[2]));
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__0 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__1[3]));
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__0 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__1[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__0 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__1[5]));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a[5]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39708 n6m_reg_0_63_0_6
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_0_6_n_0),
        .DOB(n6m_reg_0_63_0_6_n_1),
        .DOC(n6m_reg_0_63_0_6_n_2),
        .DOD(n6m_reg_0_63_0_6_n_3),
        .DOE(n6m_reg_0_63_0_6_n_4),
        .DOF(n6m_reg_0_63_0_6_n_5),
        .DOG(n6m_reg_0_63_0_6_n_6),
        .DOH(NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_0_6_i_1
       (.I0(n8[0]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_0),
        .I4(n8[16]),
        .I5(n6m_reg_0_63_14_20_n_2),
        .O(inf4_s[0]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_0_6_i_2
       (.I0(n8[1]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_1),
        .I4(n8[17]),
        .I5(n6m_reg_0_63_14_20_n_3),
        .O(inf4_s[1]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_0_6_i_3
       (.I0(n8[2]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_2),
        .I4(n8[18]),
        .I5(n6m_reg_0_63_14_20_n_4),
        .O(inf4_s[2]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_0_6_i_4
       (.I0(n8[3]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_3),
        .I4(n8[19]),
        .I5(n6m_reg_0_63_14_20_n_5),
        .O(inf4_s[3]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_0_6_i_5
       (.I0(n8[4]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_4),
        .I4(n8[20]),
        .I5(n6m_reg_0_63_14_20_n_6),
        .O(inf4_s[4]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_0_6_i_6
       (.I0(n8[5]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_5),
        .I4(n8[21]),
        .I5(n6m_reg_0_63_21_27_n_0),
        .O(inf4_s[5]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_0_6_i_7
       (.I0(n8[6]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_6),
        .I4(n8[22]),
        .I5(n6m_reg_0_63_21_27_n_1),
        .O(inf4_s[6]));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39709 n6m_reg_0_63_14_20
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_14_20_n_0),
        .DOB(n6m_reg_0_63_14_20_n_1),
        .DOC(n6m_reg_0_63_14_20_n_2),
        .DOD(n6m_reg_0_63_14_20_n_3),
        .DOE(n6m_reg_0_63_14_20_n_4),
        .DOF(n6m_reg_0_63_14_20_n_5),
        .DOG(n6m_reg_0_63_14_20_n_6),
        .DOH(NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_14_20_i_1
       (.I0(n8[14]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_0),
        .I4(n8[30]),
        .I5(n6m_reg_0_63_28_31_n_2),
        .O(inf4_s[14]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_14_20_i_2
       (.I0(n8[15]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_1),
        .I4(n8[31]),
        .I5(n6m_reg_0_63_28_31_n_3),
        .O(inf4_s[15]));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39710 n6m_reg_0_63_21_27
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_21_27_n_0),
        .DOB(n6m_reg_0_63_21_27_n_1),
        .DOC(n6m_reg_0_63_21_27_n_2),
        .DOD(n6m_reg_0_63_21_27_n_3),
        .DOE(n6m_reg_0_63_21_27_n_4),
        .DOF(n6m_reg_0_63_21_27_n_5),
        .DOG(n6m_reg_0_63_21_27_n_6),
        .DOH(NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39711 n6m_reg_0_63_28_31
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_28_31_n_0),
        .DOB(n6m_reg_0_63_28_31_n_1),
        .DOC(n6m_reg_0_63_28_31_n_2),
        .DOD(n6m_reg_0_63_28_31_n_3),
        .DOE(NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39712 n6m_reg_0_63_7_13
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_7_13_n_0),
        .DOB(n6m_reg_0_63_7_13_n_1),
        .DOC(n6m_reg_0_63_7_13_n_2),
        .DOD(n6m_reg_0_63_7_13_n_3),
        .DOE(n6m_reg_0_63_7_13_n_4),
        .DOF(n6m_reg_0_63_7_13_n_5),
        .DOG(n6m_reg_0_63_7_13_n_6),
        .DOH(NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_7_13_i_1
       (.I0(n8[7]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_0),
        .I4(n8[23]),
        .I5(n6m_reg_0_63_21_27_n_2),
        .O(inf4_s[7]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_7_13_i_2
       (.I0(n8[8]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_1),
        .I4(n8[24]),
        .I5(n6m_reg_0_63_21_27_n_3),
        .O(inf4_s[8]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_7_13_i_3
       (.I0(n8[9]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_2),
        .I4(n8[25]),
        .I5(n6m_reg_0_63_21_27_n_4),
        .O(inf4_s[9]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_7_13_i_4
       (.I0(n8[10]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_3),
        .I4(n8[26]),
        .I5(n6m_reg_0_63_21_27_n_5),
        .O(inf4_s[10]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_7_13_i_5
       (.I0(n8[11]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_4),
        .I4(n8[27]),
        .I5(n6m_reg_0_63_21_27_n_6),
        .O(inf4_s[11]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_7_13_i_6
       (.I0(n8[12]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_5),
        .I4(n8[28]),
        .I5(n6m_reg_0_63_28_31_n_0),
        .O(inf4_s[12]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n6m_reg_0_63_7_13_i_7
       (.I0(n8[13]),
        .I1(n12),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_6),
        .I4(n8[29]),
        .I5(n6m_reg_0_63_28_31_n_1),
        .O(inf4_s[13]));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39713 n8m_reg_0_63_0_6
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n8[0]),
        .DOB(n8[1]),
        .DOC(n8[2]),
        .DOD(n8[3]),
        .DOE(n8[4]),
        .DOF(n8[5]),
        .DOG(n8[6]),
        .DOH(NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39714 n8m_reg_0_63_14_20
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n8[14]),
        .DOB(n8[15]),
        .DOC(n8[16]),
        .DOD(n8[17]),
        .DOE(n8[18]),
        .DOF(n8[19]),
        .DOG(n8[20]),
        .DOH(NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39715 n8m_reg_0_63_21_27
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n8[21]),
        .DOB(n8[22]),
        .DOC(n8[23]),
        .DOD(n8[24]),
        .DOE(n8[25]),
        .DOF(n8[26]),
        .DOG(n8[27]),
        .DOH(NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39716 n8m_reg_0_63_28_31
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n8[28]),
        .DOB(n8[29]),
        .DOC(n8[30]),
        .DOD(n8[31]),
        .DOE(NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s27/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39717 n8m_reg_0_63_7_13
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n8[7]),
        .DOB(n8[8]),
        .DOC(n8[9]),
        .DOD(n8[10]),
        .DOE(n8[11]),
        .DOF(n8[12]),
        .DOG(n8[13]),
        .DOH(NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_27" *) 
module switch_elements_cf_fft_512_8_27_24
   (\n9_reg[0]_0 ,
    s1_3,
    rst_i,
    enable_i,
    clk_i,
    i8,
    i1);
  output \n9_reg[0]_0 ;
  output [15:0]s1_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [0:0]i8;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [5:0]n2__2;
  wire [5:0]n3_reg;
  wire n6m_reg_0_63_0_6_n_0;
  wire n6m_reg_0_63_0_6_n_1;
  wire n6m_reg_0_63_0_6_n_2;
  wire n6m_reg_0_63_0_6_n_3;
  wire n6m_reg_0_63_0_6_n_4;
  wire n6m_reg_0_63_0_6_n_5;
  wire n6m_reg_0_63_0_6_n_6;
  wire n6m_reg_0_63_14_20_n_0;
  wire n6m_reg_0_63_14_20_n_1;
  wire n6m_reg_0_63_14_20_n_2;
  wire n6m_reg_0_63_14_20_n_3;
  wire n6m_reg_0_63_14_20_n_4;
  wire n6m_reg_0_63_14_20_n_5;
  wire n6m_reg_0_63_14_20_n_6;
  wire n6m_reg_0_63_21_27_n_0;
  wire n6m_reg_0_63_21_27_n_1;
  wire n6m_reg_0_63_21_27_n_2;
  wire n6m_reg_0_63_21_27_n_3;
  wire n6m_reg_0_63_21_27_n_4;
  wire n6m_reg_0_63_21_27_n_5;
  wire n6m_reg_0_63_21_27_n_6;
  wire n6m_reg_0_63_28_31_n_0;
  wire n6m_reg_0_63_28_31_n_1;
  wire n6m_reg_0_63_28_31_n_2;
  wire n6m_reg_0_63_28_31_n_3;
  wire n6m_reg_0_63_7_13_n_0;
  wire n6m_reg_0_63_7_13_n_1;
  wire n6m_reg_0_63_7_13_n_2;
  wire n6m_reg_0_63_7_13_n_3;
  wire n6m_reg_0_63_7_13_n_4;
  wire n6m_reg_0_63_7_13_n_5;
  wire n6m_reg_0_63_7_13_n_6;
  wire [5:0]n8a;
  wire [5:0]n8a__0;
  wire n8m_reg_0_63_0_6_n_0;
  wire n8m_reg_0_63_0_6_n_1;
  wire n8m_reg_0_63_0_6_n_2;
  wire n8m_reg_0_63_0_6_n_3;
  wire n8m_reg_0_63_0_6_n_4;
  wire n8m_reg_0_63_0_6_n_5;
  wire n8m_reg_0_63_0_6_n_6;
  wire n8m_reg_0_63_14_20_n_0;
  wire n8m_reg_0_63_14_20_n_1;
  wire n8m_reg_0_63_14_20_n_2;
  wire n8m_reg_0_63_14_20_n_3;
  wire n8m_reg_0_63_14_20_n_4;
  wire n8m_reg_0_63_14_20_n_5;
  wire n8m_reg_0_63_14_20_n_6;
  wire n8m_reg_0_63_21_27_n_0;
  wire n8m_reg_0_63_21_27_n_1;
  wire n8m_reg_0_63_21_27_n_2;
  wire n8m_reg_0_63_21_27_n_3;
  wire n8m_reg_0_63_21_27_n_4;
  wire n8m_reg_0_63_21_27_n_5;
  wire n8m_reg_0_63_21_27_n_6;
  wire n8m_reg_0_63_28_31_n_0;
  wire n8m_reg_0_63_28_31_n_1;
  wire n8m_reg_0_63_28_31_n_2;
  wire n8m_reg_0_63_28_31_n_3;
  wire n8m_reg_0_63_7_13_n_0;
  wire n8m_reg_0_63_7_13_n_1;
  wire n8m_reg_0_63_7_13_n_2;
  wire n8m_reg_0_63_7_13_n_3;
  wire n8m_reg_0_63_7_13_n_4;
  wire n8m_reg_0_63_7_13_n_5;
  wire n8m_reg_0_63_7_13_n_6;
  wire \n9_reg[0]_0 ;
  wire rst_i;
  wire [15:0]s1_3;
  wire NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED;

  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__0_i_1__7
       (.I0(n8m_reg_0_63_14_20_n_0),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_0),
        .I4(n8m_reg_0_63_28_31_n_2),
        .I5(n6m_reg_0_63_28_31_n_2),
        .O(s1_3[14]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__1_i_1__7
       (.I0(n8m_reg_0_63_7_13_n_6),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_6),
        .I4(n8m_reg_0_63_28_31_n_1),
        .I5(n6m_reg_0_63_28_31_n_1),
        .O(s1_3[13]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__2_i_1__7
       (.I0(n8m_reg_0_63_7_13_n_5),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_5),
        .I4(n8m_reg_0_63_28_31_n_0),
        .I5(n6m_reg_0_63_28_31_n_0),
        .O(s1_3[12]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__3_i_1__7
       (.I0(n8m_reg_0_63_7_13_n_4),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_4),
        .I4(n8m_reg_0_63_21_27_n_6),
        .I5(n6m_reg_0_63_21_27_n_6),
        .O(s1_3[11]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__4_i_1__7
       (.I0(n8m_reg_0_63_7_13_n_3),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_3),
        .I4(n8m_reg_0_63_21_27_n_5),
        .I5(n6m_reg_0_63_21_27_n_5),
        .O(s1_3[10]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__5_i_1__7
       (.I0(n8m_reg_0_63_7_13_n_2),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_2),
        .I4(n8m_reg_0_63_21_27_n_4),
        .I5(n6m_reg_0_63_21_27_n_4),
        .O(s1_3[9]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__6_i_1__7
       (.I0(n8m_reg_0_63_7_13_n_1),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_1),
        .I4(n8m_reg_0_63_21_27_n_3),
        .I5(n6m_reg_0_63_21_27_n_3),
        .O(s1_3[8]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22_i_1__7
       (.I0(n8m_reg_0_63_14_20_n_1),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_1),
        .I4(n8m_reg_0_63_28_31_n_3),
        .I5(n6m_reg_0_63_28_31_n_3),
        .O(s1_3[15]));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__18 
       (.I0(n3_reg[0]),
        .O(n2__2[0]));
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__18 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__2[1]));
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__18 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__2[2]));
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__18 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__2[3]));
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__18 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__2[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__18 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__2[5]));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__2[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__2[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__2[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__2[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__2[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__2[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[0]_i_1__7 
       (.I0(n8m_reg_0_63_0_6_n_0),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_0),
        .I4(n8m_reg_0_63_14_20_n_2),
        .I5(n6m_reg_0_63_14_20_n_2),
        .O(s1_3[0]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[1]_i_1__7 
       (.I0(n8m_reg_0_63_0_6_n_1),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_1),
        .I4(n8m_reg_0_63_14_20_n_3),
        .I5(n6m_reg_0_63_14_20_n_3),
        .O(s1_3[1]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[2]_i_1__7 
       (.I0(n8m_reg_0_63_0_6_n_2),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_2),
        .I4(n8m_reg_0_63_14_20_n_4),
        .I5(n6m_reg_0_63_14_20_n_4),
        .O(s1_3[2]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[3]_i_1__7 
       (.I0(n8m_reg_0_63_0_6_n_3),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_3),
        .I4(n8m_reg_0_63_14_20_n_5),
        .I5(n6m_reg_0_63_14_20_n_5),
        .O(s1_3[3]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[4]_i_1__7 
       (.I0(n8m_reg_0_63_0_6_n_4),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_4),
        .I4(n8m_reg_0_63_14_20_n_6),
        .I5(n6m_reg_0_63_14_20_n_6),
        .O(s1_3[4]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[5]_i_1__7 
       (.I0(n8m_reg_0_63_0_6_n_5),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_5),
        .I4(n8m_reg_0_63_21_27_n_0),
        .I5(n6m_reg_0_63_21_27_n_0),
        .O(s1_3[5]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[6]_i_1__7 
       (.I0(n8m_reg_0_63_0_6_n_6),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_6),
        .I4(n8m_reg_0_63_21_27_n_1),
        .I5(n6m_reg_0_63_21_27_n_1),
        .O(s1_3[6]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[7]_i_1__7 
       (.I0(n8m_reg_0_63_7_13_n_0),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_0),
        .I4(n8m_reg_0_63_21_27_n_2),
        .I5(n6m_reg_0_63_21_27_n_2),
        .O(s1_3[7]));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a[5]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s27/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_UNIQ_BASE_ n6m_reg_0_63_0_6
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_0_6_n_0),
        .DOB(n6m_reg_0_63_0_6_n_1),
        .DOC(n6m_reg_0_63_0_6_n_2),
        .DOD(n6m_reg_0_63_0_6_n_3),
        .DOE(n6m_reg_0_63_0_6_n_4),
        .DOF(n6m_reg_0_63_0_6_n_5),
        .DOG(n6m_reg_0_63_0_6_n_6),
        .DOH(NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s27/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39684 n6m_reg_0_63_14_20
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_14_20_n_0),
        .DOB(n6m_reg_0_63_14_20_n_1),
        .DOC(n6m_reg_0_63_14_20_n_2),
        .DOD(n6m_reg_0_63_14_20_n_3),
        .DOE(n6m_reg_0_63_14_20_n_4),
        .DOF(n6m_reg_0_63_14_20_n_5),
        .DOG(n6m_reg_0_63_14_20_n_6),
        .DOH(NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s27/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39685 n6m_reg_0_63_21_27
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_21_27_n_0),
        .DOB(n6m_reg_0_63_21_27_n_1),
        .DOC(n6m_reg_0_63_21_27_n_2),
        .DOD(n6m_reg_0_63_21_27_n_3),
        .DOE(n6m_reg_0_63_21_27_n_4),
        .DOF(n6m_reg_0_63_21_27_n_5),
        .DOG(n6m_reg_0_63_21_27_n_6),
        .DOH(NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s27/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39686 n6m_reg_0_63_28_31
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_28_31_n_0),
        .DOB(n6m_reg_0_63_28_31_n_1),
        .DOC(n6m_reg_0_63_28_31_n_2),
        .DOD(n6m_reg_0_63_28_31_n_3),
        .DOE(NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s27/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39687 n6m_reg_0_63_7_13
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_7_13_n_0),
        .DOB(n6m_reg_0_63_7_13_n_1),
        .DOC(n6m_reg_0_63_7_13_n_2),
        .DOD(n6m_reg_0_63_7_13_n_3),
        .DOE(n6m_reg_0_63_7_13_n_4),
        .DOF(n6m_reg_0_63_7_13_n_5),
        .DOG(n6m_reg_0_63_7_13_n_6),
        .DOH(NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s27/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39688 n8m_reg_0_63_0_6
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n8m_reg_0_63_0_6_n_0),
        .DOB(n8m_reg_0_63_0_6_n_1),
        .DOC(n8m_reg_0_63_0_6_n_2),
        .DOD(n8m_reg_0_63_0_6_n_3),
        .DOE(n8m_reg_0_63_0_6_n_4),
        .DOF(n8m_reg_0_63_0_6_n_5),
        .DOG(n8m_reg_0_63_0_6_n_6),
        .DOH(NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s27/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39689 n8m_reg_0_63_14_20
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n8m_reg_0_63_14_20_n_0),
        .DOB(n8m_reg_0_63_14_20_n_1),
        .DOC(n8m_reg_0_63_14_20_n_2),
        .DOD(n8m_reg_0_63_14_20_n_3),
        .DOE(n8m_reg_0_63_14_20_n_4),
        .DOF(n8m_reg_0_63_14_20_n_5),
        .DOG(n8m_reg_0_63_14_20_n_6),
        .DOH(NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s27/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39690 n8m_reg_0_63_21_27
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n8m_reg_0_63_21_27_n_0),
        .DOB(n8m_reg_0_63_21_27_n_1),
        .DOC(n8m_reg_0_63_21_27_n_2),
        .DOD(n8m_reg_0_63_21_27_n_3),
        .DOE(n8m_reg_0_63_21_27_n_4),
        .DOF(n8m_reg_0_63_21_27_n_5),
        .DOG(n8m_reg_0_63_21_27_n_6),
        .DOH(NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s27/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39691 n8m_reg_0_63_28_31
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n8m_reg_0_63_28_31_n_0),
        .DOB(n8m_reg_0_63_28_31_n_1),
        .DOC(n8m_reg_0_63_28_31_n_2),
        .DOD(n8m_reg_0_63_28_31_n_3),
        .DOE(NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s1/s27/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39692 n8m_reg_0_63_7_13
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n8m_reg_0_63_7_13_n_0),
        .DOB(n8m_reg_0_63_7_13_n_1),
        .DOC(n8m_reg_0_63_7_13_n_2),
        .DOD(n8m_reg_0_63_7_13_n_3),
        .DOE(n8m_reg_0_63_7_13_n_4),
        .DOF(n8m_reg_0_63_7_13_n_5),
        .DOG(n8m_reg_0_63_7_13_n_6),
        .DOH(NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(1'b1),
        .Q(\n9_reg[0]_0 ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_27" *) 
module switch_elements_cf_fft_512_8_27_3
   (\n9_reg[0]_0 ,
    s7_3,
    rst_i,
    enable_i,
    clk_i,
    i8,
    i1);
  output \n9_reg[0]_0 ;
  output [15:0]s7_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [0:0]i8;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [5:0]n2__1;
  wire [5:0]n3_reg;
  wire n6m_reg_0_63_0_6_n_0;
  wire n6m_reg_0_63_0_6_n_1;
  wire n6m_reg_0_63_0_6_n_2;
  wire n6m_reg_0_63_0_6_n_3;
  wire n6m_reg_0_63_0_6_n_4;
  wire n6m_reg_0_63_0_6_n_5;
  wire n6m_reg_0_63_0_6_n_6;
  wire n6m_reg_0_63_14_20_n_0;
  wire n6m_reg_0_63_14_20_n_1;
  wire n6m_reg_0_63_14_20_n_2;
  wire n6m_reg_0_63_14_20_n_3;
  wire n6m_reg_0_63_14_20_n_4;
  wire n6m_reg_0_63_14_20_n_5;
  wire n6m_reg_0_63_14_20_n_6;
  wire n6m_reg_0_63_21_27_n_0;
  wire n6m_reg_0_63_21_27_n_1;
  wire n6m_reg_0_63_21_27_n_2;
  wire n6m_reg_0_63_21_27_n_3;
  wire n6m_reg_0_63_21_27_n_4;
  wire n6m_reg_0_63_21_27_n_5;
  wire n6m_reg_0_63_21_27_n_6;
  wire n6m_reg_0_63_28_31_n_0;
  wire n6m_reg_0_63_28_31_n_1;
  wire n6m_reg_0_63_28_31_n_2;
  wire n6m_reg_0_63_28_31_n_3;
  wire n6m_reg_0_63_7_13_n_0;
  wire n6m_reg_0_63_7_13_n_1;
  wire n6m_reg_0_63_7_13_n_2;
  wire n6m_reg_0_63_7_13_n_3;
  wire n6m_reg_0_63_7_13_n_4;
  wire n6m_reg_0_63_7_13_n_5;
  wire n6m_reg_0_63_7_13_n_6;
  wire [31:0]n8;
  wire [5:0]n8a;
  wire [5:0]n8a__0;
  wire \n9_reg[0]_0 ;
  wire rst_i;
  wire [15:0]s7_3;
  wire NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED;

  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__0_i_1__4
       (.I0(n8[14]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_0),
        .I4(n8[30]),
        .I5(n6m_reg_0_63_28_31_n_2),
        .O(s7_3[14]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__1_i_1__4
       (.I0(n8[13]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_6),
        .I4(n8[29]),
        .I5(n6m_reg_0_63_28_31_n_1),
        .O(s7_3[13]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__2_i_1__4
       (.I0(n8[12]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_5),
        .I4(n8[28]),
        .I5(n6m_reg_0_63_28_31_n_0),
        .O(s7_3[12]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__3_i_1__4
       (.I0(n8[11]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_4),
        .I4(n8[27]),
        .I5(n6m_reg_0_63_21_27_n_6),
        .O(s7_3[11]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__4_i_1__4
       (.I0(n8[10]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_3),
        .I4(n8[26]),
        .I5(n6m_reg_0_63_21_27_n_5),
        .O(s7_3[10]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__5_i_1__4
       (.I0(n8[9]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_2),
        .I4(n8[25]),
        .I5(n6m_reg_0_63_21_27_n_4),
        .O(s7_3[9]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__6_i_1__4
       (.I0(n8[8]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_1),
        .I4(n8[24]),
        .I5(n6m_reg_0_63_21_27_n_3),
        .O(s7_3[8]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22_i_1__4
       (.I0(n8[15]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_1),
        .I4(n8[31]),
        .I5(n6m_reg_0_63_28_31_n_3),
        .O(s7_3[15]));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__12 
       (.I0(n3_reg[0]),
        .O(n2__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__12 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__1[1]));
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__12 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__1[2]));
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__12 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__1[3]));
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__12 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__1[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__12 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__1[5]));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[0]_i_1__4 
       (.I0(n8[0]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_0),
        .I4(n8[16]),
        .I5(n6m_reg_0_63_14_20_n_2),
        .O(s7_3[0]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[1]_i_1__4 
       (.I0(n8[1]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_1),
        .I4(n8[17]),
        .I5(n6m_reg_0_63_14_20_n_3),
        .O(s7_3[1]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[2]_i_1__4 
       (.I0(n8[2]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_2),
        .I4(n8[18]),
        .I5(n6m_reg_0_63_14_20_n_4),
        .O(s7_3[2]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[3]_i_1__4 
       (.I0(n8[3]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_3),
        .I4(n8[19]),
        .I5(n6m_reg_0_63_14_20_n_5),
        .O(s7_3[3]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[4]_i_1__4 
       (.I0(n8[4]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_4),
        .I4(n8[20]),
        .I5(n6m_reg_0_63_14_20_n_6),
        .O(s7_3[4]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[5]_i_1__4 
       (.I0(n8[5]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_5),
        .I4(n8[21]),
        .I5(n6m_reg_0_63_21_27_n_0),
        .O(s7_3[5]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[6]_i_1__4 
       (.I0(n8[6]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_6),
        .I4(n8[22]),
        .I5(n6m_reg_0_63_21_27_n_1),
        .O(s7_3[6]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[7]_i_1__4 
       (.I0(n8[7]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_0),
        .I4(n8[23]),
        .I5(n6m_reg_0_63_21_27_n_2),
        .O(s7_3[7]));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a[5]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39873 n6m_reg_0_63_0_6
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_0_6_n_0),
        .DOB(n6m_reg_0_63_0_6_n_1),
        .DOC(n6m_reg_0_63_0_6_n_2),
        .DOD(n6m_reg_0_63_0_6_n_3),
        .DOE(n6m_reg_0_63_0_6_n_4),
        .DOF(n6m_reg_0_63_0_6_n_5),
        .DOG(n6m_reg_0_63_0_6_n_6),
        .DOH(NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39874 n6m_reg_0_63_14_20
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_14_20_n_0),
        .DOB(n6m_reg_0_63_14_20_n_1),
        .DOC(n6m_reg_0_63_14_20_n_2),
        .DOD(n6m_reg_0_63_14_20_n_3),
        .DOE(n6m_reg_0_63_14_20_n_4),
        .DOF(n6m_reg_0_63_14_20_n_5),
        .DOG(n6m_reg_0_63_14_20_n_6),
        .DOH(NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39875 n6m_reg_0_63_21_27
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_21_27_n_0),
        .DOB(n6m_reg_0_63_21_27_n_1),
        .DOC(n6m_reg_0_63_21_27_n_2),
        .DOD(n6m_reg_0_63_21_27_n_3),
        .DOE(n6m_reg_0_63_21_27_n_4),
        .DOF(n6m_reg_0_63_21_27_n_5),
        .DOG(n6m_reg_0_63_21_27_n_6),
        .DOH(NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39876 n6m_reg_0_63_28_31
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_28_31_n_0),
        .DOB(n6m_reg_0_63_28_31_n_1),
        .DOC(n6m_reg_0_63_28_31_n_2),
        .DOD(n6m_reg_0_63_28_31_n_3),
        .DOE(NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39877 n6m_reg_0_63_7_13
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_7_13_n_0),
        .DOB(n6m_reg_0_63_7_13_n_1),
        .DOC(n6m_reg_0_63_7_13_n_2),
        .DOD(n6m_reg_0_63_7_13_n_3),
        .DOE(n6m_reg_0_63_7_13_n_4),
        .DOF(n6m_reg_0_63_7_13_n_5),
        .DOG(n6m_reg_0_63_7_13_n_6),
        .DOH(NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39878 n8m_reg_0_63_0_6
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n8[0]),
        .DOB(n8[1]),
        .DOC(n8[2]),
        .DOD(n8[3]),
        .DOE(n8[4]),
        .DOF(n8[5]),
        .DOG(n8[6]),
        .DOH(NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39879 n8m_reg_0_63_14_20
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n8[14]),
        .DOB(n8[15]),
        .DOC(n8[16]),
        .DOD(n8[17]),
        .DOE(n8[18]),
        .DOF(n8[19]),
        .DOG(n8[20]),
        .DOH(NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39880 n8m_reg_0_63_21_27
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n8[21]),
        .DOB(n8[22]),
        .DOC(n8[23]),
        .DOD(n8[24]),
        .DOE(n8[25]),
        .DOF(n8[26]),
        .DOG(n8[27]),
        .DOH(NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39881 n8m_reg_0_63_28_31
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n8[28]),
        .DOB(n8[29]),
        .DOC(n8[30]),
        .DOD(n8[31]),
        .DOE(NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39882 n8m_reg_0_63_7_13
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n8[7]),
        .DOB(n8[8]),
        .DOC(n8[9]),
        .DOD(n8[10]),
        .DOE(n8[11]),
        .DOF(n8[12]),
        .DOG(n8[13]),
        .DOH(NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(1'b1),
        .Q(\n9_reg[0]_0 ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_27" *) 
module switch_elements_cf_fft_512_8_27_6
   (\n9_reg[0]_0 ,
    s6_3,
    rst_i,
    enable_i,
    clk_i,
    i8,
    i1);
  output \n9_reg[0]_0 ;
  output [15:0]s6_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [0:0]i8;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [5:0]n2__1;
  wire [5:0]n3_reg;
  wire n6m_reg_0_63_0_6_n_0;
  wire n6m_reg_0_63_0_6_n_1;
  wire n6m_reg_0_63_0_6_n_2;
  wire n6m_reg_0_63_0_6_n_3;
  wire n6m_reg_0_63_0_6_n_4;
  wire n6m_reg_0_63_0_6_n_5;
  wire n6m_reg_0_63_0_6_n_6;
  wire n6m_reg_0_63_14_20_n_0;
  wire n6m_reg_0_63_14_20_n_1;
  wire n6m_reg_0_63_14_20_n_2;
  wire n6m_reg_0_63_14_20_n_3;
  wire n6m_reg_0_63_14_20_n_4;
  wire n6m_reg_0_63_14_20_n_5;
  wire n6m_reg_0_63_14_20_n_6;
  wire n6m_reg_0_63_21_27_n_0;
  wire n6m_reg_0_63_21_27_n_1;
  wire n6m_reg_0_63_21_27_n_2;
  wire n6m_reg_0_63_21_27_n_3;
  wire n6m_reg_0_63_21_27_n_4;
  wire n6m_reg_0_63_21_27_n_5;
  wire n6m_reg_0_63_21_27_n_6;
  wire n6m_reg_0_63_28_31_n_0;
  wire n6m_reg_0_63_28_31_n_1;
  wire n6m_reg_0_63_28_31_n_2;
  wire n6m_reg_0_63_28_31_n_3;
  wire n6m_reg_0_63_7_13_n_0;
  wire n6m_reg_0_63_7_13_n_1;
  wire n6m_reg_0_63_7_13_n_2;
  wire n6m_reg_0_63_7_13_n_3;
  wire n6m_reg_0_63_7_13_n_4;
  wire n6m_reg_0_63_7_13_n_5;
  wire n6m_reg_0_63_7_13_n_6;
  wire [31:0]n8;
  wire [5:0]n8a;
  wire [5:0]n8a__0;
  wire \n9_reg[0]_0 ;
  wire rst_i;
  wire [15:0]s6_3;
  wire NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED;

  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__0_i_1__3
       (.I0(n8[14]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_0),
        .I4(n8[30]),
        .I5(n6m_reg_0_63_28_31_n_2),
        .O(s6_3[14]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__1_i_1__3
       (.I0(n8[13]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_6),
        .I4(n8[29]),
        .I5(n6m_reg_0_63_28_31_n_1),
        .O(s6_3[13]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__2_i_1__3
       (.I0(n8[12]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_5),
        .I4(n8[28]),
        .I5(n6m_reg_0_63_28_31_n_0),
        .O(s6_3[12]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__3_i_1__3
       (.I0(n8[11]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_4),
        .I4(n8[27]),
        .I5(n6m_reg_0_63_21_27_n_6),
        .O(s6_3[11]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__4_i_1__3
       (.I0(n8[10]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_3),
        .I4(n8[26]),
        .I5(n6m_reg_0_63_21_27_n_5),
        .O(s6_3[10]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__5_i_1__3
       (.I0(n8[9]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_2),
        .I4(n8[25]),
        .I5(n6m_reg_0_63_21_27_n_4),
        .O(s6_3[9]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__6_i_1__3
       (.I0(n8[8]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_1),
        .I4(n8[24]),
        .I5(n6m_reg_0_63_21_27_n_3),
        .O(s6_3[8]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22_i_1__3
       (.I0(n8[15]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_1),
        .I4(n8[31]),
        .I5(n6m_reg_0_63_28_31_n_3),
        .O(s6_3[15]));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__10 
       (.I0(n3_reg[0]),
        .O(n2__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__10 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__1[1]));
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__10 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__1[2]));
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__10 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__1[3]));
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__10 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__1[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__10 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__1[5]));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[0]_i_1__3 
       (.I0(n8[0]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_0),
        .I4(n8[16]),
        .I5(n6m_reg_0_63_14_20_n_2),
        .O(s6_3[0]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[1]_i_1__3 
       (.I0(n8[1]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_1),
        .I4(n8[17]),
        .I5(n6m_reg_0_63_14_20_n_3),
        .O(s6_3[1]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[2]_i_1__3 
       (.I0(n8[2]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_2),
        .I4(n8[18]),
        .I5(n6m_reg_0_63_14_20_n_4),
        .O(s6_3[2]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[3]_i_1__3 
       (.I0(n8[3]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_3),
        .I4(n8[19]),
        .I5(n6m_reg_0_63_14_20_n_5),
        .O(s6_3[3]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[4]_i_1__3 
       (.I0(n8[4]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_4),
        .I4(n8[20]),
        .I5(n6m_reg_0_63_14_20_n_6),
        .O(s6_3[4]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[5]_i_1__3 
       (.I0(n8[5]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_5),
        .I4(n8[21]),
        .I5(n6m_reg_0_63_21_27_n_0),
        .O(s6_3[5]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[6]_i_1__3 
       (.I0(n8[6]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_6),
        .I4(n8[22]),
        .I5(n6m_reg_0_63_21_27_n_1),
        .O(s6_3[6]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[7]_i_1__3 
       (.I0(n8[7]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_0),
        .I4(n8[23]),
        .I5(n6m_reg_0_63_21_27_n_2),
        .O(s6_3[7]));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a[5]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39848 n6m_reg_0_63_0_6
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_0_6_n_0),
        .DOB(n6m_reg_0_63_0_6_n_1),
        .DOC(n6m_reg_0_63_0_6_n_2),
        .DOD(n6m_reg_0_63_0_6_n_3),
        .DOE(n6m_reg_0_63_0_6_n_4),
        .DOF(n6m_reg_0_63_0_6_n_5),
        .DOG(n6m_reg_0_63_0_6_n_6),
        .DOH(NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39849 n6m_reg_0_63_14_20
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_14_20_n_0),
        .DOB(n6m_reg_0_63_14_20_n_1),
        .DOC(n6m_reg_0_63_14_20_n_2),
        .DOD(n6m_reg_0_63_14_20_n_3),
        .DOE(n6m_reg_0_63_14_20_n_4),
        .DOF(n6m_reg_0_63_14_20_n_5),
        .DOG(n6m_reg_0_63_14_20_n_6),
        .DOH(NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39850 n6m_reg_0_63_21_27
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_21_27_n_0),
        .DOB(n6m_reg_0_63_21_27_n_1),
        .DOC(n6m_reg_0_63_21_27_n_2),
        .DOD(n6m_reg_0_63_21_27_n_3),
        .DOE(n6m_reg_0_63_21_27_n_4),
        .DOF(n6m_reg_0_63_21_27_n_5),
        .DOG(n6m_reg_0_63_21_27_n_6),
        .DOH(NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39851 n6m_reg_0_63_28_31
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_28_31_n_0),
        .DOB(n6m_reg_0_63_28_31_n_1),
        .DOC(n6m_reg_0_63_28_31_n_2),
        .DOD(n6m_reg_0_63_28_31_n_3),
        .DOE(NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39852 n6m_reg_0_63_7_13
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_7_13_n_0),
        .DOB(n6m_reg_0_63_7_13_n_1),
        .DOC(n6m_reg_0_63_7_13_n_2),
        .DOD(n6m_reg_0_63_7_13_n_3),
        .DOE(n6m_reg_0_63_7_13_n_4),
        .DOF(n6m_reg_0_63_7_13_n_5),
        .DOG(n6m_reg_0_63_7_13_n_6),
        .DOH(NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39853 n8m_reg_0_63_0_6
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n8[0]),
        .DOB(n8[1]),
        .DOC(n8[2]),
        .DOD(n8[3]),
        .DOE(n8[4]),
        .DOF(n8[5]),
        .DOG(n8[6]),
        .DOH(NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39854 n8m_reg_0_63_14_20
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n8[14]),
        .DOB(n8[15]),
        .DOC(n8[16]),
        .DOD(n8[17]),
        .DOE(n8[18]),
        .DOF(n8[19]),
        .DOG(n8[20]),
        .DOH(NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39855 n8m_reg_0_63_21_27
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n8[21]),
        .DOB(n8[22]),
        .DOC(n8[23]),
        .DOD(n8[24]),
        .DOE(n8[25]),
        .DOF(n8[26]),
        .DOG(n8[27]),
        .DOH(NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39856 n8m_reg_0_63_28_31
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n8[28]),
        .DOB(n8[29]),
        .DOC(n8[30]),
        .DOD(n8[31]),
        .DOE(NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39857 n8m_reg_0_63_7_13
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n8[7]),
        .DOB(n8[8]),
        .DOC(n8[9]),
        .DOD(n8[10]),
        .DOE(n8[11]),
        .DOF(n8[12]),
        .DOG(n8[13]),
        .DOH(NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(1'b1),
        .Q(\n9_reg[0]_0 ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_27" *) 
module switch_elements_cf_fft_512_8_27_9
   (\n9_reg[0]_0 ,
    s5_3,
    rst_i,
    enable_i,
    clk_i,
    i8,
    i1);
  output \n9_reg[0]_0 ;
  output [15:0]s5_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [0:0]i8;
  input [29:0]i1;

  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [0:0]i8;
  wire [5:0]n2__1;
  wire [5:0]n3_reg;
  wire n6m_reg_0_63_0_6_n_0;
  wire n6m_reg_0_63_0_6_n_1;
  wire n6m_reg_0_63_0_6_n_2;
  wire n6m_reg_0_63_0_6_n_3;
  wire n6m_reg_0_63_0_6_n_4;
  wire n6m_reg_0_63_0_6_n_5;
  wire n6m_reg_0_63_0_6_n_6;
  wire n6m_reg_0_63_14_20_n_0;
  wire n6m_reg_0_63_14_20_n_1;
  wire n6m_reg_0_63_14_20_n_2;
  wire n6m_reg_0_63_14_20_n_3;
  wire n6m_reg_0_63_14_20_n_4;
  wire n6m_reg_0_63_14_20_n_5;
  wire n6m_reg_0_63_14_20_n_6;
  wire n6m_reg_0_63_21_27_n_0;
  wire n6m_reg_0_63_21_27_n_1;
  wire n6m_reg_0_63_21_27_n_2;
  wire n6m_reg_0_63_21_27_n_3;
  wire n6m_reg_0_63_21_27_n_4;
  wire n6m_reg_0_63_21_27_n_5;
  wire n6m_reg_0_63_21_27_n_6;
  wire n6m_reg_0_63_28_31_n_0;
  wire n6m_reg_0_63_28_31_n_1;
  wire n6m_reg_0_63_28_31_n_2;
  wire n6m_reg_0_63_28_31_n_3;
  wire n6m_reg_0_63_7_13_n_0;
  wire n6m_reg_0_63_7_13_n_1;
  wire n6m_reg_0_63_7_13_n_2;
  wire n6m_reg_0_63_7_13_n_3;
  wire n6m_reg_0_63_7_13_n_4;
  wire n6m_reg_0_63_7_13_n_5;
  wire n6m_reg_0_63_7_13_n_6;
  wire [31:0]n8;
  wire [5:0]n8a;
  wire [5:0]n8a__0;
  wire \n9_reg[0]_0 ;
  wire rst_i;
  wire [15:0]s5_3;
  wire NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED;

  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__0_i_1__2
       (.I0(n8[14]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_0),
        .I4(n8[30]),
        .I5(n6m_reg_0_63_28_31_n_2),
        .O(s5_3[14]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__1_i_1__2
       (.I0(n8[13]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_6),
        .I4(n8[29]),
        .I5(n6m_reg_0_63_28_31_n_1),
        .O(s5_3[13]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__2_i_1__2
       (.I0(n8[12]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_5),
        .I4(n8[28]),
        .I5(n6m_reg_0_63_28_31_n_0),
        .O(s5_3[12]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__3_i_1__2
       (.I0(n8[11]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_4),
        .I4(n8[27]),
        .I5(n6m_reg_0_63_21_27_n_6),
        .O(s5_3[11]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__4_i_1__2
       (.I0(n8[10]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_3),
        .I4(n8[26]),
        .I5(n6m_reg_0_63_21_27_n_5),
        .O(s5_3[10]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__5_i_1__2
       (.I0(n8[9]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_2),
        .I4(n8[25]),
        .I5(n6m_reg_0_63_21_27_n_4),
        .O(s5_3[9]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22__6_i_1__2
       (.I0(n8[8]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_1),
        .I4(n8[24]),
        .I5(n6m_reg_0_63_21_27_n_3),
        .O(s5_3[8]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    n22_i_1__2
       (.I0(n8[15]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_14_20_n_1),
        .I4(n8[31]),
        .I5(n6m_reg_0_63_28_31_n_3),
        .O(s5_3[15]));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__8 
       (.I0(n3_reg[0]),
        .O(n2__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__8 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__1[1]));
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__8 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__1[2]));
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__8 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__1[3]));
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__8 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__1[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__8 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__1[5]));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[0]_i_1__2 
       (.I0(n8[0]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_0),
        .I4(n8[16]),
        .I5(n6m_reg_0_63_14_20_n_2),
        .O(s5_3[0]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[1]_i_1__2 
       (.I0(n8[1]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_1),
        .I4(n8[17]),
        .I5(n6m_reg_0_63_14_20_n_3),
        .O(s5_3[1]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[2]_i_1__2 
       (.I0(n8[2]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_2),
        .I4(n8[18]),
        .I5(n6m_reg_0_63_14_20_n_4),
        .O(s5_3[2]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[3]_i_1__2 
       (.I0(n8[3]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_3),
        .I4(n8[19]),
        .I5(n6m_reg_0_63_14_20_n_5),
        .O(s5_3[3]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[4]_i_1__2 
       (.I0(n8[4]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_4),
        .I4(n8[20]),
        .I5(n6m_reg_0_63_14_20_n_6),
        .O(s5_3[4]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[5]_i_1__2 
       (.I0(n8[5]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_5),
        .I4(n8[21]),
        .I5(n6m_reg_0_63_21_27_n_0),
        .O(s5_3[5]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[6]_i_1__2 
       (.I0(n8[6]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_0_6_n_6),
        .I4(n8[22]),
        .I5(n6m_reg_0_63_21_27_n_1),
        .O(s5_3[6]));
  LUT6 #(
    .INIT(64'hBF8FB383BC8CB080)) 
    \n4[7]_i_1__2 
       (.I0(n8[7]),
        .I1(\n9_reg[0]_0 ),
        .I2(i8),
        .I3(n6m_reg_0_63_7_13_n_0),
        .I4(n8[23]),
        .I5(n6m_reg_0_63_21_27_n_2),
        .O(s5_3[7]));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a__0[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a__0[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a__0[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a__0[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a__0[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a__0[5]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a[0]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a[1]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a[2]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a[3]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a[4]),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a[5]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39823 n6m_reg_0_63_0_6
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_0_6_n_0),
        .DOB(n6m_reg_0_63_0_6_n_1),
        .DOC(n6m_reg_0_63_0_6_n_2),
        .DOD(n6m_reg_0_63_0_6_n_3),
        .DOE(n6m_reg_0_63_0_6_n_4),
        .DOF(n6m_reg_0_63_0_6_n_5),
        .DOG(n6m_reg_0_63_0_6_n_6),
        .DOH(NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39824 n6m_reg_0_63_14_20
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_14_20_n_0),
        .DOB(n6m_reg_0_63_14_20_n_1),
        .DOC(n6m_reg_0_63_14_20_n_2),
        .DOD(n6m_reg_0_63_14_20_n_3),
        .DOE(n6m_reg_0_63_14_20_n_4),
        .DOF(n6m_reg_0_63_14_20_n_5),
        .DOG(n6m_reg_0_63_14_20_n_6),
        .DOH(NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39825 n6m_reg_0_63_21_27
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_21_27_n_0),
        .DOB(n6m_reg_0_63_21_27_n_1),
        .DOC(n6m_reg_0_63_21_27_n_2),
        .DOD(n6m_reg_0_63_21_27_n_3),
        .DOE(n6m_reg_0_63_21_27_n_4),
        .DOF(n6m_reg_0_63_21_27_n_5),
        .DOG(n6m_reg_0_63_21_27_n_6),
        .DOH(NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39826 n6m_reg_0_63_28_31
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_28_31_n_0),
        .DOB(n6m_reg_0_63_28_31_n_1),
        .DOC(n6m_reg_0_63_28_31_n_2),
        .DOD(n6m_reg_0_63_28_31_n_3),
        .DOE(NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39827 n6m_reg_0_63_7_13
       (.ADDRA(n8a),
        .ADDRB(n8a),
        .ADDRC(n8a),
        .ADDRD(n8a),
        .ADDRE(n8a),
        .ADDRF(n8a),
        .ADDRG(n8a),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_7_13_n_0),
        .DOB(n6m_reg_0_63_7_13_n_1),
        .DOC(n6m_reg_0_63_7_13_n_2),
        .DOD(n6m_reg_0_63_7_13_n_3),
        .DOE(n6m_reg_0_63_7_13_n_4),
        .DOF(n6m_reg_0_63_7_13_n_5),
        .DOG(n6m_reg_0_63_7_13_n_6),
        .DOH(NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39828 n8m_reg_0_63_0_6
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[15]),
        .DIB(i1[0]),
        .DIC(i1[1]),
        .DID(i1[2]),
        .DIE(i1[3]),
        .DIF(i1[4]),
        .DIG(i1[5]),
        .DIH(1'b0),
        .DOA(n8[0]),
        .DOB(n8[1]),
        .DOC(n8[2]),
        .DOD(n8[3]),
        .DOE(n8[4]),
        .DOF(n8[5]),
        .DOG(n8[6]),
        .DOH(NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39829 n8m_reg_0_63_14_20
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[13]),
        .DIB(i1[14]),
        .DIC(i1[15]),
        .DID(i1[16]),
        .DIE(i1[17]),
        .DIF(i1[18]),
        .DIG(i1[19]),
        .DIH(1'b0),
        .DOA(n8[14]),
        .DOB(n8[15]),
        .DOC(n8[16]),
        .DOD(n8[17]),
        .DOE(n8[18]),
        .DOF(n8[19]),
        .DOG(n8[20]),
        .DOH(NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39830 n8m_reg_0_63_21_27
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[20]),
        .DIB(i1[21]),
        .DIC(i1[22]),
        .DID(i1[7]),
        .DIE(i1[23]),
        .DIF(i1[24]),
        .DIG(i1[25]),
        .DIH(1'b0),
        .DOA(n8[21]),
        .DOB(n8[22]),
        .DOC(n8[23]),
        .DOD(n8[24]),
        .DOE(n8[25]),
        .DOF(n8[26]),
        .DOG(n8[27]),
        .DOH(NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39831 n8m_reg_0_63_28_31
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[26]),
        .DIB(i1[27]),
        .DIC(i1[28]),
        .DID(i1[29]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n8[28]),
        .DOB(n8[29]),
        .DOC(n8[30]),
        .DOD(n8[31]),
        .DOE(NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "s29/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39832 n8m_reg_0_63_7_13
       (.ADDRA(n8a__0),
        .ADDRB(n8a__0),
        .ADDRC(n8a__0),
        .ADDRD(n8a__0),
        .ADDRE(n8a__0),
        .ADDRF(n8a__0),
        .ADDRG(n8a__0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i1[6]),
        .DIB(i1[7]),
        .DIC(i1[8]),
        .DID(i1[9]),
        .DIE(i1[10]),
        .DIF(i1[11]),
        .DIG(i1[12]),
        .DIH(1'b0),
        .DOA(n8[7]),
        .DOB(n8[8]),
        .DOC(n8[9]),
        .DOD(n8[10]),
        .DOE(n8[11]),
        .DOF(n8[12]),
        .DOG(n8[13]),
        .DOH(NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(1'b1),
        .Q(\n9_reg[0]_0 ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_3" *) 
module switch_elements_cf_fft_512_8_3
   (\n5_reg[0] ,
    n4,
    clk_i,
    i2,
    i8,
    \n1_reg[15] ,
    enable_i,
    rst_i);
  output [15:0]\n5_reg[0] ;
  output n4;
  input clk_i;
  input [31:0]i2;
  input [0:0]i8;
  input \n1_reg[15] ;
  input [0:0]enable_i;
  input rst_i;

  wire clk_i;
  wire [0:0]enable_i;
  wire [31:0]i2;
  wire [0:0]i8;
  wire [31:0]n11;
  wire [6:0]n11a_1;
  wire \n1_reg[15] ;
  wire [6:0]n2__1;
  wire \n3[6]_i_2__8_n_0 ;
  wire [6:0]n3_reg;
  wire n4;
  wire \n5[0]_i_2__8_n_0 ;
  wire [15:0]\n5_reg[0] ;
  wire \n9a_reg_n_0_[0] ;
  wire \n9a_reg_n_0_[1] ;
  wire \n9a_reg_n_0_[2] ;
  wire \n9a_reg_n_0_[3] ;
  wire \n9a_reg_n_0_[4] ;
  wire \n9a_reg_n_0_[5] ;
  wire n9m_reg_0_63_0_6_n_0;
  wire n9m_reg_0_63_0_6_n_1;
  wire n9m_reg_0_63_0_6_n_2;
  wire n9m_reg_0_63_0_6_n_3;
  wire n9m_reg_0_63_0_6_n_4;
  wire n9m_reg_0_63_0_6_n_5;
  wire n9m_reg_0_63_0_6_n_6;
  wire n9m_reg_0_63_14_20_n_0;
  wire n9m_reg_0_63_14_20_n_1;
  wire n9m_reg_0_63_14_20_n_2;
  wire n9m_reg_0_63_14_20_n_3;
  wire n9m_reg_0_63_14_20_n_4;
  wire n9m_reg_0_63_14_20_n_5;
  wire n9m_reg_0_63_14_20_n_6;
  wire n9m_reg_0_63_21_27_n_0;
  wire n9m_reg_0_63_21_27_n_1;
  wire n9m_reg_0_63_21_27_n_2;
  wire n9m_reg_0_63_21_27_n_3;
  wire n9m_reg_0_63_21_27_n_4;
  wire n9m_reg_0_63_21_27_n_5;
  wire n9m_reg_0_63_21_27_n_6;
  wire n9m_reg_0_63_28_31_n_0;
  wire n9m_reg_0_63_28_31_n_1;
  wire n9m_reg_0_63_28_31_n_2;
  wire n9m_reg_0_63_28_31_n_3;
  wire n9m_reg_0_63_7_13_n_0;
  wire n9m_reg_0_63_7_13_n_1;
  wire n9m_reg_0_63_7_13_n_2;
  wire n9m_reg_0_63_7_13_n_3;
  wire n9m_reg_0_63_7_13_n_4;
  wire n9m_reg_0_63_7_13_n_5;
  wire n9m_reg_0_63_7_13_n_6;
  wire n9m_reg_64_127_0_6_n_0;
  wire n9m_reg_64_127_0_6_n_1;
  wire n9m_reg_64_127_0_6_n_2;
  wire n9m_reg_64_127_0_6_n_3;
  wire n9m_reg_64_127_0_6_n_4;
  wire n9m_reg_64_127_0_6_n_5;
  wire n9m_reg_64_127_0_6_n_6;
  wire n9m_reg_64_127_14_20_n_0;
  wire n9m_reg_64_127_14_20_n_1;
  wire n9m_reg_64_127_14_20_n_2;
  wire n9m_reg_64_127_14_20_n_3;
  wire n9m_reg_64_127_14_20_n_4;
  wire n9m_reg_64_127_14_20_n_5;
  wire n9m_reg_64_127_14_20_n_6;
  wire n9m_reg_64_127_21_27_n_0;
  wire n9m_reg_64_127_21_27_n_1;
  wire n9m_reg_64_127_21_27_n_2;
  wire n9m_reg_64_127_21_27_n_3;
  wire n9m_reg_64_127_21_27_n_4;
  wire n9m_reg_64_127_21_27_n_5;
  wire n9m_reg_64_127_21_27_n_6;
  wire n9m_reg_64_127_28_31_n_0;
  wire n9m_reg_64_127_28_31_n_1;
  wire n9m_reg_64_127_28_31_n_2;
  wire n9m_reg_64_127_28_31_n_3;
  wire n9m_reg_64_127_7_13_n_0;
  wire n9m_reg_64_127_7_13_n_1;
  wire n9m_reg_64_127_7_13_n_2;
  wire n9m_reg_64_127_7_13_n_3;
  wire n9m_reg_64_127_7_13_n_4;
  wire n9m_reg_64_127_7_13_n_5;
  wire n9m_reg_64_127_7_13_n_6;
  wire [31:0]p_0_in;
  wire rst_i;
  wire NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED;
  wire NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED;
  wire NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED;

  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39918 n11m_reg_0_63_0_6
       (.ADDRA({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRB({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRC({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRD({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRE({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRF({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRG({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[0]),
        .DIB(i2[1]),
        .DIC(i2[2]),
        .DID(i2[3]),
        .DIE(i2[4]),
        .DIF(i2[5]),
        .DIG(i2[6]),
        .DIH(1'b0),
        .DOA(n11[0]),
        .DOB(n11[1]),
        .DOC(n11[2]),
        .DOD(n11[3]),
        .DOE(n11[4]),
        .DOF(n11[5]),
        .DOG(n11[6]),
        .DOH(NLW_n11m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39919 n11m_reg_0_63_14_20
       (.ADDRA({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRB({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRC({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRD({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRE({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRF({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRG({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[14]),
        .DIB(i2[15]),
        .DIC(i2[16]),
        .DID(i2[17]),
        .DIE(i2[18]),
        .DIF(i2[19]),
        .DIG(i2[20]),
        .DIH(1'b0),
        .DOA(n11[14]),
        .DOB(n11[15]),
        .DOC(n11[16]),
        .DOD(n11[17]),
        .DOE(n11[18]),
        .DOF(n11[19]),
        .DOG(n11[20]),
        .DOH(NLW_n11m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39920 n11m_reg_0_63_21_27
       (.ADDRA({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRB({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRC({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRD({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRE({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRF({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRG({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[21]),
        .DIB(i2[22]),
        .DIC(i2[23]),
        .DID(i2[24]),
        .DIE(i2[25]),
        .DIF(i2[26]),
        .DIG(i2[27]),
        .DIH(1'b0),
        .DOA(n11[21]),
        .DOB(n11[22]),
        .DOC(n11[23]),
        .DOD(n11[24]),
        .DOE(n11[25]),
        .DOF(n11[26]),
        .DOG(n11[27]),
        .DOH(NLW_n11m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39921 n11m_reg_0_63_28_31
       (.ADDRA({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRB({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRC({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRD({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRE({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRF({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRG({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[28]),
        .DIB(i2[29]),
        .DIC(i2[30]),
        .DID(i2[31]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n11[28]),
        .DOB(n11[29]),
        .DOC(n11[30]),
        .DOD(n11[31]),
        .DOE(NLW_n11m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n11m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n11m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n11m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n11m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39922 n11m_reg_0_63_7_13
       (.ADDRA({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRB({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRC({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRD({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRE({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRF({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRG({\n9a_reg_n_0_[5] ,\n9a_reg_n_0_[4] ,\n9a_reg_n_0_[3] ,\n9a_reg_n_0_[2] ,\n9a_reg_n_0_[1] ,\n9a_reg_n_0_[0] }),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[7]),
        .DIB(i2[8]),
        .DIC(i2[9]),
        .DID(i2[10]),
        .DIE(i2[11]),
        .DIF(i2[12]),
        .DIG(i2[13]),
        .DIH(1'b0),
        .DOA(n11[7]),
        .DOB(n11[8]),
        .DOC(n11[9]),
        .DOD(n11[10]),
        .DOE(n11[11]),
        .DOF(n11[12]),
        .DOG(n11[13]),
        .DOH(NLW_n11m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[0]_i_2__6 
       (.I0(n11[16]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_14_20_n_2),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_14_20_n_2),
        .O(p_0_in[16]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[0]_i_3__6 
       (.I0(n11[0]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_0_6_n_0),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_0_6_n_0),
        .O(p_0_in[0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[10]_i_2__6 
       (.I0(n11[26]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_21_27_n_5),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_21_27_n_5),
        .O(p_0_in[26]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[10]_i_3__6 
       (.I0(n11[10]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_7_13_n_3),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_7_13_n_3),
        .O(p_0_in[10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[11]_i_2__6 
       (.I0(n11[27]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_21_27_n_6),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_21_27_n_6),
        .O(p_0_in[27]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[11]_i_3__6 
       (.I0(n11[11]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_7_13_n_4),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_7_13_n_4),
        .O(p_0_in[11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[12]_i_2__6 
       (.I0(n11[28]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_28_31_n_0),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_28_31_n_0),
        .O(p_0_in[28]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[12]_i_3__6 
       (.I0(n11[12]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_7_13_n_5),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_7_13_n_5),
        .O(p_0_in[12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[13]_i_2__6 
       (.I0(n11[29]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_28_31_n_1),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_28_31_n_1),
        .O(p_0_in[29]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[13]_i_3__6 
       (.I0(n11[13]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_7_13_n_6),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_7_13_n_6),
        .O(p_0_in[13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[14]_i_2__6 
       (.I0(n11[30]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_28_31_n_2),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_28_31_n_2),
        .O(p_0_in[30]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[14]_i_3__6 
       (.I0(n11[14]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_14_20_n_0),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_14_20_n_0),
        .O(p_0_in[14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[15]_i_2__6 
       (.I0(n11[31]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_28_31_n_3),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_28_31_n_3),
        .O(p_0_in[31]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[15]_i_3__6 
       (.I0(n11[15]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_14_20_n_1),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_14_20_n_1),
        .O(p_0_in[15]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[1]_i_2__6 
       (.I0(n11[17]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_14_20_n_3),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_14_20_n_3),
        .O(p_0_in[17]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[1]_i_3__6 
       (.I0(n11[1]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_0_6_n_1),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_0_6_n_1),
        .O(p_0_in[1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[2]_i_2__6 
       (.I0(n11[18]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_14_20_n_4),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_14_20_n_4),
        .O(p_0_in[18]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[2]_i_3__6 
       (.I0(n11[2]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_0_6_n_2),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_0_6_n_2),
        .O(p_0_in[2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[3]_i_2__6 
       (.I0(n11[19]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_14_20_n_5),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_14_20_n_5),
        .O(p_0_in[19]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[3]_i_3__6 
       (.I0(n11[3]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_0_6_n_3),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_0_6_n_3),
        .O(p_0_in[3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[4]_i_2__6 
       (.I0(n11[20]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_14_20_n_6),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_14_20_n_6),
        .O(p_0_in[20]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[4]_i_3__6 
       (.I0(n11[4]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_0_6_n_4),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_0_6_n_4),
        .O(p_0_in[4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[5]_i_2__6 
       (.I0(n11[21]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_21_27_n_0),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_21_27_n_0),
        .O(p_0_in[21]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[5]_i_3__6 
       (.I0(n11[5]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_0_6_n_5),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_0_6_n_5),
        .O(p_0_in[5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[6]_i_2__6 
       (.I0(n11[22]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_21_27_n_1),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_21_27_n_1),
        .O(p_0_in[22]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[6]_i_3__6 
       (.I0(n11[6]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_0_6_n_6),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_0_6_n_6),
        .O(p_0_in[6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[7]_i_2__6 
       (.I0(n11[23]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_21_27_n_2),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_21_27_n_2),
        .O(p_0_in[23]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[7]_i_3__6 
       (.I0(n11[7]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_7_13_n_0),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_7_13_n_0),
        .O(p_0_in[7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[8]_i_2__6 
       (.I0(n11[24]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_21_27_n_3),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_21_27_n_3),
        .O(p_0_in[24]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[8]_i_3__6 
       (.I0(n11[8]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_7_13_n_1),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_7_13_n_1),
        .O(p_0_in[8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[9]_i_2__6 
       (.I0(n11[25]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_21_27_n_4),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_21_27_n_4),
        .O(p_0_in[25]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \n1[9]_i_3__6 
       (.I0(n11[9]),
        .I1(\n1_reg[15] ),
        .I2(n9m_reg_64_127_7_13_n_2),
        .I3(n11a_1[6]),
        .I4(n9m_reg_0_63_7_13_n_2),
        .O(p_0_in[9]));
  MUXF7 \n1_reg[0]_i_1 
       (.I0(p_0_in[16]),
        .I1(p_0_in[0]),
        .O(\n5_reg[0] [0]),
        .S(i8));
  MUXF7 \n1_reg[10]_i_1 
       (.I0(p_0_in[26]),
        .I1(p_0_in[10]),
        .O(\n5_reg[0] [10]),
        .S(i8));
  MUXF7 \n1_reg[11]_i_1 
       (.I0(p_0_in[27]),
        .I1(p_0_in[11]),
        .O(\n5_reg[0] [11]),
        .S(i8));
  MUXF7 \n1_reg[12]_i_1 
       (.I0(p_0_in[28]),
        .I1(p_0_in[12]),
        .O(\n5_reg[0] [12]),
        .S(i8));
  MUXF7 \n1_reg[13]_i_1 
       (.I0(p_0_in[29]),
        .I1(p_0_in[13]),
        .O(\n5_reg[0] [13]),
        .S(i8));
  MUXF7 \n1_reg[14]_i_1 
       (.I0(p_0_in[30]),
        .I1(p_0_in[14]),
        .O(\n5_reg[0] [14]),
        .S(i8));
  MUXF7 \n1_reg[15]_i_1 
       (.I0(p_0_in[31]),
        .I1(p_0_in[15]),
        .O(\n5_reg[0] [15]),
        .S(i8));
  MUXF7 \n1_reg[1]_i_1 
       (.I0(p_0_in[17]),
        .I1(p_0_in[1]),
        .O(\n5_reg[0] [1]),
        .S(i8));
  MUXF7 \n1_reg[2]_i_1 
       (.I0(p_0_in[18]),
        .I1(p_0_in[2]),
        .O(\n5_reg[0] [2]),
        .S(i8));
  MUXF7 \n1_reg[3]_i_1 
       (.I0(p_0_in[19]),
        .I1(p_0_in[3]),
        .O(\n5_reg[0] [3]),
        .S(i8));
  MUXF7 \n1_reg[4]_i_1 
       (.I0(p_0_in[20]),
        .I1(p_0_in[4]),
        .O(\n5_reg[0] [4]),
        .S(i8));
  MUXF7 \n1_reg[5]_i_1 
       (.I0(p_0_in[21]),
        .I1(p_0_in[5]),
        .O(\n5_reg[0] [5]),
        .S(i8));
  MUXF7 \n1_reg[6]_i_1 
       (.I0(p_0_in[22]),
        .I1(p_0_in[6]),
        .O(\n5_reg[0] [6]),
        .S(i8));
  MUXF7 \n1_reg[7]_i_1 
       (.I0(p_0_in[23]),
        .I1(p_0_in[7]),
        .O(\n5_reg[0] [7]),
        .S(i8));
  MUXF7 \n1_reg[8]_i_1 
       (.I0(p_0_in[24]),
        .I1(p_0_in[8]),
        .O(\n5_reg[0] [8]),
        .S(i8));
  MUXF7 \n1_reg[9]_i_1 
       (.I0(p_0_in[25]),
        .I1(p_0_in[9]),
        .O(\n5_reg[0] [9]),
        .S(i8));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__17 
       (.I0(n3_reg[0]),
        .O(n2__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair235" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__17 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__1[1]));
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__17 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__1[2]));
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__17 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__1[3]));
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__17 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__1[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__17 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__1[5]));
  LUT3 #(
    .INIT(8'hD2)) 
    \n3[6]_i_1__8 
       (.I0(n3_reg[5]),
        .I1(\n3[6]_i_2__8_n_0 ),
        .I2(n3_reg[6]),
        .O(n2__1[6]));
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \n3[6]_i_2__8 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(\n3[6]_i_2__8_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__1[6]),
        .Q(n3_reg[6]),
        .R(rst_i));
  (* SOFT_HLUTNM = "soft_lutpair235" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \n5[0]_i_1__8 
       (.I0(n3_reg[0]),
        .I1(\n5[0]_i_2__8_n_0 ),
        .I2(i8),
        .O(n4));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \n5[0]_i_2__8 
       (.I0(n3_reg[3]),
        .I1(n3_reg[4]),
        .I2(n3_reg[1]),
        .I3(n3_reg[2]),
        .I4(n3_reg[6]),
        .I5(n3_reg[5]),
        .O(\n5[0]_i_2__8_n_0 ));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(\n9a_reg_n_0_[0] ),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(\n9a_reg_n_0_[1] ),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(\n9a_reg_n_0_[2] ),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(\n9a_reg_n_0_[3] ),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(\n9a_reg_n_0_[4] ),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(\n9a_reg_n_0_[5] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n11a_1[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n11a_1[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n11a_1[2]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n11a_1[3]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n11a_1[4]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n11a_1[5]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n9a_reg_rep[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[6]),
        .Q(n11a_1[6]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39923 n9m_reg_0_63_0_6
       (.ADDRA(n11a_1[5:0]),
        .ADDRB(n11a_1[5:0]),
        .ADDRC(n11a_1[5:0]),
        .ADDRD(n11a_1[5:0]),
        .ADDRE(n11a_1[5:0]),
        .ADDRF(n11a_1[5:0]),
        .ADDRG(n11a_1[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[0]),
        .DIB(i2[1]),
        .DIC(i2[2]),
        .DID(i2[3]),
        .DIE(i2[4]),
        .DIF(i2[5]),
        .DIG(i2[6]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_0_6_n_0),
        .DOB(n9m_reg_0_63_0_6_n_1),
        .DOC(n9m_reg_0_63_0_6_n_2),
        .DOD(n9m_reg_0_63_0_6_n_3),
        .DOE(n9m_reg_0_63_0_6_n_4),
        .DOF(n9m_reg_0_63_0_6_n_5),
        .DOG(n9m_reg_0_63_0_6_n_6),
        .DOH(NLW_n9m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39924 n9m_reg_0_63_14_20
       (.ADDRA(n11a_1[5:0]),
        .ADDRB(n11a_1[5:0]),
        .ADDRC(n11a_1[5:0]),
        .ADDRD(n11a_1[5:0]),
        .ADDRE(n11a_1[5:0]),
        .ADDRF(n11a_1[5:0]),
        .ADDRG(n11a_1[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[14]),
        .DIB(i2[15]),
        .DIC(i2[16]),
        .DID(i2[17]),
        .DIE(i2[18]),
        .DIF(i2[19]),
        .DIG(i2[20]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_14_20_n_0),
        .DOB(n9m_reg_0_63_14_20_n_1),
        .DOC(n9m_reg_0_63_14_20_n_2),
        .DOD(n9m_reg_0_63_14_20_n_3),
        .DOE(n9m_reg_0_63_14_20_n_4),
        .DOF(n9m_reg_0_63_14_20_n_5),
        .DOG(n9m_reg_0_63_14_20_n_6),
        .DOH(NLW_n9m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39925 n9m_reg_0_63_21_27
       (.ADDRA(n11a_1[5:0]),
        .ADDRB(n11a_1[5:0]),
        .ADDRC(n11a_1[5:0]),
        .ADDRD(n11a_1[5:0]),
        .ADDRE(n11a_1[5:0]),
        .ADDRF(n11a_1[5:0]),
        .ADDRG(n11a_1[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[21]),
        .DIB(i2[22]),
        .DIC(i2[23]),
        .DID(i2[24]),
        .DIE(i2[25]),
        .DIF(i2[26]),
        .DIG(i2[27]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_21_27_n_0),
        .DOB(n9m_reg_0_63_21_27_n_1),
        .DOC(n9m_reg_0_63_21_27_n_2),
        .DOD(n9m_reg_0_63_21_27_n_3),
        .DOE(n9m_reg_0_63_21_27_n_4),
        .DOF(n9m_reg_0_63_21_27_n_5),
        .DOG(n9m_reg_0_63_21_27_n_6),
        .DOH(NLW_n9m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39926 n9m_reg_0_63_28_31
       (.ADDRA(n11a_1[5:0]),
        .ADDRB(n11a_1[5:0]),
        .ADDRC(n11a_1[5:0]),
        .ADDRD(n11a_1[5:0]),
        .ADDRE(n11a_1[5:0]),
        .ADDRF(n11a_1[5:0]),
        .ADDRG(n11a_1[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[28]),
        .DIB(i2[29]),
        .DIC(i2[30]),
        .DID(i2[31]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_28_31_n_0),
        .DOB(n9m_reg_0_63_28_31_n_1),
        .DOC(n9m_reg_0_63_28_31_n_2),
        .DOD(n9m_reg_0_63_28_31_n_3),
        .DOE(NLW_n9m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n9m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39927 n9m_reg_0_63_7_13
       (.ADDRA(n11a_1[5:0]),
        .ADDRB(n11a_1[5:0]),
        .ADDRC(n11a_1[5:0]),
        .ADDRD(n11a_1[5:0]),
        .ADDRE(n11a_1[5:0]),
        .ADDRF(n11a_1[5:0]),
        .ADDRG(n11a_1[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[7]),
        .DIB(i2[8]),
        .DIC(i2[9]),
        .DID(i2[10]),
        .DIE(i2[11]),
        .DIF(i2[12]),
        .DIG(i2[13]),
        .DIH(1'b0),
        .DOA(n9m_reg_0_63_7_13_n_0),
        .DOB(n9m_reg_0_63_7_13_n_1),
        .DOC(n9m_reg_0_63_7_13_n_2),
        .DOD(n9m_reg_0_63_7_13_n_3),
        .DOE(n9m_reg_0_63_7_13_n_4),
        .DOF(n9m_reg_0_63_7_13_n_5),
        .DOG(n9m_reg_0_63_7_13_n_6),
        .DOH(NLW_n9m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(enable_i));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39928 n9m_reg_64_127_0_6
       (.ADDRA(n11a_1[5:0]),
        .ADDRB(n11a_1[5:0]),
        .ADDRC(n11a_1[5:0]),
        .ADDRD(n11a_1[5:0]),
        .ADDRE(n11a_1[5:0]),
        .ADDRF(n11a_1[5:0]),
        .ADDRG(n11a_1[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[0]),
        .DIB(i2[1]),
        .DIC(i2[2]),
        .DID(i2[3]),
        .DIE(i2[4]),
        .DIF(i2[5]),
        .DIG(i2[6]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_0_6_n_0),
        .DOB(n9m_reg_64_127_0_6_n_1),
        .DOC(n9m_reg_64_127_0_6_n_2),
        .DOD(n9m_reg_64_127_0_6_n_3),
        .DOE(n9m_reg_64_127_0_6_n_4),
        .DOF(n9m_reg_64_127_0_6_n_5),
        .DOG(n9m_reg_64_127_0_6_n_6),
        .DOH(NLW_n9m_reg_64_127_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39929 n9m_reg_64_127_14_20
       (.ADDRA(n11a_1[5:0]),
        .ADDRB(n11a_1[5:0]),
        .ADDRC(n11a_1[5:0]),
        .ADDRD(n11a_1[5:0]),
        .ADDRE(n11a_1[5:0]),
        .ADDRF(n11a_1[5:0]),
        .ADDRG(n11a_1[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[14]),
        .DIB(i2[15]),
        .DIC(i2[16]),
        .DID(i2[17]),
        .DIE(i2[18]),
        .DIF(i2[19]),
        .DIG(i2[20]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_14_20_n_0),
        .DOB(n9m_reg_64_127_14_20_n_1),
        .DOC(n9m_reg_64_127_14_20_n_2),
        .DOD(n9m_reg_64_127_14_20_n_3),
        .DOE(n9m_reg_64_127_14_20_n_4),
        .DOF(n9m_reg_64_127_14_20_n_5),
        .DOG(n9m_reg_64_127_14_20_n_6),
        .DOH(NLW_n9m_reg_64_127_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39930 n9m_reg_64_127_21_27
       (.ADDRA(n11a_1[5:0]),
        .ADDRB(n11a_1[5:0]),
        .ADDRC(n11a_1[5:0]),
        .ADDRD(n11a_1[5:0]),
        .ADDRE(n11a_1[5:0]),
        .ADDRF(n11a_1[5:0]),
        .ADDRG(n11a_1[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[21]),
        .DIB(i2[22]),
        .DIC(i2[23]),
        .DID(i2[24]),
        .DIE(i2[25]),
        .DIF(i2[26]),
        .DIG(i2[27]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_21_27_n_0),
        .DOB(n9m_reg_64_127_21_27_n_1),
        .DOC(n9m_reg_64_127_21_27_n_2),
        .DOD(n9m_reg_64_127_21_27_n_3),
        .DOE(n9m_reg_64_127_21_27_n_4),
        .DOF(n9m_reg_64_127_21_27_n_5),
        .DOG(n9m_reg_64_127_21_27_n_6),
        .DOH(NLW_n9m_reg_64_127_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39931 n9m_reg_64_127_28_31
       (.ADDRA(n11a_1[5:0]),
        .ADDRB(n11a_1[5:0]),
        .ADDRC(n11a_1[5:0]),
        .ADDRD(n11a_1[5:0]),
        .ADDRE(n11a_1[5:0]),
        .ADDRF(n11a_1[5:0]),
        .ADDRG(n11a_1[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[28]),
        .DIB(i2[29]),
        .DIC(i2[30]),
        .DID(i2[31]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_28_31_n_0),
        .DOB(n9m_reg_64_127_28_31_n_1),
        .DOC(n9m_reg_64_127_28_31_n_2),
        .DOD(n9m_reg_64_127_28_31_n_3),
        .DOE(NLW_n9m_reg_64_127_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n9m_reg_64_127_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n9m_reg_64_127_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n9m_reg_64_127_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s15/n9m" *) 
  (* ram_addr_begin = "64" *) 
  (* ram_addr_end = "127" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39932 n9m_reg_64_127_7_13
       (.ADDRA(n11a_1[5:0]),
        .ADDRB(n11a_1[5:0]),
        .ADDRC(n11a_1[5:0]),
        .ADDRD(n11a_1[5:0]),
        .ADDRE(n11a_1[5:0]),
        .ADDRF(n11a_1[5:0]),
        .ADDRG(n11a_1[5:0]),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[7]),
        .DIB(i2[8]),
        .DIC(i2[9]),
        .DID(i2[10]),
        .DIE(i2[11]),
        .DIF(i2[12]),
        .DIG(i2[13]),
        .DIH(1'b0),
        .DOA(n9m_reg_64_127_7_13_n_0),
        .DOB(n9m_reg_64_127_7_13_n_1),
        .DOC(n9m_reg_64_127_7_13_n_2),
        .DOD(n9m_reg_64_127_7_13_n_3),
        .DOE(n9m_reg_64_127_7_13_n_4),
        .DOF(n9m_reg_64_127_7_13_n_5),
        .DOG(n9m_reg_64_127_7_13_n_6),
        .DOH(NLW_n9m_reg_64_127_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_31" *) 
module switch_elements_cf_fft_512_8_31
   (i8,
    rst_i,
    enable_i,
    n4,
    clk_i);
  output [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input n4;
  input clk_i;

  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire n4;
  wire rst_i;

  FDRE #(
    .INIT(1'b0)) 
    \n5_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n4),
        .Q(i8),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_31" *) 
module switch_elements_cf_fft_512_8_31_0
   (i8,
    rst_i,
    enable_i,
    n4,
    clk_i);
  output [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input n4;
  input clk_i;

  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire n4;
  wire rst_i;

  FDRE #(
    .INIT(1'b0)) 
    \n5_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n4),
        .Q(i8),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_31" *) 
module switch_elements_cf_fft_512_8_31_1
   (i8,
    rst_i,
    enable_i,
    n4,
    clk_i);
  output [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input n4;
  input clk_i;

  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire n4;
  wire rst_i;

  FDRE #(
    .INIT(1'b0)) 
    \n5_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n4),
        .Q(i8),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_31" *) 
module switch_elements_cf_fft_512_8_31_10
   (i8,
    rst_i,
    enable_i,
    n4,
    clk_i);
  output [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input n4;
  input clk_i;

  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire n4;
  wire rst_i;

  FDRE #(
    .INIT(1'b0)) 
    \n5_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n4),
        .Q(i8),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_31" *) 
module switch_elements_cf_fft_512_8_31_13
   (i8,
    rst_i,
    enable_i,
    n4,
    clk_i);
  output [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input n4;
  input clk_i;

  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire n4;
  wire rst_i;

  FDRE #(
    .INIT(1'b0)) 
    \n5_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n4),
        .Q(i8),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_31" *) 
module switch_elements_cf_fft_512_8_31_16
   (i8,
    rst_i,
    enable_i,
    n4,
    clk_i);
  output [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input n4;
  input clk_i;

  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire n4;
  wire rst_i;

  FDRE #(
    .INIT(1'b0)) 
    \n5_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n4),
        .Q(i8),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_31" *) 
module switch_elements_cf_fft_512_8_31_19
   (i8,
    rst_i,
    enable_i,
    n4,
    clk_i);
  output [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input n4;
  input clk_i;

  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire n4;
  wire rst_i;

  FDRE #(
    .INIT(1'b0)) 
    \n5_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n4),
        .Q(i8),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_31" *) 
module switch_elements_cf_fft_512_8_31_23
   (i8,
    rst_i,
    enable_i,
    n4,
    clk_i);
  output [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input n4;
  input clk_i;

  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire n4;
  wire rst_i;

  FDRE #(
    .INIT(1'b0)) 
    \n5_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n4),
        .Q(i8),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_31" *) 
module switch_elements_cf_fft_512_8_31_4
   (i8,
    rst_i,
    enable_i,
    n4,
    clk_i);
  output [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input n4;
  input clk_i;

  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire n4;
  wire rst_i;

  FDRE #(
    .INIT(1'b0)) 
    \n5_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n4),
        .Q(i8),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_31" *) 
module switch_elements_cf_fft_512_8_31_7
   (i8,
    rst_i,
    enable_i,
    n4,
    clk_i);
  output [0:0]i8;
  input rst_i;
  input [0:0]enable_i;
  input n4;
  input clk_i;

  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire n4;
  wire rst_i;

  FDRE #(
    .INIT(1'b0)) 
    \n5_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n4),
        .Q(i8),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_37" *) 
module switch_elements_cf_fft_512_8_37
   (i1,
    enable_i,
    clk_i,
    rst_i,
    i3,
    i2);
  output [29:0]i1;
  input [0:0]enable_i;
  input clk_i;
  input rst_i;
  input [15:0]i3;
  input [15:0]i2;

  wire [6:6]B;
  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [15:0]i2;
  wire [15:0]i3;
  wire [7:0]n10;
  wire n14__21_carry__0_i_1_n_0;
  wire n14__21_carry__0_i_2__0_n_0;
  wire n14__21_carry__0_i_3_n_0;
  wire n14__21_carry__0_i_4__0_n_0;
  wire n14__21_carry__0_n_14;
  wire n14__21_carry__0_n_15;
  wire n14__21_carry__0_n_5;
  wire n14__21_carry__0_n_7;
  wire n14__21_carry_i_10__0_n_0;
  wire n14__21_carry_i_11_n_0;
  wire n14__21_carry_i_12_n_0;
  wire n14__21_carry_i_13_n_0;
  wire n14__21_carry_i_14_n_0;
  wire n14__21_carry_i_1__0_n_0;
  wire n14__21_carry_i_2__0_n_0;
  wire n14__21_carry_i_3__0_n_0;
  wire n14__21_carry_i_4__0_n_0;
  wire n14__21_carry_i_5__0_n_0;
  wire n14__21_carry_i_6_n_0;
  wire n14__21_carry_i_7_n_0;
  wire n14__21_carry_i_8__0_n_0;
  wire n14__21_carry_i_9_n_0;
  wire n14__21_carry_n_0;
  wire n14__21_carry_n_1;
  wire n14__21_carry_n_10;
  wire n14__21_carry_n_11;
  wire n14__21_carry_n_12;
  wire n14__21_carry_n_13;
  wire n14__21_carry_n_14;
  wire n14__21_carry_n_2;
  wire n14__21_carry_n_3;
  wire n14__21_carry_n_4;
  wire n14__21_carry_n_5;
  wire n14__21_carry_n_6;
  wire n14__21_carry_n_7;
  wire n14__21_carry_n_8;
  wire n14__21_carry_n_9;
  wire n14__47_carry_i_10_n_0;
  wire n14__47_carry_i_11_n_0;
  wire n14__47_carry_i_12_n_0;
  wire n14__47_carry_i_1__0_n_0;
  wire n14__47_carry_i_2__0_n_0;
  wire n14__47_carry_i_3_n_0;
  wire n14__47_carry_i_4_n_0;
  wire n14__47_carry_i_5_n_0;
  wire n14__47_carry_i_6__0_n_0;
  wire n14__47_carry_i_7_n_0;
  wire n14__47_carry_i_8_n_0;
  wire n14__47_carry_i_9_n_0;
  wire n14__47_carry_n_1;
  wire n14__47_carry_n_10;
  wire n14__47_carry_n_11;
  wire n14__47_carry_n_12;
  wire n14__47_carry_n_13;
  wire n14__47_carry_n_14;
  wire n14__47_carry_n_15;
  wire n14__47_carry_n_2;
  wire n14__47_carry_n_3;
  wire n14__47_carry_n_4;
  wire n14__47_carry_n_5;
  wire n14__47_carry_n_6;
  wire n14__47_carry_n_7;
  wire n14__47_carry_n_8;
  wire n14__47_carry_n_9;
  wire n14__67_carry__0_i_1__0_n_0;
  wire n14__67_carry__0_i_2__0_n_0;
  wire n14__67_carry__0_i_3__0_n_0;
  wire n14__67_carry__0_i_4__0_n_0;
  wire n14__67_carry__0_i_5__0_n_0;
  wire n14__67_carry__0_i_6__0_n_0;
  wire n14__67_carry__0_i_7__0_n_0;
  wire n14__67_carry__0_n_5;
  wire n14__67_carry__0_n_6;
  wire n14__67_carry__0_n_7;
  wire n14__67_carry_i_10__0_n_0;
  wire n14__67_carry_i_11__0_n_0;
  wire n14__67_carry_i_12__0_n_0;
  wire n14__67_carry_i_13__0_n_0;
  wire n14__67_carry_i_14__0_n_0;
  wire n14__67_carry_i_15__0_n_0;
  wire n14__67_carry_i_1__0_n_0;
  wire n14__67_carry_i_2__0_n_0;
  wire n14__67_carry_i_3__0_n_0;
  wire n14__67_carry_i_4__0_n_0;
  wire n14__67_carry_i_5__0_n_0;
  wire n14__67_carry_i_6__0_n_0;
  wire n14__67_carry_i_7__0_n_0;
  wire n14__67_carry_i_8__0_n_0;
  wire n14__67_carry_i_9__0_n_0;
  wire n14__67_carry_n_0;
  wire n14__67_carry_n_1;
  wire n14__67_carry_n_2;
  wire n14__67_carry_n_3;
  wire n14__67_carry_n_4;
  wire n14__67_carry_n_5;
  wire n14__67_carry_n_6;
  wire n14__67_carry_n_7;
  wire n14_carry__0_i_1__0_n_0;
  wire n14_carry__0_i_2__0_n_0;
  wire n14_carry__0_i_3_n_0;
  wire n14_carry__0_i_4__0_n_0;
  wire n14_carry__0_n_14;
  wire n14_carry__0_n_15;
  wire n14_carry__0_n_5;
  wire n14_carry__0_n_7;
  wire n14_carry_i_10__0_n_0;
  wire n14_carry_i_11__0_n_0;
  wire n14_carry_i_12__0_n_0;
  wire n14_carry_i_13_n_0;
  wire n14_carry_i_14_n_0;
  wire n14_carry_i_15_n_0;
  wire n14_carry_i_1__0_n_0;
  wire n14_carry_i_2__0_n_0;
  wire n14_carry_i_3__0_n_0;
  wire n14_carry_i_4__0_n_0;
  wire n14_carry_i_5__0_n_0;
  wire n14_carry_i_6__0_n_0;
  wire n14_carry_i_7_n_0;
  wire n14_carry_i_8_n_0;
  wire n14_carry_i_9__0_n_0;
  wire n14_carry_n_0;
  wire n14_carry_n_1;
  wire n14_carry_n_10;
  wire n14_carry_n_11;
  wire n14_carry_n_12;
  wire n14_carry_n_15;
  wire n14_carry_n_2;
  wire n14_carry_n_3;
  wire n14_carry_n_4;
  wire n14_carry_n_5;
  wire n14_carry_n_6;
  wire n14_carry_n_7;
  wire n14_carry_n_8;
  wire n14_carry_n_9;
  wire [7:0]n15;
  wire \n16_reg_n_0_[0] ;
  wire \n16_reg_n_0_[1] ;
  wire \n16_reg_n_0_[2] ;
  wire \n16_reg_n_0_[3] ;
  wire \n16_reg_n_0_[4] ;
  wire \n16_reg_n_0_[5] ;
  wire \n16_reg_n_0_[6] ;
  wire \n16_reg_n_0_[7] ;
  wire \n1_reg_n_0_[0] ;
  wire \n1_reg_n_0_[1] ;
  wire \n1_reg_n_0_[2] ;
  wire \n1_reg_n_0_[3] ;
  wire \n1_reg_n_0_[4] ;
  wire \n1_reg_n_0_[5] ;
  wire \n1_reg_n_0_[6] ;
  wire \n1_reg_n_0_[7] ;
  wire [7:0]n2;
  wire [7:0]n202_out;
  wire [7:0]n21;
  wire \n21[7]_i_2_n_0 ;
  wire \n21[7]_i_3_n_0 ;
  wire \n21[7]_i_4_n_0 ;
  wire \n21[7]_i_5_n_0 ;
  wire \n21[7]_i_6_n_0 ;
  wire \n21[7]_i_7_n_0 ;
  wire \n21[7]_i_8_n_0 ;
  wire \n21[7]_i_9_n_0 ;
  wire \n21_reg[7]_i_1__2_n_1 ;
  wire \n21_reg[7]_i_1__2_n_2 ;
  wire \n21_reg[7]_i_1__2_n_3 ;
  wire \n21_reg[7]_i_1__2_n_4 ;
  wire \n21_reg[7]_i_1__2_n_5 ;
  wire \n21_reg[7]_i_1__2_n_6 ;
  wire \n21_reg[7]_i_1__2_n_7 ;
  wire n22__0_n_0;
  wire n22__1_n_0;
  wire n22__2_n_0;
  wire n22__3_n_0;
  wire n22__4_n_0;
  wire n22__5_n_0;
  wire n22__6_n_0;
  wire n22_n_0;
  wire n25__17_carry__0_i_1_n_0;
  wire n25__17_carry__0_i_2__0_n_0;
  wire n25__17_carry__0_i_3_n_0;
  wire n25__17_carry__0_i_4__0_n_0;
  wire n25__17_carry__0_n_14;
  wire n25__17_carry__0_n_15;
  wire n25__17_carry__0_n_5;
  wire n25__17_carry__0_n_7;
  wire n25__17_carry_i_10__0_n_0;
  wire n25__17_carry_i_11_n_0;
  wire n25__17_carry_i_12_n_0;
  wire n25__17_carry_i_13_n_0;
  wire n25__17_carry_i_14_n_0;
  wire n25__17_carry_i_1__0_n_0;
  wire n25__17_carry_i_2__0_n_0;
  wire n25__17_carry_i_3__0_n_0;
  wire n25__17_carry_i_4__0_n_0;
  wire n25__17_carry_i_5__0_n_0;
  wire n25__17_carry_i_6_n_0;
  wire n25__17_carry_i_7_n_0;
  wire n25__17_carry_i_8__0_n_0;
  wire n25__17_carry_i_9_n_0;
  wire n25__17_carry_n_0;
  wire n25__17_carry_n_1;
  wire n25__17_carry_n_10;
  wire n25__17_carry_n_11;
  wire n25__17_carry_n_12;
  wire n25__17_carry_n_13;
  wire n25__17_carry_n_14;
  wire n25__17_carry_n_2;
  wire n25__17_carry_n_3;
  wire n25__17_carry_n_4;
  wire n25__17_carry_n_5;
  wire n25__17_carry_n_6;
  wire n25__17_carry_n_7;
  wire n25__17_carry_n_8;
  wire n25__17_carry_n_9;
  wire n25__47_carry_i_10_n_0;
  wire n25__47_carry_i_11_n_0;
  wire n25__47_carry_i_12_n_0;
  wire n25__47_carry_i_1__0_n_0;
  wire n25__47_carry_i_2__0_n_0;
  wire n25__47_carry_i_3_n_0;
  wire n25__47_carry_i_4_n_0;
  wire n25__47_carry_i_5_n_0;
  wire n25__47_carry_i_6__0_n_0;
  wire n25__47_carry_i_7_n_0;
  wire n25__47_carry_i_8_n_0;
  wire n25__47_carry_i_9_n_0;
  wire n25__47_carry_n_1;
  wire n25__47_carry_n_10;
  wire n25__47_carry_n_11;
  wire n25__47_carry_n_12;
  wire n25__47_carry_n_13;
  wire n25__47_carry_n_14;
  wire n25__47_carry_n_15;
  wire n25__47_carry_n_2;
  wire n25__47_carry_n_3;
  wire n25__47_carry_n_4;
  wire n25__47_carry_n_5;
  wire n25__47_carry_n_6;
  wire n25__47_carry_n_7;
  wire n25__47_carry_n_8;
  wire n25__47_carry_n_9;
  wire n25__67_carry__0_i_1__0_n_0;
  wire n25__67_carry__0_i_2__0_n_0;
  wire n25__67_carry__0_i_3__0_n_0;
  wire n25__67_carry__0_i_4__0_n_0;
  wire n25__67_carry__0_i_5__0_n_0;
  wire n25__67_carry__0_i_6__0_n_0;
  wire n25__67_carry__0_i_7__0_n_0;
  wire n25__67_carry__0_n_5;
  wire n25__67_carry__0_n_6;
  wire n25__67_carry__0_n_7;
  wire n25__67_carry_i_10__0_n_0;
  wire n25__67_carry_i_11__0_n_0;
  wire n25__67_carry_i_12__0_n_0;
  wire n25__67_carry_i_13__0_n_0;
  wire n25__67_carry_i_14__0_n_0;
  wire n25__67_carry_i_15__0_n_0;
  wire n25__67_carry_i_1__0_n_0;
  wire n25__67_carry_i_2__0_n_0;
  wire n25__67_carry_i_3__0_n_0;
  wire n25__67_carry_i_4__0_n_0;
  wire n25__67_carry_i_5__0_n_0;
  wire n25__67_carry_i_6__0_n_0;
  wire n25__67_carry_i_7__0_n_0;
  wire n25__67_carry_i_8__0_n_0;
  wire n25__67_carry_i_9__0_n_0;
  wire n25__67_carry_n_0;
  wire n25__67_carry_n_1;
  wire n25__67_carry_n_2;
  wire n25__67_carry_n_3;
  wire n25__67_carry_n_4;
  wire n25__67_carry_n_5;
  wire n25__67_carry_n_6;
  wire n25__67_carry_n_7;
  wire n25_carry__0_i_1__0_n_0;
  wire n25_carry__0_i_2__0_n_0;
  wire n25_carry__0_i_3_n_0;
  wire n25_carry__0_i_4__0_n_0;
  wire n25_carry__0_n_14;
  wire n25_carry__0_n_15;
  wire n25_carry__0_n_5;
  wire n25_carry__0_n_7;
  wire n25_carry_i_10__0_n_0;
  wire n25_carry_i_11__0_n_0;
  wire n25_carry_i_12__0_n_0;
  wire n25_carry_i_13_n_0;
  wire n25_carry_i_14_n_0;
  wire n25_carry_i_15_n_0;
  wire n25_carry_i_1__0_n_0;
  wire n25_carry_i_2__0_n_0;
  wire n25_carry_i_3__0_n_0;
  wire n25_carry_i_4__0_n_0;
  wire n25_carry_i_5__0_n_0;
  wire n25_carry_i_6__0_n_0;
  wire n25_carry_i_7_n_0;
  wire n25_carry_i_8_n_0;
  wire n25_carry_i_9__0_n_0;
  wire n25_carry_n_0;
  wire n25_carry_n_1;
  wire n25_carry_n_10;
  wire n25_carry_n_11;
  wire n25_carry_n_12;
  wire n25_carry_n_15;
  wire n25_carry_n_2;
  wire n25_carry_n_3;
  wire n25_carry_n_4;
  wire n25_carry_n_5;
  wire n25_carry_n_6;
  wire n25_carry_n_7;
  wire n25_carry_n_8;
  wire n25_carry_n_9;
  wire [7:0]n26;
  wire [7:0]n27;
  wire [7:0]n29;
  wire [7:7]n30;
  wire [7:0]n31;
  wire \n33[10]_i_1__6_n_0 ;
  wire \n33[11]_i_1__6_n_0 ;
  wire \n33[12]_i_1__6_n_0 ;
  wire \n33[12]_i_2__6_n_0 ;
  wire \n33[13]_i_1__6_n_0 ;
  wire \n33[14]_i_1__6_n_0 ;
  wire \n33[14]_i_2__6_n_0 ;
  wire \n33[15]_i_2__6_n_0 ;
  wire \n33[2]_i_1__6_n_0 ;
  wire \n33[3]_i_1__6_n_0 ;
  wire \n33[4]_i_1__6_n_0 ;
  wire \n33[4]_i_2__6_n_0 ;
  wire \n33[5]_i_1__6_n_0 ;
  wire \n33[6]_i_1__6_n_0 ;
  wire \n33[6]_i_2__6_n_0 ;
  wire \n33[7]_i_2__6_n_0 ;
  wire \n33[9]_i_1__6_n_0 ;
  wire [7:0]n341_out;
  wire [7:1]n350_out;
  wire \n37[12]_i_2__6_n_0 ;
  wire \n37[14]_i_2__6_n_0 ;
  wire \n37[15]_i_2__6_n_0 ;
  wire \n37[4]_i_2__6_n_0 ;
  wire \n37[6]_i_2__6_n_0 ;
  wire \n37[7]_i_2__6_n_0 ;
  wire [7:0]n4;
  wire \n7_reg_n_0_[0] ;
  wire \n7_reg_n_0_[1] ;
  wire \n7_reg_n_0_[2] ;
  wire \n7_reg_n_0_[3] ;
  wire \n7_reg_n_0_[4] ;
  wire \n7_reg_n_0_[5] ;
  wire \n7_reg_n_0_[6] ;
  wire \n7_reg_n_0_[7] ;
  wire \n8_reg_n_0_[0] ;
  wire \n8_reg_n_0_[1] ;
  wire \n8_reg_n_0_[2] ;
  wire \n8_reg_n_0_[3] ;
  wire \n8_reg_n_0_[4] ;
  wire \n8_reg_n_0_[5] ;
  wire \n8_reg_n_0_[6] ;
  wire \n8_reg_n_0_[7] ;
  wire \n9_reg_n_0_[0] ;
  wire \n9_reg_n_0_[1] ;
  wire \n9_reg_n_0_[2] ;
  wire \n9_reg_n_0_[3] ;
  wire \n9_reg_n_0_[4] ;
  wire \n9_reg_n_0_[5] ;
  wire \n9_reg_n_0_[6] ;
  wire \n9_reg_n_0_[7] ;
  wire rst_i;
  wire [0:0]NLW_n14__21_carry_O_UNCONNECTED;
  wire [7:1]NLW_n14__21_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n14__21_carry__0_O_UNCONNECTED;
  wire [7:7]NLW_n14__47_carry_CO_UNCONNECTED;
  wire [3:0]NLW_n14__67_carry_O_UNCONNECTED;
  wire [7:3]NLW_n14__67_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n14__67_carry__0_O_UNCONNECTED;
  wire [2:1]NLW_n14_carry_O_UNCONNECTED;
  wire [7:1]NLW_n14_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n14_carry__0_O_UNCONNECTED;
  wire [7:7]\NLW_n21_reg[7]_i_1__2_CO_UNCONNECTED ;
  wire [0:0]NLW_n25__17_carry_O_UNCONNECTED;
  wire [7:1]NLW_n25__17_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n25__17_carry__0_O_UNCONNECTED;
  wire [7:7]NLW_n25__47_carry_CO_UNCONNECTED;
  wire [3:0]NLW_n25__67_carry_O_UNCONNECTED;
  wire [7:3]NLW_n25__67_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n25__67_carry__0_O_UNCONNECTED;
  wire [2:1]NLW_n25_carry_O_UNCONNECTED;
  wire [7:1]NLW_n25_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n25_carry__0_O_UNCONNECTED;

  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[0] ),
        .Q(n10[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[1] ),
        .Q(n10[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[2] ),
        .Q(n10[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[3] ),
        .Q(n10[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[4] ),
        .Q(n10[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[5] ),
        .Q(n10[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[6] ),
        .Q(n10[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[7] ),
        .Q(n10[7]),
        .R(rst_i));
  FDSE #(
    .INIT(1'b0)) 
    \n11_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(1'b0),
        .Q(B),
        .S(enable_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__21_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__21_carry_n_0,n14__21_carry_n_1,n14__21_carry_n_2,n14__21_carry_n_3,n14__21_carry_n_4,n14__21_carry_n_5,n14__21_carry_n_6,n14__21_carry_n_7}),
        .DI({n14_carry_i_1__0_n_0,n14__21_carry_i_1__0_n_0,n14__21_carry_i_2__0_n_0,n14__21_carry_i_3__0_n_0,n14__21_carry_i_4__0_n_0,n14__21_carry_i_5__0_n_0,n14__21_carry_i_6_n_0,1'b0}),
        .O({n14__21_carry_n_8,n14__21_carry_n_9,n14__21_carry_n_10,n14__21_carry_n_11,n14__21_carry_n_12,n14__21_carry_n_13,n14__21_carry_n_14,NLW_n14__21_carry_O_UNCONNECTED[0]}),
        .S({n14__21_carry_i_7_n_0,n14__21_carry_i_8__0_n_0,n14__21_carry_i_9_n_0,n14__21_carry_i_10__0_n_0,n14__21_carry_i_11_n_0,n14__21_carry_i_12_n_0,n14__21_carry_i_13_n_0,n14__21_carry_i_14_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__21_carry__0
       (.CI(n14__21_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__21_carry__0_CO_UNCONNECTED[7:3],n14__21_carry__0_n_5,NLW_n14__21_carry__0_CO_UNCONNECTED[1],n14__21_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14__21_carry__0_i_1_n_0,n14__21_carry__0_i_2__0_n_0}),
        .O({NLW_n14__21_carry__0_O_UNCONNECTED[7:2],n14__21_carry__0_n_14,n14__21_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n14__21_carry__0_i_3_n_0,n14__21_carry__0_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h40)) 
    n14__21_carry__0_i_1
       (.I0(n22_n_0),
        .I1(B),
        .I2(n22__0_n_0),
        .O(n14__21_carry__0_i_1_n_0));
  LUT4 #(
    .INIT(16'h80C8)) 
    n14__21_carry__0_i_2__0
       (.I0(n22__1_n_0),
        .I1(B),
        .I2(n22__0_n_0),
        .I3(n22_n_0),
        .O(n14__21_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h37)) 
    n14__21_carry__0_i_3
       (.I0(n22__0_n_0),
        .I1(B),
        .I2(n22_n_0),
        .O(n14__21_carry__0_i_3_n_0));
  LUT4 #(
    .INIT(16'h4FDF)) 
    n14__21_carry__0_i_4__0
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(B),
        .I3(n22_n_0),
        .O(n14__21_carry__0_i_4__0_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n14__21_carry_i_10__0
       (.I0(n22__5_n_0),
        .I1(n22__3_n_0),
        .I2(B),
        .I3(n22__4_n_0),
        .I4(n22__2_n_0),
        .O(n14__21_carry_i_10__0_n_0));
  LUT5 #(
    .INIT(32'h66009600)) 
    n14__21_carry_i_11
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__5_n_0),
        .I3(B),
        .I4(n22__6_n_0),
        .O(n14__21_carry_i_11_n_0));
  LUT4 #(
    .INIT(16'h9060)) 
    n14__21_carry_i_12
       (.I0(n22__6_n_0),
        .I1(n22__5_n_0),
        .I2(B),
        .I3(n22__4_n_0),
        .O(n14__21_carry_i_12_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n14__21_carry_i_13
       (.I0(n22__5_n_0),
        .I1(B),
        .I2(n22__6_n_0),
        .O(n14__21_carry_i_13_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__21_carry_i_14
       (.I0(B),
        .I1(n22__6_n_0),
        .O(n14__21_carry_i_14_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n14__21_carry_i_1__0
       (.I0(n22__3_n_0),
        .I1(B),
        .I2(n22__2_n_0),
        .I3(n22__1_n_0),
        .O(n14__21_carry_i_1__0_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n14__21_carry_i_2__0
       (.I0(n22__4_n_0),
        .I1(B),
        .I2(n22__3_n_0),
        .I3(n22__2_n_0),
        .O(n14__21_carry_i_2__0_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n14__21_carry_i_3__0
       (.I0(n22__5_n_0),
        .I1(B),
        .I2(n22__4_n_0),
        .I3(n22__3_n_0),
        .O(n14__21_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h8448)) 
    n14__21_carry_i_4__0
       (.I0(n22__4_n_0),
        .I1(B),
        .I2(n22__5_n_0),
        .I3(n22__3_n_0),
        .O(n14__21_carry_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n14__21_carry_i_5__0
       (.I0(n22__5_n_0),
        .I1(B),
        .I2(n22__6_n_0),
        .O(n14__21_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__21_carry_i_6
       (.I0(B),
        .I1(n22__5_n_0),
        .O(n14__21_carry_i_6_n_0));
  LUT5 #(
    .INIT(32'h95656595)) 
    n14__21_carry_i_7
       (.I0(n14_carry_i_1__0_n_0),
        .I1(n22__0_n_0),
        .I2(B),
        .I3(n22__1_n_0),
        .I4(n22_n_0),
        .O(n14__21_carry_i_7_n_0));
  (* HLUTNM = "lutpair106" *) 
  LUT5 #(
    .INIT(32'h4C8004C8)) 
    n14__21_carry_i_8__0
       (.I0(n22__2_n_0),
        .I1(B),
        .I2(n22__1_n_0),
        .I3(n22__0_n_0),
        .I4(n22__3_n_0),
        .O(n14__21_carry_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n14__21_carry_i_9
       (.I0(n22__4_n_0),
        .I1(n22__2_n_0),
        .I2(B),
        .I3(n22__3_n_0),
        .I4(n22__1_n_0),
        .O(n14__21_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__47_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__47_carry_CO_UNCONNECTED[7],n14__47_carry_n_1,n14__47_carry_n_2,n14__47_carry_n_3,n14__47_carry_n_4,n14__47_carry_n_5,n14__47_carry_n_6,n14__47_carry_n_7}),
        .DI({1'b0,n14__47_carry_i_1__0_n_0,n14__47_carry_i_2__0_n_0,n14__47_carry_i_3_n_0,n14__47_carry_i_4_n_0,1'b1,1'b0,1'b1}),
        .O({n14__47_carry_n_8,n14__47_carry_n_9,n14__47_carry_n_10,n14__47_carry_n_11,n14__47_carry_n_12,n14__47_carry_n_13,n14__47_carry_n_14,n14__47_carry_n_15}),
        .S({n14__47_carry_i_5_n_0,n14__47_carry_i_6__0_n_0,n14__47_carry_i_7_n_0,n14__47_carry_i_8_n_0,n14__47_carry_i_9_n_0,n14__47_carry_i_10_n_0,n14__47_carry_i_11_n_0,n14__47_carry_i_12_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n14__47_carry_i_10
       (.I0(B),
        .I1(n22__3_n_0),
        .O(n14__47_carry_i_10_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__47_carry_i_11
       (.I0(B),
        .I1(n22__4_n_0),
        .O(n14__47_carry_i_11_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n14__47_carry_i_12
       (.I0(n22__5_n_0),
        .I1(B),
        .O(n14__47_carry_i_12_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__47_carry_i_1__0
       (.I0(B),
        .I1(n22__0_n_0),
        .O(n14__47_carry_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__47_carry_i_2__0
       (.I0(B),
        .I1(n22__1_n_0),
        .O(n14__47_carry_i_2__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__47_carry_i_3
       (.I0(B),
        .I1(n22__2_n_0),
        .O(n14__47_carry_i_3_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__47_carry_i_4
       (.I0(B),
        .I1(n22__3_n_0),
        .O(n14__47_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n14__47_carry_i_5
       (.I0(n22_n_0),
        .I1(B),
        .O(n14__47_carry_i_5_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n14__47_carry_i_6__0
       (.I0(n22__0_n_0),
        .I1(B),
        .I2(n22_n_0),
        .O(n14__47_carry_i_6__0_n_0));
  LUT3 #(
    .INIT(8'hB7)) 
    n14__47_carry_i_7
       (.I0(n22__1_n_0),
        .I1(B),
        .I2(n22__0_n_0),
        .O(n14__47_carry_i_7_n_0));
  LUT3 #(
    .INIT(8'hB7)) 
    n14__47_carry_i_8
       (.I0(n22__2_n_0),
        .I1(B),
        .I2(n22__1_n_0),
        .O(n14__47_carry_i_8_n_0));
  LUT3 #(
    .INIT(8'hB7)) 
    n14__47_carry_i_9
       (.I0(n22__3_n_0),
        .I1(B),
        .I2(n22__2_n_0),
        .O(n14__47_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__67_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__67_carry_n_0,n14__67_carry_n_1,n14__67_carry_n_2,n14__67_carry_n_3,n14__67_carry_n_4,n14__67_carry_n_5,n14__67_carry_n_6,n14__67_carry_n_7}),
        .DI({n14__67_carry_i_1__0_n_0,n14__67_carry_i_2__0_n_0,n14__67_carry_i_3__0_n_0,n14__67_carry_i_4__0_n_0,n14__67_carry_i_5__0_n_0,n14__67_carry_i_6__0_n_0,n14__67_carry_i_7__0_n_0,1'b0}),
        .O({n15[3:0],NLW_n14__67_carry_O_UNCONNECTED[3:0]}),
        .S({n14__67_carry_i_8__0_n_0,n14__67_carry_i_9__0_n_0,n14__67_carry_i_10__0_n_0,n14__67_carry_i_11__0_n_0,n14__67_carry_i_12__0_n_0,n14__67_carry_i_13__0_n_0,n14__67_carry_i_14__0_n_0,n14__67_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__67_carry__0
       (.CI(n14__67_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__67_carry__0_CO_UNCONNECTED[7:3],n14__67_carry__0_n_5,n14__67_carry__0_n_6,n14__67_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n14__67_carry__0_i_1__0_n_0,n14__67_carry__0_i_2__0_n_0,n14__67_carry__0_i_3__0_n_0}),
        .O({NLW_n14__67_carry__0_O_UNCONNECTED[7:4],n15[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n14__67_carry__0_i_4__0_n_0,n14__67_carry__0_i_5__0_n_0,n14__67_carry__0_i_6__0_n_0,n14__67_carry__0_i_7__0_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry__0_i_1__0
       (.I0(n14__21_carry__0_n_14),
        .I1(n14__47_carry_n_10),
        .O(n14__67_carry__0_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry__0_i_2__0
       (.I0(n14__21_carry__0_n_15),
        .I1(n14__47_carry_n_11),
        .O(n14__67_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14__67_carry__0_i_3__0
       (.I0(n14__47_carry_n_12),
        .I1(n14__21_carry_n_8),
        .I2(n14_carry__0_n_5),
        .O(n14__67_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n14__67_carry__0_i_4__0
       (.I0(n14__21_carry__0_n_5),
        .I1(n14__47_carry_n_9),
        .I2(n14__47_carry_n_8),
        .O(n14__67_carry__0_i_4__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__67_carry__0_i_5__0
       (.I0(n14__21_carry__0_n_14),
        .I1(n14__47_carry_n_10),
        .I2(n14__47_carry_n_9),
        .I3(n14__21_carry__0_n_5),
        .O(n14__67_carry__0_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__67_carry__0_i_6__0
       (.I0(n14__21_carry__0_n_15),
        .I1(n14__47_carry_n_11),
        .I2(n14__47_carry_n_10),
        .I3(n14__21_carry__0_n_14),
        .O(n14__67_carry__0_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n14__67_carry__0_i_7__0
       (.I0(n14_carry__0_n_5),
        .I1(n14__21_carry_n_8),
        .I2(n14__47_carry_n_12),
        .I3(n14__47_carry_n_11),
        .I4(n14__21_carry__0_n_15),
        .O(n14__67_carry__0_i_7__0_n_0));
  (* HLUTNM = "lutpair70" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__67_carry_i_10__0
       (.I0(n14__47_carry_n_14),
        .I1(n14__21_carry_n_10),
        .I2(n14_carry__0_n_15),
        .I3(n14__67_carry_i_3__0_n_0),
        .O(n14__67_carry_i_10__0_n_0));
  (* HLUTNM = "lutpair69" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__67_carry_i_11__0
       (.I0(n14__47_carry_n_15),
        .I1(n14__21_carry_n_11),
        .I2(n14_carry_n_8),
        .I3(n14__67_carry_i_4__0_n_0),
        .O(n14__67_carry_i_11__0_n_0));
  (* HLUTNM = "lutpair68" *) 
  LUT5 #(
    .INIT(32'h78878778)) 
    n14__67_carry_i_12__0
       (.I0(B),
        .I1(n22__6_n_0),
        .I2(n14__21_carry_n_12),
        .I3(n14_carry_n_9),
        .I4(n14__67_carry_i_5__0_n_0),
        .O(n14__67_carry_i_12__0_n_0));
  (* HLUTNM = "lutpair107" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n14__67_carry_i_13__0
       (.I0(n14__21_carry_n_13),
        .I1(n14_carry_n_10),
        .I2(n14_carry_n_11),
        .I3(n14__21_carry_n_14),
        .O(n14__67_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__67_carry_i_14__0
       (.I0(n14_carry_n_12),
        .I1(n14_carry_n_15),
        .I2(n14__21_carry_n_14),
        .I3(n14_carry_n_11),
        .O(n14__67_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n14__67_carry_i_15__0
       (.I0(n14_carry_n_12),
        .I1(n14_carry_n_15),
        .O(n14__67_carry_i_15__0_n_0));
  (* HLUTNM = "lutpair71" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__67_carry_i_1__0
       (.I0(n14__47_carry_n_13),
        .I1(n14__21_carry_n_9),
        .I2(n14_carry__0_n_14),
        .O(n14__67_carry_i_1__0_n_0));
  (* HLUTNM = "lutpair70" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__67_carry_i_2__0
       (.I0(n14__47_carry_n_14),
        .I1(n14__21_carry_n_10),
        .I2(n14_carry__0_n_15),
        .O(n14__67_carry_i_2__0_n_0));
  (* HLUTNM = "lutpair69" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__67_carry_i_3__0
       (.I0(n14__47_carry_n_15),
        .I1(n14__21_carry_n_11),
        .I2(n14_carry_n_8),
        .O(n14__67_carry_i_3__0_n_0));
  (* HLUTNM = "lutpair68" *) 
  LUT4 #(
    .INIT(16'hF880)) 
    n14__67_carry_i_4__0
       (.I0(B),
        .I1(n22__6_n_0),
        .I2(n14__21_carry_n_12),
        .I3(n14_carry_n_9),
        .O(n14__67_carry_i_4__0_n_0));
  (* HLUTNM = "lutpair107" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry_i_5__0
       (.I0(n14__21_carry_n_13),
        .I1(n14_carry_n_10),
        .O(n14__67_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry_i_6__0
       (.I0(n14_carry_n_11),
        .I1(n14__21_carry_n_14),
        .O(n14__67_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry_i_7__0
       (.I0(n14_carry_n_12),
        .I1(n14_carry_n_15),
        .O(n14__67_carry_i_7__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n14__67_carry_i_8__0
       (.I0(n14__67_carry_i_1__0_n_0),
        .I1(n14__21_carry_n_8),
        .I2(n14__47_carry_n_12),
        .I3(n14_carry__0_n_5),
        .O(n14__67_carry_i_8__0_n_0));
  (* HLUTNM = "lutpair71" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__67_carry_i_9__0
       (.I0(n14__47_carry_n_13),
        .I1(n14__21_carry_n_9),
        .I2(n14_carry__0_n_14),
        .I3(n14__67_carry_i_2__0_n_0),
        .O(n14__67_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14_carry_n_0,n14_carry_n_1,n14_carry_n_2,n14_carry_n_3,n14_carry_n_4,n14_carry_n_5,n14_carry_n_6,n14_carry_n_7}),
        .DI({n14_carry_i_1__0_n_0,n14_carry_i_2__0_n_0,n14_carry_i_3__0_n_0,n14_carry_i_4__0_n_0,n14_carry_i_5__0_n_0,n14_carry_i_6__0_n_0,n14_carry_i_7_n_0,1'b0}),
        .O({n14_carry_n_8,n14_carry_n_9,n14_carry_n_10,n14_carry_n_11,n14_carry_n_12,NLW_n14_carry_O_UNCONNECTED[2:1],n14_carry_n_15}),
        .S({n14_carry_i_8_n_0,n14_carry_i_9__0_n_0,n14_carry_i_10__0_n_0,n14_carry_i_11__0_n_0,n14_carry_i_12__0_n_0,n14_carry_i_13_n_0,n14_carry_i_14_n_0,n14_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14_carry__0
       (.CI(n14_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14_carry__0_CO_UNCONNECTED[7:3],n14_carry__0_n_5,NLW_n14_carry__0_CO_UNCONNECTED[1],n14_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14_carry__0_i_1__0_n_0,n14_carry__0_i_2__0_n_0}),
        .O({NLW_n14_carry__0_O_UNCONNECTED[7:2],n14_carry__0_n_14,n14_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n14_carry__0_i_3_n_0,n14_carry__0_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h40)) 
    n14_carry__0_i_1__0
       (.I0(n22_n_0),
        .I1(B),
        .I2(n22__0_n_0),
        .O(n14_carry__0_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h80C8)) 
    n14_carry__0_i_2__0
       (.I0(n22__1_n_0),
        .I1(B),
        .I2(n22__0_n_0),
        .I3(n22_n_0),
        .O(n14_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h37)) 
    n14_carry__0_i_3
       (.I0(n22__0_n_0),
        .I1(B),
        .I2(n22_n_0),
        .O(n14_carry__0_i_3_n_0));
  LUT4 #(
    .INIT(16'h4FDF)) 
    n14_carry__0_i_4__0
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(B),
        .I3(n22_n_0),
        .O(n14_carry__0_i_4__0_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n14_carry_i_10__0
       (.I0(n22__4_n_0),
        .I1(n22__2_n_0),
        .I2(B),
        .I3(n22__3_n_0),
        .I4(n22__1_n_0),
        .O(n14_carry_i_10__0_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n14_carry_i_11__0
       (.I0(n22__5_n_0),
        .I1(n22__3_n_0),
        .I2(B),
        .I3(n22__4_n_0),
        .I4(n22__2_n_0),
        .O(n14_carry_i_11__0_n_0));
  LUT5 #(
    .INIT(32'h66009600)) 
    n14_carry_i_12__0
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__5_n_0),
        .I3(B),
        .I4(n22__6_n_0),
        .O(n14_carry_i_12__0_n_0));
  LUT4 #(
    .INIT(16'h9060)) 
    n14_carry_i_13
       (.I0(n22__6_n_0),
        .I1(n22__5_n_0),
        .I2(B),
        .I3(n22__4_n_0),
        .O(n14_carry_i_13_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n14_carry_i_14
       (.I0(n22__5_n_0),
        .I1(B),
        .I2(n22__6_n_0),
        .O(n14_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14_carry_i_15
       (.I0(B),
        .I1(n22__6_n_0),
        .O(n14_carry_i_15_n_0));
  (* HLUTNM = "lutpair106" *) 
  LUT4 #(
    .INIT(16'hC880)) 
    n14_carry_i_1__0
       (.I0(n22__2_n_0),
        .I1(B),
        .I2(n22__1_n_0),
        .I3(n22__0_n_0),
        .O(n14_carry_i_1__0_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n14_carry_i_2__0
       (.I0(n22__3_n_0),
        .I1(B),
        .I2(n22__2_n_0),
        .I3(n22__1_n_0),
        .O(n14_carry_i_2__0_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n14_carry_i_3__0
       (.I0(n22__4_n_0),
        .I1(B),
        .I2(n22__3_n_0),
        .I3(n22__2_n_0),
        .O(n14_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n14_carry_i_4__0
       (.I0(n22__5_n_0),
        .I1(B),
        .I2(n22__4_n_0),
        .I3(n22__3_n_0),
        .O(n14_carry_i_4__0_n_0));
  LUT4 #(
    .INIT(16'h8448)) 
    n14_carry_i_5__0
       (.I0(n22__4_n_0),
        .I1(B),
        .I2(n22__5_n_0),
        .I3(n22__3_n_0),
        .O(n14_carry_i_5__0_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n14_carry_i_6__0
       (.I0(n22__5_n_0),
        .I1(B),
        .I2(n22__6_n_0),
        .O(n14_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14_carry_i_7
       (.I0(B),
        .I1(n22__5_n_0),
        .O(n14_carry_i_7_n_0));
  LUT5 #(
    .INIT(32'h95656595)) 
    n14_carry_i_8
       (.I0(n14_carry_i_1__0_n_0),
        .I1(n22__0_n_0),
        .I2(B),
        .I3(n22__1_n_0),
        .I4(n22_n_0),
        .O(n14_carry_i_8_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n14_carry_i_9__0
       (.I0(n22__3_n_0),
        .I1(n22__1_n_0),
        .I2(B),
        .I3(n22__2_n_0),
        .I4(n22__0_n_0),
        .O(n14_carry_i_9__0_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[0]),
        .Q(\n16_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[1]),
        .Q(\n16_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[2]),
        .Q(\n16_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[3]),
        .Q(\n16_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[4]),
        .Q(\n16_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[5]),
        .Q(\n16_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[6]),
        .Q(\n16_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[7]),
        .Q(\n16_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[0]),
        .Q(\n1_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[10]),
        .Q(n2[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[11]),
        .Q(n2[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[12]),
        .Q(n2[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[13]),
        .Q(n2[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[14]),
        .Q(n2[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[15]),
        .Q(n2[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[1]),
        .Q(\n1_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[2]),
        .Q(\n1_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[3]),
        .Q(\n1_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[4]),
        .Q(\n1_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[5]),
        .Q(\n1_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[6]),
        .Q(\n1_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[7]),
        .Q(\n1_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[8]),
        .Q(n2[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i2[9]),
        .Q(n2[1]),
        .R(rst_i));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_2 
       (.I0(\n16_reg_n_0_[7] ),
        .O(\n21[7]_i_2_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_3 
       (.I0(\n16_reg_n_0_[6] ),
        .O(\n21[7]_i_3_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_4 
       (.I0(\n16_reg_n_0_[5] ),
        .O(\n21[7]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_5 
       (.I0(\n16_reg_n_0_[4] ),
        .O(\n21[7]_i_5_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_6 
       (.I0(\n16_reg_n_0_[3] ),
        .O(\n21[7]_i_6_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_7 
       (.I0(\n16_reg_n_0_[2] ),
        .O(\n21[7]_i_7_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_8 
       (.I0(\n16_reg_n_0_[1] ),
        .O(\n21[7]_i_8_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_9 
       (.I0(\n16_reg_n_0_[0] ),
        .O(\n21[7]_i_9_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[0]),
        .Q(n21[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[1]),
        .Q(n21[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[2]),
        .Q(n21[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[3]),
        .Q(n21[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[4]),
        .Q(n21[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[5]),
        .Q(n21[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[6]),
        .Q(n21[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[7]),
        .Q(n21[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n21_reg[7]_i_1__2 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\NLW_n21_reg[7]_i_1__2_CO_UNCONNECTED [7],\n21_reg[7]_i_1__2_n_1 ,\n21_reg[7]_i_1__2_n_2 ,\n21_reg[7]_i_1__2_n_3 ,\n21_reg[7]_i_1__2_n_4 ,\n21_reg[7]_i_1__2_n_5 ,\n21_reg[7]_i_1__2_n_6 ,\n21_reg[7]_i_1__2_n_7 }),
        .DI({1'b0,\n16_reg_n_0_[6] ,\n16_reg_n_0_[5] ,\n16_reg_n_0_[4] ,\n16_reg_n_0_[3] ,\n16_reg_n_0_[2] ,\n16_reg_n_0_[1] ,\n16_reg_n_0_[0] }),
        .O(n202_out),
        .S({\n21[7]_i_2_n_0 ,\n21[7]_i_3_n_0 ,\n21[7]_i_4_n_0 ,\n21[7]_i_5_n_0 ,\n21[7]_i_6_n_0 ,\n21[7]_i_7_n_0 ,\n21[7]_i_8_n_0 ,\n21[7]_i_9_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    n22
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[15]),
        .Q(n22_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__0
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[14]),
        .Q(n22__0_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__1
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[13]),
        .Q(n22__1_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__2
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[12]),
        .Q(n22__2_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__3
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[11]),
        .Q(n22__3_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__4
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[10]),
        .Q(n22__4_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__5
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[9]),
        .Q(n22__5_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__6
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[8]),
        .Q(n22__6_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__17_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__17_carry_n_0,n25__17_carry_n_1,n25__17_carry_n_2,n25__17_carry_n_3,n25__17_carry_n_4,n25__17_carry_n_5,n25__17_carry_n_6,n25__17_carry_n_7}),
        .DI({n25_carry_i_1__0_n_0,n25__17_carry_i_1__0_n_0,n25__17_carry_i_2__0_n_0,n25__17_carry_i_3__0_n_0,n25__17_carry_i_4__0_n_0,n25__17_carry_i_5__0_n_0,n25__17_carry_i_6_n_0,1'b0}),
        .O({n25__17_carry_n_8,n25__17_carry_n_9,n25__17_carry_n_10,n25__17_carry_n_11,n25__17_carry_n_12,n25__17_carry_n_13,n25__17_carry_n_14,NLW_n25__17_carry_O_UNCONNECTED[0]}),
        .S({n25__17_carry_i_7_n_0,n25__17_carry_i_8__0_n_0,n25__17_carry_i_9_n_0,n25__17_carry_i_10__0_n_0,n25__17_carry_i_11_n_0,n25__17_carry_i_12_n_0,n25__17_carry_i_13_n_0,n25__17_carry_i_14_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__17_carry__0
       (.CI(n25__17_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__17_carry__0_CO_UNCONNECTED[7:3],n25__17_carry__0_n_5,NLW_n25__17_carry__0_CO_UNCONNECTED[1],n25__17_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25__17_carry__0_i_1_n_0,n25__17_carry__0_i_2__0_n_0}),
        .O({NLW_n25__17_carry__0_O_UNCONNECTED[7:2],n25__17_carry__0_n_14,n25__17_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n25__17_carry__0_i_3_n_0,n25__17_carry__0_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h40)) 
    n25__17_carry__0_i_1
       (.I0(n4[7]),
        .I1(B),
        .I2(n4[6]),
        .O(n25__17_carry__0_i_1_n_0));
  LUT4 #(
    .INIT(16'h80C8)) 
    n25__17_carry__0_i_2__0
       (.I0(n4[5]),
        .I1(B),
        .I2(n4[6]),
        .I3(n4[7]),
        .O(n25__17_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h37)) 
    n25__17_carry__0_i_3
       (.I0(n4[6]),
        .I1(B),
        .I2(n4[7]),
        .O(n25__17_carry__0_i_3_n_0));
  LUT4 #(
    .INIT(16'h4FDF)) 
    n25__17_carry__0_i_4__0
       (.I0(n4[5]),
        .I1(n4[6]),
        .I2(B),
        .I3(n4[7]),
        .O(n25__17_carry__0_i_4__0_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n25__17_carry_i_10__0
       (.I0(n4[1]),
        .I1(n4[3]),
        .I2(B),
        .I3(n4[2]),
        .I4(n4[4]),
        .O(n25__17_carry_i_10__0_n_0));
  LUT5 #(
    .INIT(32'h66009600)) 
    n25__17_carry_i_11
       (.I0(n4[2]),
        .I1(n4[3]),
        .I2(n4[1]),
        .I3(B),
        .I4(n4[0]),
        .O(n25__17_carry_i_11_n_0));
  LUT4 #(
    .INIT(16'h9060)) 
    n25__17_carry_i_12
       (.I0(n4[0]),
        .I1(n4[1]),
        .I2(B),
        .I3(n4[2]),
        .O(n25__17_carry_i_12_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n25__17_carry_i_13
       (.I0(n4[1]),
        .I1(B),
        .I2(n4[0]),
        .O(n25__17_carry_i_13_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__17_carry_i_14
       (.I0(B),
        .I1(n4[0]),
        .O(n25__17_carry_i_14_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n25__17_carry_i_1__0
       (.I0(n4[3]),
        .I1(B),
        .I2(n4[4]),
        .I3(n4[5]),
        .O(n25__17_carry_i_1__0_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n25__17_carry_i_2__0
       (.I0(n4[2]),
        .I1(B),
        .I2(n4[3]),
        .I3(n4[4]),
        .O(n25__17_carry_i_2__0_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n25__17_carry_i_3__0
       (.I0(n4[1]),
        .I1(B),
        .I2(n4[2]),
        .I3(n4[3]),
        .O(n25__17_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h8448)) 
    n25__17_carry_i_4__0
       (.I0(n4[2]),
        .I1(B),
        .I2(n4[1]),
        .I3(n4[3]),
        .O(n25__17_carry_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n25__17_carry_i_5__0
       (.I0(n4[1]),
        .I1(B),
        .I2(n4[0]),
        .O(n25__17_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__17_carry_i_6
       (.I0(B),
        .I1(n4[1]),
        .O(n25__17_carry_i_6_n_0));
  LUT5 #(
    .INIT(32'h95656595)) 
    n25__17_carry_i_7
       (.I0(n25_carry_i_1__0_n_0),
        .I1(n4[6]),
        .I2(B),
        .I3(n4[5]),
        .I4(n4[7]),
        .O(n25__17_carry_i_7_n_0));
  (* HLUTNM = "lutpair104" *) 
  LUT5 #(
    .INIT(32'h4C8004C8)) 
    n25__17_carry_i_8__0
       (.I0(n4[4]),
        .I1(B),
        .I2(n4[5]),
        .I3(n4[6]),
        .I4(n4[3]),
        .O(n25__17_carry_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n25__17_carry_i_9
       (.I0(n4[2]),
        .I1(n4[4]),
        .I2(B),
        .I3(n4[3]),
        .I4(n4[5]),
        .O(n25__17_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__47_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__47_carry_CO_UNCONNECTED[7],n25__47_carry_n_1,n25__47_carry_n_2,n25__47_carry_n_3,n25__47_carry_n_4,n25__47_carry_n_5,n25__47_carry_n_6,n25__47_carry_n_7}),
        .DI({1'b0,n25__47_carry_i_1__0_n_0,n25__47_carry_i_2__0_n_0,n25__47_carry_i_3_n_0,n25__47_carry_i_4_n_0,1'b1,1'b0,1'b1}),
        .O({n25__47_carry_n_8,n25__47_carry_n_9,n25__47_carry_n_10,n25__47_carry_n_11,n25__47_carry_n_12,n25__47_carry_n_13,n25__47_carry_n_14,n25__47_carry_n_15}),
        .S({n25__47_carry_i_5_n_0,n25__47_carry_i_6__0_n_0,n25__47_carry_i_7_n_0,n25__47_carry_i_8_n_0,n25__47_carry_i_9_n_0,n25__47_carry_i_10_n_0,n25__47_carry_i_11_n_0,n25__47_carry_i_12_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n25__47_carry_i_10
       (.I0(B),
        .I1(n4[3]),
        .O(n25__47_carry_i_10_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__47_carry_i_11
       (.I0(B),
        .I1(n4[2]),
        .O(n25__47_carry_i_11_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n25__47_carry_i_12
       (.I0(n4[1]),
        .I1(B),
        .O(n25__47_carry_i_12_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__47_carry_i_1__0
       (.I0(B),
        .I1(n4[6]),
        .O(n25__47_carry_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__47_carry_i_2__0
       (.I0(B),
        .I1(n4[5]),
        .O(n25__47_carry_i_2__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__47_carry_i_3
       (.I0(B),
        .I1(n4[4]),
        .O(n25__47_carry_i_3_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__47_carry_i_4
       (.I0(B),
        .I1(n4[3]),
        .O(n25__47_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n25__47_carry_i_5
       (.I0(n4[7]),
        .I1(B),
        .O(n25__47_carry_i_5_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n25__47_carry_i_6__0
       (.I0(n4[6]),
        .I1(B),
        .I2(n4[7]),
        .O(n25__47_carry_i_6__0_n_0));
  LUT3 #(
    .INIT(8'hB7)) 
    n25__47_carry_i_7
       (.I0(n4[5]),
        .I1(B),
        .I2(n4[6]),
        .O(n25__47_carry_i_7_n_0));
  LUT3 #(
    .INIT(8'hB7)) 
    n25__47_carry_i_8
       (.I0(n4[4]),
        .I1(B),
        .I2(n4[5]),
        .O(n25__47_carry_i_8_n_0));
  LUT3 #(
    .INIT(8'hB7)) 
    n25__47_carry_i_9
       (.I0(n4[3]),
        .I1(B),
        .I2(n4[4]),
        .O(n25__47_carry_i_9_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__67_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__67_carry_n_0,n25__67_carry_n_1,n25__67_carry_n_2,n25__67_carry_n_3,n25__67_carry_n_4,n25__67_carry_n_5,n25__67_carry_n_6,n25__67_carry_n_7}),
        .DI({n25__67_carry_i_1__0_n_0,n25__67_carry_i_2__0_n_0,n25__67_carry_i_3__0_n_0,n25__67_carry_i_4__0_n_0,n25__67_carry_i_5__0_n_0,n25__67_carry_i_6__0_n_0,n25__67_carry_i_7__0_n_0,1'b0}),
        .O({n26[3:0],NLW_n25__67_carry_O_UNCONNECTED[3:0]}),
        .S({n25__67_carry_i_8__0_n_0,n25__67_carry_i_9__0_n_0,n25__67_carry_i_10__0_n_0,n25__67_carry_i_11__0_n_0,n25__67_carry_i_12__0_n_0,n25__67_carry_i_13__0_n_0,n25__67_carry_i_14__0_n_0,n25__67_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__67_carry__0
       (.CI(n25__67_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__67_carry__0_CO_UNCONNECTED[7:3],n25__67_carry__0_n_5,n25__67_carry__0_n_6,n25__67_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n25__67_carry__0_i_1__0_n_0,n25__67_carry__0_i_2__0_n_0,n25__67_carry__0_i_3__0_n_0}),
        .O({NLW_n25__67_carry__0_O_UNCONNECTED[7:4],n26[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n25__67_carry__0_i_4__0_n_0,n25__67_carry__0_i_5__0_n_0,n25__67_carry__0_i_6__0_n_0,n25__67_carry__0_i_7__0_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry__0_i_1__0
       (.I0(n25__17_carry__0_n_14),
        .I1(n25__47_carry_n_10),
        .O(n25__67_carry__0_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry__0_i_2__0
       (.I0(n25__17_carry__0_n_15),
        .I1(n25__47_carry_n_11),
        .O(n25__67_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25__67_carry__0_i_3__0
       (.I0(n25__47_carry_n_12),
        .I1(n25__17_carry_n_8),
        .I2(n25_carry__0_n_5),
        .O(n25__67_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n25__67_carry__0_i_4__0
       (.I0(n25__17_carry__0_n_5),
        .I1(n25__47_carry_n_9),
        .I2(n25__47_carry_n_8),
        .O(n25__67_carry__0_i_4__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__67_carry__0_i_5__0
       (.I0(n25__17_carry__0_n_14),
        .I1(n25__47_carry_n_10),
        .I2(n25__47_carry_n_9),
        .I3(n25__17_carry__0_n_5),
        .O(n25__67_carry__0_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__67_carry__0_i_6__0
       (.I0(n25__17_carry__0_n_15),
        .I1(n25__47_carry_n_11),
        .I2(n25__47_carry_n_10),
        .I3(n25__17_carry__0_n_14),
        .O(n25__67_carry__0_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n25__67_carry__0_i_7__0
       (.I0(n25_carry__0_n_5),
        .I1(n25__17_carry_n_8),
        .I2(n25__47_carry_n_12),
        .I3(n25__47_carry_n_11),
        .I4(n25__17_carry__0_n_15),
        .O(n25__67_carry__0_i_7__0_n_0));
  (* HLUTNM = "lutpair66" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__67_carry_i_10__0
       (.I0(n25__47_carry_n_14),
        .I1(n25__17_carry_n_10),
        .I2(n25_carry__0_n_15),
        .I3(n25__67_carry_i_3__0_n_0),
        .O(n25__67_carry_i_10__0_n_0));
  (* HLUTNM = "lutpair65" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__67_carry_i_11__0
       (.I0(n25__47_carry_n_15),
        .I1(n25__17_carry_n_11),
        .I2(n25_carry_n_8),
        .I3(n25__67_carry_i_4__0_n_0),
        .O(n25__67_carry_i_11__0_n_0));
  (* HLUTNM = "lutpair64" *) 
  LUT5 #(
    .INIT(32'h78878778)) 
    n25__67_carry_i_12__0
       (.I0(B),
        .I1(n4[0]),
        .I2(n25__17_carry_n_12),
        .I3(n25_carry_n_9),
        .I4(n25__67_carry_i_5__0_n_0),
        .O(n25__67_carry_i_12__0_n_0));
  (* HLUTNM = "lutpair105" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n25__67_carry_i_13__0
       (.I0(n25__17_carry_n_13),
        .I1(n25_carry_n_10),
        .I2(n25_carry_n_11),
        .I3(n25__17_carry_n_14),
        .O(n25__67_carry_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__67_carry_i_14__0
       (.I0(n25_carry_n_12),
        .I1(n25_carry_n_15),
        .I2(n25__17_carry_n_14),
        .I3(n25_carry_n_11),
        .O(n25__67_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n25__67_carry_i_15__0
       (.I0(n25_carry_n_12),
        .I1(n25_carry_n_15),
        .O(n25__67_carry_i_15__0_n_0));
  (* HLUTNM = "lutpair67" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__67_carry_i_1__0
       (.I0(n25__47_carry_n_13),
        .I1(n25__17_carry_n_9),
        .I2(n25_carry__0_n_14),
        .O(n25__67_carry_i_1__0_n_0));
  (* HLUTNM = "lutpair66" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__67_carry_i_2__0
       (.I0(n25__47_carry_n_14),
        .I1(n25__17_carry_n_10),
        .I2(n25_carry__0_n_15),
        .O(n25__67_carry_i_2__0_n_0));
  (* HLUTNM = "lutpair65" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__67_carry_i_3__0
       (.I0(n25__47_carry_n_15),
        .I1(n25__17_carry_n_11),
        .I2(n25_carry_n_8),
        .O(n25__67_carry_i_3__0_n_0));
  (* HLUTNM = "lutpair64" *) 
  LUT4 #(
    .INIT(16'hF880)) 
    n25__67_carry_i_4__0
       (.I0(B),
        .I1(n4[0]),
        .I2(n25__17_carry_n_12),
        .I3(n25_carry_n_9),
        .O(n25__67_carry_i_4__0_n_0));
  (* HLUTNM = "lutpair105" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry_i_5__0
       (.I0(n25__17_carry_n_13),
        .I1(n25_carry_n_10),
        .O(n25__67_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry_i_6__0
       (.I0(n25_carry_n_11),
        .I1(n25__17_carry_n_14),
        .O(n25__67_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry_i_7__0
       (.I0(n25_carry_n_12),
        .I1(n25_carry_n_15),
        .O(n25__67_carry_i_7__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n25__67_carry_i_8__0
       (.I0(n25__67_carry_i_1__0_n_0),
        .I1(n25__17_carry_n_8),
        .I2(n25__47_carry_n_12),
        .I3(n25_carry__0_n_5),
        .O(n25__67_carry_i_8__0_n_0));
  (* HLUTNM = "lutpair67" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__67_carry_i_9__0
       (.I0(n25__47_carry_n_13),
        .I1(n25__17_carry_n_9),
        .I2(n25_carry__0_n_14),
        .I3(n25__67_carry_i_2__0_n_0),
        .O(n25__67_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25_carry_n_0,n25_carry_n_1,n25_carry_n_2,n25_carry_n_3,n25_carry_n_4,n25_carry_n_5,n25_carry_n_6,n25_carry_n_7}),
        .DI({n25_carry_i_1__0_n_0,n25_carry_i_2__0_n_0,n25_carry_i_3__0_n_0,n25_carry_i_4__0_n_0,n25_carry_i_5__0_n_0,n25_carry_i_6__0_n_0,n25_carry_i_7_n_0,1'b0}),
        .O({n25_carry_n_8,n25_carry_n_9,n25_carry_n_10,n25_carry_n_11,n25_carry_n_12,NLW_n25_carry_O_UNCONNECTED[2:1],n25_carry_n_15}),
        .S({n25_carry_i_8_n_0,n25_carry_i_9__0_n_0,n25_carry_i_10__0_n_0,n25_carry_i_11__0_n_0,n25_carry_i_12__0_n_0,n25_carry_i_13_n_0,n25_carry_i_14_n_0,n25_carry_i_15_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25_carry__0
       (.CI(n25_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25_carry__0_CO_UNCONNECTED[7:3],n25_carry__0_n_5,NLW_n25_carry__0_CO_UNCONNECTED[1],n25_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25_carry__0_i_1__0_n_0,n25_carry__0_i_2__0_n_0}),
        .O({NLW_n25_carry__0_O_UNCONNECTED[7:2],n25_carry__0_n_14,n25_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n25_carry__0_i_3_n_0,n25_carry__0_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h40)) 
    n25_carry__0_i_1__0
       (.I0(n4[7]),
        .I1(B),
        .I2(n4[6]),
        .O(n25_carry__0_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h80C8)) 
    n25_carry__0_i_2__0
       (.I0(n4[5]),
        .I1(B),
        .I2(n4[6]),
        .I3(n4[7]),
        .O(n25_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h37)) 
    n25_carry__0_i_3
       (.I0(n4[6]),
        .I1(B),
        .I2(n4[7]),
        .O(n25_carry__0_i_3_n_0));
  LUT4 #(
    .INIT(16'h4FDF)) 
    n25_carry__0_i_4__0
       (.I0(n4[5]),
        .I1(n4[6]),
        .I2(B),
        .I3(n4[7]),
        .O(n25_carry__0_i_4__0_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n25_carry_i_10__0
       (.I0(n4[2]),
        .I1(n4[4]),
        .I2(B),
        .I3(n4[3]),
        .I4(n4[5]),
        .O(n25_carry_i_10__0_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n25_carry_i_11__0
       (.I0(n4[1]),
        .I1(n4[3]),
        .I2(B),
        .I3(n4[2]),
        .I4(n4[4]),
        .O(n25_carry_i_11__0_n_0));
  LUT5 #(
    .INIT(32'h66009600)) 
    n25_carry_i_12__0
       (.I0(n4[2]),
        .I1(n4[3]),
        .I2(n4[1]),
        .I3(B),
        .I4(n4[0]),
        .O(n25_carry_i_12__0_n_0));
  LUT4 #(
    .INIT(16'h9060)) 
    n25_carry_i_13
       (.I0(n4[0]),
        .I1(n4[1]),
        .I2(B),
        .I3(n4[2]),
        .O(n25_carry_i_13_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n25_carry_i_14
       (.I0(n4[1]),
        .I1(B),
        .I2(n4[0]),
        .O(n25_carry_i_14_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25_carry_i_15
       (.I0(B),
        .I1(n4[0]),
        .O(n25_carry_i_15_n_0));
  (* HLUTNM = "lutpair104" *) 
  LUT4 #(
    .INIT(16'hC880)) 
    n25_carry_i_1__0
       (.I0(n4[4]),
        .I1(B),
        .I2(n4[5]),
        .I3(n4[6]),
        .O(n25_carry_i_1__0_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n25_carry_i_2__0
       (.I0(n4[3]),
        .I1(B),
        .I2(n4[4]),
        .I3(n4[5]),
        .O(n25_carry_i_2__0_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n25_carry_i_3__0
       (.I0(n4[2]),
        .I1(B),
        .I2(n4[3]),
        .I3(n4[4]),
        .O(n25_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n25_carry_i_4__0
       (.I0(n4[1]),
        .I1(B),
        .I2(n4[2]),
        .I3(n4[3]),
        .O(n25_carry_i_4__0_n_0));
  LUT4 #(
    .INIT(16'h8448)) 
    n25_carry_i_5__0
       (.I0(n4[2]),
        .I1(B),
        .I2(n4[1]),
        .I3(n4[3]),
        .O(n25_carry_i_5__0_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n25_carry_i_6__0
       (.I0(n4[1]),
        .I1(B),
        .I2(n4[0]),
        .O(n25_carry_i_6__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25_carry_i_7
       (.I0(B),
        .I1(n4[1]),
        .O(n25_carry_i_7_n_0));
  LUT5 #(
    .INIT(32'h95656595)) 
    n25_carry_i_8
       (.I0(n25_carry_i_1__0_n_0),
        .I1(n4[6]),
        .I2(B),
        .I3(n4[5]),
        .I4(n4[7]),
        .O(n25_carry_i_8_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n25_carry_i_9__0
       (.I0(n4[3]),
        .I1(n4[5]),
        .I2(B),
        .I3(n4[4]),
        .I4(n4[6]),
        .O(n25_carry_i_9__0_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[0]),
        .Q(n27[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[1]),
        .Q(n27[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[2]),
        .Q(n27[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[3]),
        .Q(n27[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[4]),
        .Q(n27[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[5]),
        .Q(n27[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[6]),
        .Q(n27[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[7]),
        .Q(n27[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[0]),
        .Q(n29[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[1]),
        .Q(n29[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[2]),
        .Q(n29[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[3]),
        .Q(n29[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[4]),
        .Q(n29[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[5]),
        .Q(n29[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[6]),
        .Q(n29[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[7]),
        .Q(n29[7]),
        .R(rst_i));
  LUT2 #(
    .INIT(4'h6)) 
    \n33[0]_i_1__6 
       (.I0(n29[0]),
        .I1(n10[0]),
        .O(n31[0]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[10]_i_1__6 
       (.I0(n21[2]),
        .I1(\n8_reg_n_0_[2] ),
        .I2(\n8_reg_n_0_[1] ),
        .I3(n21[1]),
        .I4(\n8_reg_n_0_[0] ),
        .I5(n21[0]),
        .O(\n33[10]_i_1__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[11]_i_1__6 
       (.I0(n21[3]),
        .I1(\n8_reg_n_0_[3] ),
        .I2(\n33[12]_i_2__6_n_0 ),
        .O(\n33[11]_i_1__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[12]_i_1__6 
       (.I0(n21[4]),
        .I1(\n8_reg_n_0_[4] ),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[3]),
        .I4(\n33[12]_i_2__6_n_0 ),
        .O(\n33[12]_i_1__6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[12]_i_2__6 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n33[12]_i_2__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[13]_i_1__6 
       (.I0(n21[5]),
        .I1(\n8_reg_n_0_[5] ),
        .I2(\n33[14]_i_2__6_n_0 ),
        .O(\n33[13]_i_1__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[14]_i_1__6 
       (.I0(n21[6]),
        .I1(\n8_reg_n_0_[6] ),
        .I2(\n8_reg_n_0_[5] ),
        .I3(n21[5]),
        .I4(\n33[14]_i_2__6_n_0 ),
        .O(\n33[14]_i_1__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[14]_i_2__6 
       (.I0(\n33[12]_i_2__6_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n33[14]_i_2__6_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[15]_i_1__6 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n33[15]_i_2__6_n_0 ),
        .O(n30));
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[15]_i_2__6 
       (.I0(\n33[14]_i_2__6_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n33[15]_i_2__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[1]_i_1__6 
       (.I0(n29[1]),
        .I1(n10[1]),
        .I2(n10[0]),
        .I3(n29[0]),
        .O(n31[1]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[2]_i_1__6 
       (.I0(n29[2]),
        .I1(n10[2]),
        .I2(n10[1]),
        .I3(n29[1]),
        .I4(n10[0]),
        .I5(n29[0]),
        .O(\n33[2]_i_1__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[3]_i_1__6 
       (.I0(n29[3]),
        .I1(n10[3]),
        .I2(\n33[4]_i_2__6_n_0 ),
        .O(\n33[3]_i_1__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[4]_i_1__6 
       (.I0(n29[4]),
        .I1(n10[4]),
        .I2(n10[3]),
        .I3(n29[3]),
        .I4(\n33[4]_i_2__6_n_0 ),
        .O(\n33[4]_i_1__6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[4]_i_2__6 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n33[4]_i_2__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[5]_i_1__6 
       (.I0(n29[5]),
        .I1(n10[5]),
        .I2(\n33[6]_i_2__6_n_0 ),
        .O(\n33[5]_i_1__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[6]_i_1__6 
       (.I0(n29[6]),
        .I1(n10[6]),
        .I2(n10[5]),
        .I3(n29[5]),
        .I4(\n33[6]_i_2__6_n_0 ),
        .O(\n33[6]_i_1__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[6]_i_2__6 
       (.I0(\n33[4]_i_2__6_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n33[6]_i_2__6_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[7]_i_1__6 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n33[7]_i_2__6_n_0 ),
        .O(n31[7]));
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[7]_i_2__6 
       (.I0(\n33[6]_i_2__6_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n33[7]_i_2__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[9]_i_1__6 
       (.I0(n21[1]),
        .I1(\n8_reg_n_0_[1] ),
        .I2(\n8_reg_n_0_[0] ),
        .I3(n21[0]),
        .O(\n33[9]_i_1__6_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[0]),
        .Q(i1[15]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[10]_i_1__6_n_0 ),
        .Q(i1[24]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[11]_i_1__6_n_0 ),
        .Q(i1[25]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[12]_i_1__6_n_0 ),
        .Q(i1[26]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[13]_i_1__6_n_0 ),
        .Q(i1[27]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[14]_i_1__6_n_0 ),
        .Q(i1[28]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n30),
        .Q(i1[29]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[1]),
        .Q(i1[16]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[2]_i_1__6_n_0 ),
        .Q(i1[17]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[3]_i_1__6_n_0 ),
        .Q(i1[18]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[4]_i_1__6_n_0 ),
        .Q(i1[19]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[5]_i_1__6_n_0 ),
        .Q(i1[20]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[6]_i_1__6_n_0 ),
        .Q(i1[21]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[7]),
        .Q(i1[22]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[9]_i_1__6_n_0 ),
        .Q(i1[23]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[10]_i_1__6 
       (.I0(\n8_reg_n_0_[1] ),
        .I1(n21[1]),
        .I2(n21[0]),
        .I3(\n8_reg_n_0_[0] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(n341_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[11]_i_1__6 
       (.I0(\n37[12]_i_2__6_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .O(n341_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[12]_i_1__6 
       (.I0(\n8_reg_n_0_[3] ),
        .I1(n21[3]),
        .I2(\n37[12]_i_2__6_n_0 ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(n341_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[12]_i_2__6 
       (.I0(\n8_reg_n_0_[0] ),
        .I1(n21[0]),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n37[12]_i_2__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[13]_i_1__6 
       (.I0(\n37[14]_i_2__6_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(n341_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[14]_i_1__6 
       (.I0(\n8_reg_n_0_[5] ),
        .I1(n21[5]),
        .I2(\n37[14]_i_2__6_n_0 ),
        .I3(n21[6]),
        .I4(\n8_reg_n_0_[6] ),
        .O(n341_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[14]_i_2__6 
       (.I0(\n37[12]_i_2__6_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n37[14]_i_2__6_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[15]_i_1__6 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n37[15]_i_2__6_n_0 ),
        .O(n341_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[15]_i_2__6 
       (.I0(\n37[14]_i_2__6_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n37[15]_i_2__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[1]_i_1__6 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .O(n350_out[1]));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[2]_i_1__6 
       (.I0(n10[1]),
        .I1(n29[1]),
        .I2(n29[0]),
        .I3(n10[0]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(n350_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[3]_i_1__6 
       (.I0(\n37[4]_i_2__6_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .O(n350_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[4]_i_1__6 
       (.I0(n10[3]),
        .I1(n29[3]),
        .I2(\n37[4]_i_2__6_n_0 ),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(n350_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[4]_i_2__6 
       (.I0(n10[0]),
        .I1(n29[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n37[4]_i_2__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[5]_i_1__6 
       (.I0(\n37[6]_i_2__6_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(n350_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[6]_i_1__6 
       (.I0(n10[5]),
        .I1(n29[5]),
        .I2(\n37[6]_i_2__6_n_0 ),
        .I3(n29[6]),
        .I4(n10[6]),
        .O(n350_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[6]_i_2__6 
       (.I0(\n37[4]_i_2__6_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n37[6]_i_2__6_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[7]_i_1__6 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n37[7]_i_2__6_n_0 ),
        .O(n350_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[7]_i_2__6 
       (.I0(\n37[6]_i_2__6_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n37[7]_i_2__6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n37[8]_i_1__3 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .O(n341_out[0]));
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[9]_i_1__6 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .O(n341_out[1]));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[2]),
        .Q(i1[9]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[3]),
        .Q(i1[10]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[4]),
        .Q(i1[11]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[5]),
        .Q(i1[12]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[6]),
        .Q(i1[13]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[7]),
        .Q(i1[14]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[1]),
        .Q(i1[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[2]),
        .Q(i1[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[3]),
        .Q(i1[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[4]),
        .Q(i1[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[5]),
        .Q(i1[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[6]),
        .Q(i1[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[7]),
        .Q(i1[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[0]),
        .Q(i1[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[1]),
        .Q(i1[8]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[0]),
        .Q(n4[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[1]),
        .Q(n4[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[2]),
        .Q(n4[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[3]),
        .Q(n4[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[4]),
        .Q(n4[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[5]),
        .Q(n4[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[6]),
        .Q(n4[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(i3[7]),
        .Q(n4[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[0]),
        .Q(\n7_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[1]),
        .Q(\n7_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[2]),
        .Q(\n7_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[3]),
        .Q(\n7_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[4]),
        .Q(\n7_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[5]),
        .Q(\n7_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[6]),
        .Q(\n7_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[7]),
        .Q(\n7_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[0] ),
        .Q(\n8_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[1] ),
        .Q(\n8_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[2] ),
        .Q(\n8_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[3] ),
        .Q(\n8_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[4] ),
        .Q(\n8_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[5] ),
        .Q(\n8_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[6] ),
        .Q(\n8_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[7] ),
        .Q(\n8_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[0] ),
        .Q(\n9_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[1] ),
        .Q(\n9_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[2] ),
        .Q(\n9_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[3] ),
        .Q(\n9_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[4] ),
        .Q(\n9_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[5] ),
        .Q(\n9_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[6] ),
        .Q(\n9_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[7] ),
        .Q(\n9_reg_n_0_[7] ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_37" *) 
module switch_elements_cf_fft_512_8_37_22
   (i1,
    enable_i,
    clk_i,
    rst_i,
    n22_0,
    \n1_reg[15]_0 ,
    \n4_reg[7]_0 );
  output [29:0]i1;
  input [0:0]enable_i;
  input clk_i;
  input rst_i;
  input [7:0]n22_0;
  input [15:0]\n1_reg[15]_0 ;
  input [7:0]\n4_reg[7]_0 ;

  wire [6:6]B;
  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [7:0]n10;
  wire n14__21_carry__0_i_1__0_n_0;
  wire n14__21_carry__0_i_2__1_n_0;
  wire n14__21_carry__0_i_3__0_n_0;
  wire n14__21_carry__0_i_4__1_n_0;
  wire n14__21_carry__0_n_14;
  wire n14__21_carry__0_n_15;
  wire n14__21_carry__0_n_5;
  wire n14__21_carry__0_n_7;
  wire n14__21_carry_i_10__1_n_0;
  wire n14__21_carry_i_11__0_n_0;
  wire n14__21_carry_i_12__0_n_0;
  wire n14__21_carry_i_13__0_n_0;
  wire n14__21_carry_i_14__0_n_0;
  wire n14__21_carry_i_1__1_n_0;
  wire n14__21_carry_i_2__1_n_0;
  wire n14__21_carry_i_3__1_n_0;
  wire n14__21_carry_i_4__1_n_0;
  wire n14__21_carry_i_5__1_n_0;
  wire n14__21_carry_i_6__0_n_0;
  wire n14__21_carry_i_7__0_n_0;
  wire n14__21_carry_i_8__1_n_0;
  wire n14__21_carry_i_9__0_n_0;
  wire n14__21_carry_n_0;
  wire n14__21_carry_n_1;
  wire n14__21_carry_n_10;
  wire n14__21_carry_n_11;
  wire n14__21_carry_n_12;
  wire n14__21_carry_n_13;
  wire n14__21_carry_n_14;
  wire n14__21_carry_n_2;
  wire n14__21_carry_n_3;
  wire n14__21_carry_n_4;
  wire n14__21_carry_n_5;
  wire n14__21_carry_n_6;
  wire n14__21_carry_n_7;
  wire n14__21_carry_n_8;
  wire n14__21_carry_n_9;
  wire n14__47_carry_i_10__0_n_0;
  wire n14__47_carry_i_11__0_n_0;
  wire n14__47_carry_i_12__0_n_0;
  wire n14__47_carry_i_1__1_n_0;
  wire n14__47_carry_i_2__1_n_0;
  wire n14__47_carry_i_3__0_n_0;
  wire n14__47_carry_i_4__0_n_0;
  wire n14__47_carry_i_5__0_n_0;
  wire n14__47_carry_i_6__1_n_0;
  wire n14__47_carry_i_7__0_n_0;
  wire n14__47_carry_i_8__0_n_0;
  wire n14__47_carry_i_9__0_n_0;
  wire n14__47_carry_n_1;
  wire n14__47_carry_n_10;
  wire n14__47_carry_n_11;
  wire n14__47_carry_n_12;
  wire n14__47_carry_n_13;
  wire n14__47_carry_n_14;
  wire n14__47_carry_n_15;
  wire n14__47_carry_n_2;
  wire n14__47_carry_n_3;
  wire n14__47_carry_n_4;
  wire n14__47_carry_n_5;
  wire n14__47_carry_n_6;
  wire n14__47_carry_n_7;
  wire n14__47_carry_n_8;
  wire n14__47_carry_n_9;
  wire n14__67_carry__0_i_1__1_n_0;
  wire n14__67_carry__0_i_2__1_n_0;
  wire n14__67_carry__0_i_3__1_n_0;
  wire n14__67_carry__0_i_4__1_n_0;
  wire n14__67_carry__0_i_5__1_n_0;
  wire n14__67_carry__0_i_6__1_n_0;
  wire n14__67_carry__0_i_7__1_n_0;
  wire n14__67_carry__0_n_5;
  wire n14__67_carry__0_n_6;
  wire n14__67_carry__0_n_7;
  wire n14__67_carry_i_10__1_n_0;
  wire n14__67_carry_i_11__1_n_0;
  wire n14__67_carry_i_12__1_n_0;
  wire n14__67_carry_i_13__1_n_0;
  wire n14__67_carry_i_14__1_n_0;
  wire n14__67_carry_i_15__1_n_0;
  wire n14__67_carry_i_1__1_n_0;
  wire n14__67_carry_i_2__1_n_0;
  wire n14__67_carry_i_3__1_n_0;
  wire n14__67_carry_i_4__1_n_0;
  wire n14__67_carry_i_5__1_n_0;
  wire n14__67_carry_i_6__1_n_0;
  wire n14__67_carry_i_7__1_n_0;
  wire n14__67_carry_i_8__1_n_0;
  wire n14__67_carry_i_9__1_n_0;
  wire n14__67_carry_n_0;
  wire n14__67_carry_n_1;
  wire n14__67_carry_n_2;
  wire n14__67_carry_n_3;
  wire n14__67_carry_n_4;
  wire n14__67_carry_n_5;
  wire n14__67_carry_n_6;
  wire n14__67_carry_n_7;
  wire n14_carry__0_i_1__1_n_0;
  wire n14_carry__0_i_2__1_n_0;
  wire n14_carry__0_i_3__0_n_0;
  wire n14_carry__0_i_4__1_n_0;
  wire n14_carry__0_n_14;
  wire n14_carry__0_n_15;
  wire n14_carry__0_n_5;
  wire n14_carry__0_n_7;
  wire n14_carry_i_10__1_n_0;
  wire n14_carry_i_11__1_n_0;
  wire n14_carry_i_12__1_n_0;
  wire n14_carry_i_13__0_n_0;
  wire n14_carry_i_14__0_n_0;
  wire n14_carry_i_15__0_n_0;
  wire n14_carry_i_1__1_n_0;
  wire n14_carry_i_2__1_n_0;
  wire n14_carry_i_3__1_n_0;
  wire n14_carry_i_4__1_n_0;
  wire n14_carry_i_5__1_n_0;
  wire n14_carry_i_6__1_n_0;
  wire n14_carry_i_7__0_n_0;
  wire n14_carry_i_8__0_n_0;
  wire n14_carry_i_9__1_n_0;
  wire n14_carry_n_0;
  wire n14_carry_n_1;
  wire n14_carry_n_10;
  wire n14_carry_n_11;
  wire n14_carry_n_12;
  wire n14_carry_n_15;
  wire n14_carry_n_2;
  wire n14_carry_n_3;
  wire n14_carry_n_4;
  wire n14_carry_n_5;
  wire n14_carry_n_6;
  wire n14_carry_n_7;
  wire n14_carry_n_8;
  wire n14_carry_n_9;
  wire [7:0]n15;
  wire \n16_reg_n_0_[0] ;
  wire \n16_reg_n_0_[1] ;
  wire \n16_reg_n_0_[2] ;
  wire \n16_reg_n_0_[3] ;
  wire \n16_reg_n_0_[4] ;
  wire \n16_reg_n_0_[5] ;
  wire \n16_reg_n_0_[6] ;
  wire \n16_reg_n_0_[7] ;
  wire [15:0]\n1_reg[15]_0 ;
  wire \n1_reg_n_0_[0] ;
  wire \n1_reg_n_0_[1] ;
  wire \n1_reg_n_0_[2] ;
  wire \n1_reg_n_0_[3] ;
  wire \n1_reg_n_0_[4] ;
  wire \n1_reg_n_0_[5] ;
  wire \n1_reg_n_0_[6] ;
  wire \n1_reg_n_0_[7] ;
  wire [7:0]n202_out;
  wire [7:0]n21;
  wire \n21[7]_i_2_n_0 ;
  wire \n21[7]_i_3_n_0 ;
  wire \n21[7]_i_4_n_0 ;
  wire \n21[7]_i_5_n_0 ;
  wire \n21[7]_i_6_n_0 ;
  wire \n21[7]_i_7_n_0 ;
  wire \n21[7]_i_8_n_0 ;
  wire \n21[7]_i_9_n_0 ;
  wire \n21_reg[7]_i_1__3_n_1 ;
  wire \n21_reg[7]_i_1__3_n_2 ;
  wire \n21_reg[7]_i_1__3_n_3 ;
  wire \n21_reg[7]_i_1__3_n_4 ;
  wire \n21_reg[7]_i_1__3_n_5 ;
  wire \n21_reg[7]_i_1__3_n_6 ;
  wire \n21_reg[7]_i_1__3_n_7 ;
  wire [7:0]n22_0;
  wire n22__0_n_0;
  wire n22__1_n_0;
  wire n22__2_n_0;
  wire n22__3_n_0;
  wire n22__4_n_0;
  wire n22__5_n_0;
  wire n22__6_n_0;
  wire n22_n_0;
  wire n25__17_carry__0_i_1__0_n_0;
  wire n25__17_carry__0_i_2__1_n_0;
  wire n25__17_carry__0_i_3__0_n_0;
  wire n25__17_carry__0_i_4__1_n_0;
  wire n25__17_carry__0_n_14;
  wire n25__17_carry__0_n_15;
  wire n25__17_carry__0_n_5;
  wire n25__17_carry__0_n_7;
  wire n25__17_carry_i_10__1_n_0;
  wire n25__17_carry_i_11__0_n_0;
  wire n25__17_carry_i_12__0_n_0;
  wire n25__17_carry_i_13__0_n_0;
  wire n25__17_carry_i_14__0_n_0;
  wire n25__17_carry_i_1__1_n_0;
  wire n25__17_carry_i_2__1_n_0;
  wire n25__17_carry_i_3__1_n_0;
  wire n25__17_carry_i_4__1_n_0;
  wire n25__17_carry_i_5__1_n_0;
  wire n25__17_carry_i_6__0_n_0;
  wire n25__17_carry_i_7__0_n_0;
  wire n25__17_carry_i_8__1_n_0;
  wire n25__17_carry_i_9__0_n_0;
  wire n25__17_carry_n_0;
  wire n25__17_carry_n_1;
  wire n25__17_carry_n_10;
  wire n25__17_carry_n_11;
  wire n25__17_carry_n_12;
  wire n25__17_carry_n_13;
  wire n25__17_carry_n_14;
  wire n25__17_carry_n_2;
  wire n25__17_carry_n_3;
  wire n25__17_carry_n_4;
  wire n25__17_carry_n_5;
  wire n25__17_carry_n_6;
  wire n25__17_carry_n_7;
  wire n25__17_carry_n_8;
  wire n25__17_carry_n_9;
  wire n25__47_carry_i_10__0_n_0;
  wire n25__47_carry_i_11__0_n_0;
  wire n25__47_carry_i_12__0_n_0;
  wire n25__47_carry_i_1__1_n_0;
  wire n25__47_carry_i_2__1_n_0;
  wire n25__47_carry_i_3__0_n_0;
  wire n25__47_carry_i_4__0_n_0;
  wire n25__47_carry_i_5__0_n_0;
  wire n25__47_carry_i_6__1_n_0;
  wire n25__47_carry_i_7__0_n_0;
  wire n25__47_carry_i_8__0_n_0;
  wire n25__47_carry_i_9__0_n_0;
  wire n25__47_carry_n_1;
  wire n25__47_carry_n_10;
  wire n25__47_carry_n_11;
  wire n25__47_carry_n_12;
  wire n25__47_carry_n_13;
  wire n25__47_carry_n_14;
  wire n25__47_carry_n_15;
  wire n25__47_carry_n_2;
  wire n25__47_carry_n_3;
  wire n25__47_carry_n_4;
  wire n25__47_carry_n_5;
  wire n25__47_carry_n_6;
  wire n25__47_carry_n_7;
  wire n25__47_carry_n_8;
  wire n25__47_carry_n_9;
  wire n25__67_carry__0_i_1__1_n_0;
  wire n25__67_carry__0_i_2__1_n_0;
  wire n25__67_carry__0_i_3__1_n_0;
  wire n25__67_carry__0_i_4__1_n_0;
  wire n25__67_carry__0_i_5__1_n_0;
  wire n25__67_carry__0_i_6__1_n_0;
  wire n25__67_carry__0_i_7__1_n_0;
  wire n25__67_carry__0_n_5;
  wire n25__67_carry__0_n_6;
  wire n25__67_carry__0_n_7;
  wire n25__67_carry_i_10__1_n_0;
  wire n25__67_carry_i_11__1_n_0;
  wire n25__67_carry_i_12__1_n_0;
  wire n25__67_carry_i_13__1_n_0;
  wire n25__67_carry_i_14__1_n_0;
  wire n25__67_carry_i_15__1_n_0;
  wire n25__67_carry_i_1__1_n_0;
  wire n25__67_carry_i_2__1_n_0;
  wire n25__67_carry_i_3__1_n_0;
  wire n25__67_carry_i_4__1_n_0;
  wire n25__67_carry_i_5__1_n_0;
  wire n25__67_carry_i_6__1_n_0;
  wire n25__67_carry_i_7__1_n_0;
  wire n25__67_carry_i_8__1_n_0;
  wire n25__67_carry_i_9__1_n_0;
  wire n25__67_carry_n_0;
  wire n25__67_carry_n_1;
  wire n25__67_carry_n_2;
  wire n25__67_carry_n_3;
  wire n25__67_carry_n_4;
  wire n25__67_carry_n_5;
  wire n25__67_carry_n_6;
  wire n25__67_carry_n_7;
  wire n25_carry__0_i_1__1_n_0;
  wire n25_carry__0_i_2__1_n_0;
  wire n25_carry__0_i_3__0_n_0;
  wire n25_carry__0_i_4__1_n_0;
  wire n25_carry__0_n_14;
  wire n25_carry__0_n_15;
  wire n25_carry__0_n_5;
  wire n25_carry__0_n_7;
  wire n25_carry_i_10__1_n_0;
  wire n25_carry_i_11__1_n_0;
  wire n25_carry_i_12__1_n_0;
  wire n25_carry_i_13__0_n_0;
  wire n25_carry_i_14__0_n_0;
  wire n25_carry_i_15__0_n_0;
  wire n25_carry_i_1__1_n_0;
  wire n25_carry_i_2__1_n_0;
  wire n25_carry_i_3__1_n_0;
  wire n25_carry_i_4__1_n_0;
  wire n25_carry_i_5__1_n_0;
  wire n25_carry_i_6__1_n_0;
  wire n25_carry_i_7__0_n_0;
  wire n25_carry_i_8__0_n_0;
  wire n25_carry_i_9__1_n_0;
  wire n25_carry_n_0;
  wire n25_carry_n_1;
  wire n25_carry_n_10;
  wire n25_carry_n_11;
  wire n25_carry_n_12;
  wire n25_carry_n_15;
  wire n25_carry_n_2;
  wire n25_carry_n_3;
  wire n25_carry_n_4;
  wire n25_carry_n_5;
  wire n25_carry_n_6;
  wire n25_carry_n_7;
  wire n25_carry_n_8;
  wire n25_carry_n_9;
  wire [7:0]n26;
  wire [7:0]n27;
  wire [7:0]n29;
  wire [7:0]n2_2;
  wire [7:7]n30;
  wire [7:0]n31;
  wire \n33[10]_i_1__7_n_0 ;
  wire \n33[11]_i_1__7_n_0 ;
  wire \n33[12]_i_1__7_n_0 ;
  wire \n33[12]_i_2__7_n_0 ;
  wire \n33[13]_i_1__7_n_0 ;
  wire \n33[14]_i_1__7_n_0 ;
  wire \n33[14]_i_2__7_n_0 ;
  wire \n33[15]_i_2__7_n_0 ;
  wire \n33[2]_i_1__7_n_0 ;
  wire \n33[3]_i_1__7_n_0 ;
  wire \n33[4]_i_1__7_n_0 ;
  wire \n33[4]_i_2__7_n_0 ;
  wire \n33[5]_i_1__7_n_0 ;
  wire \n33[6]_i_1__7_n_0 ;
  wire \n33[6]_i_2__7_n_0 ;
  wire \n33[7]_i_2__7_n_0 ;
  wire \n33[9]_i_1__7_n_0 ;
  wire [7:0]n341_out;
  wire [7:1]n350_out;
  wire \n37[12]_i_2__7_n_0 ;
  wire \n37[14]_i_2__7_n_0 ;
  wire \n37[15]_i_2__7_n_0 ;
  wire \n37[4]_i_2__7_n_0 ;
  wire \n37[6]_i_2__7_n_0 ;
  wire \n37[7]_i_2__7_n_0 ;
  wire [7:0]\n4_reg[7]_0 ;
  wire \n4_reg_n_0_[0] ;
  wire \n4_reg_n_0_[1] ;
  wire \n4_reg_n_0_[2] ;
  wire \n4_reg_n_0_[3] ;
  wire \n4_reg_n_0_[4] ;
  wire \n4_reg_n_0_[5] ;
  wire \n4_reg_n_0_[6] ;
  wire \n4_reg_n_0_[7] ;
  wire \n7_reg_n_0_[0] ;
  wire \n7_reg_n_0_[1] ;
  wire \n7_reg_n_0_[2] ;
  wire \n7_reg_n_0_[3] ;
  wire \n7_reg_n_0_[4] ;
  wire \n7_reg_n_0_[5] ;
  wire \n7_reg_n_0_[6] ;
  wire \n7_reg_n_0_[7] ;
  wire \n8_reg_n_0_[0] ;
  wire \n8_reg_n_0_[1] ;
  wire \n8_reg_n_0_[2] ;
  wire \n8_reg_n_0_[3] ;
  wire \n8_reg_n_0_[4] ;
  wire \n8_reg_n_0_[5] ;
  wire \n8_reg_n_0_[6] ;
  wire \n8_reg_n_0_[7] ;
  wire \n9_reg_n_0_[0] ;
  wire \n9_reg_n_0_[1] ;
  wire \n9_reg_n_0_[2] ;
  wire \n9_reg_n_0_[3] ;
  wire \n9_reg_n_0_[4] ;
  wire \n9_reg_n_0_[5] ;
  wire \n9_reg_n_0_[6] ;
  wire \n9_reg_n_0_[7] ;
  wire rst_i;
  wire [0:0]NLW_n14__21_carry_O_UNCONNECTED;
  wire [7:1]NLW_n14__21_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n14__21_carry__0_O_UNCONNECTED;
  wire [7:7]NLW_n14__47_carry_CO_UNCONNECTED;
  wire [3:0]NLW_n14__67_carry_O_UNCONNECTED;
  wire [7:3]NLW_n14__67_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n14__67_carry__0_O_UNCONNECTED;
  wire [2:1]NLW_n14_carry_O_UNCONNECTED;
  wire [7:1]NLW_n14_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n14_carry__0_O_UNCONNECTED;
  wire [7:7]\NLW_n21_reg[7]_i_1__3_CO_UNCONNECTED ;
  wire [0:0]NLW_n25__17_carry_O_UNCONNECTED;
  wire [7:1]NLW_n25__17_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n25__17_carry__0_O_UNCONNECTED;
  wire [7:7]NLW_n25__47_carry_CO_UNCONNECTED;
  wire [3:0]NLW_n25__67_carry_O_UNCONNECTED;
  wire [7:3]NLW_n25__67_carry__0_CO_UNCONNECTED;
  wire [7:4]NLW_n25__67_carry__0_O_UNCONNECTED;
  wire [2:1]NLW_n25_carry_O_UNCONNECTED;
  wire [7:1]NLW_n25_carry__0_CO_UNCONNECTED;
  wire [7:2]NLW_n25_carry__0_O_UNCONNECTED;

  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[0] ),
        .Q(n10[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[1] ),
        .Q(n10[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[2] ),
        .Q(n10[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[3] ),
        .Q(n10[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[4] ),
        .Q(n10[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[5] ),
        .Q(n10[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[6] ),
        .Q(n10[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[7] ),
        .Q(n10[7]),
        .R(rst_i));
  FDSE #(
    .INIT(1'b0)) 
    \n11_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(1'b0),
        .Q(B),
        .S(enable_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__21_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__21_carry_n_0,n14__21_carry_n_1,n14__21_carry_n_2,n14__21_carry_n_3,n14__21_carry_n_4,n14__21_carry_n_5,n14__21_carry_n_6,n14__21_carry_n_7}),
        .DI({n14_carry_i_1__1_n_0,n14__21_carry_i_1__1_n_0,n14__21_carry_i_2__1_n_0,n14__21_carry_i_3__1_n_0,n14__21_carry_i_4__1_n_0,n14__21_carry_i_5__1_n_0,n14__21_carry_i_6__0_n_0,1'b0}),
        .O({n14__21_carry_n_8,n14__21_carry_n_9,n14__21_carry_n_10,n14__21_carry_n_11,n14__21_carry_n_12,n14__21_carry_n_13,n14__21_carry_n_14,NLW_n14__21_carry_O_UNCONNECTED[0]}),
        .S({n14__21_carry_i_7__0_n_0,n14__21_carry_i_8__1_n_0,n14__21_carry_i_9__0_n_0,n14__21_carry_i_10__1_n_0,n14__21_carry_i_11__0_n_0,n14__21_carry_i_12__0_n_0,n14__21_carry_i_13__0_n_0,n14__21_carry_i_14__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__21_carry__0
       (.CI(n14__21_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__21_carry__0_CO_UNCONNECTED[7:3],n14__21_carry__0_n_5,NLW_n14__21_carry__0_CO_UNCONNECTED[1],n14__21_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14__21_carry__0_i_1__0_n_0,n14__21_carry__0_i_2__1_n_0}),
        .O({NLW_n14__21_carry__0_O_UNCONNECTED[7:2],n14__21_carry__0_n_14,n14__21_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n14__21_carry__0_i_3__0_n_0,n14__21_carry__0_i_4__1_n_0}));
  LUT3 #(
    .INIT(8'h40)) 
    n14__21_carry__0_i_1__0
       (.I0(n22_n_0),
        .I1(B),
        .I2(n22__0_n_0),
        .O(n14__21_carry__0_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h80C8)) 
    n14__21_carry__0_i_2__1
       (.I0(n22__1_n_0),
        .I1(B),
        .I2(n22__0_n_0),
        .I3(n22_n_0),
        .O(n14__21_carry__0_i_2__1_n_0));
  LUT3 #(
    .INIT(8'h37)) 
    n14__21_carry__0_i_3__0
       (.I0(n22__0_n_0),
        .I1(B),
        .I2(n22_n_0),
        .O(n14__21_carry__0_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h4FDF)) 
    n14__21_carry__0_i_4__1
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(B),
        .I3(n22_n_0),
        .O(n14__21_carry__0_i_4__1_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n14__21_carry_i_10__1
       (.I0(n22__5_n_0),
        .I1(n22__3_n_0),
        .I2(B),
        .I3(n22__4_n_0),
        .I4(n22__2_n_0),
        .O(n14__21_carry_i_10__1_n_0));
  LUT5 #(
    .INIT(32'h66009600)) 
    n14__21_carry_i_11__0
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__5_n_0),
        .I3(B),
        .I4(n22__6_n_0),
        .O(n14__21_carry_i_11__0_n_0));
  LUT4 #(
    .INIT(16'h9060)) 
    n14__21_carry_i_12__0
       (.I0(n22__6_n_0),
        .I1(n22__5_n_0),
        .I2(B),
        .I3(n22__4_n_0),
        .O(n14__21_carry_i_12__0_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n14__21_carry_i_13__0
       (.I0(n22__5_n_0),
        .I1(B),
        .I2(n22__6_n_0),
        .O(n14__21_carry_i_13__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__21_carry_i_14__0
       (.I0(B),
        .I1(n22__6_n_0),
        .O(n14__21_carry_i_14__0_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n14__21_carry_i_1__1
       (.I0(n22__3_n_0),
        .I1(B),
        .I2(n22__2_n_0),
        .I3(n22__1_n_0),
        .O(n14__21_carry_i_1__1_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n14__21_carry_i_2__1
       (.I0(n22__4_n_0),
        .I1(B),
        .I2(n22__3_n_0),
        .I3(n22__2_n_0),
        .O(n14__21_carry_i_2__1_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n14__21_carry_i_3__1
       (.I0(n22__5_n_0),
        .I1(B),
        .I2(n22__4_n_0),
        .I3(n22__3_n_0),
        .O(n14__21_carry_i_3__1_n_0));
  LUT4 #(
    .INIT(16'h8448)) 
    n14__21_carry_i_4__1
       (.I0(n22__4_n_0),
        .I1(B),
        .I2(n22__5_n_0),
        .I3(n22__3_n_0),
        .O(n14__21_carry_i_4__1_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n14__21_carry_i_5__1
       (.I0(n22__5_n_0),
        .I1(B),
        .I2(n22__6_n_0),
        .O(n14__21_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__21_carry_i_6__0
       (.I0(B),
        .I1(n22__5_n_0),
        .O(n14__21_carry_i_6__0_n_0));
  LUT5 #(
    .INIT(32'h95656595)) 
    n14__21_carry_i_7__0
       (.I0(n14_carry_i_1__1_n_0),
        .I1(n22__0_n_0),
        .I2(B),
        .I3(n22__1_n_0),
        .I4(n22_n_0),
        .O(n14__21_carry_i_7__0_n_0));
  (* HLUTNM = "lutpair110" *) 
  LUT5 #(
    .INIT(32'h4C8004C8)) 
    n14__21_carry_i_8__1
       (.I0(n22__2_n_0),
        .I1(B),
        .I2(n22__1_n_0),
        .I3(n22__0_n_0),
        .I4(n22__3_n_0),
        .O(n14__21_carry_i_8__1_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n14__21_carry_i_9__0
       (.I0(n22__4_n_0),
        .I1(n22__2_n_0),
        .I2(B),
        .I3(n22__3_n_0),
        .I4(n22__1_n_0),
        .O(n14__21_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__47_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__47_carry_CO_UNCONNECTED[7],n14__47_carry_n_1,n14__47_carry_n_2,n14__47_carry_n_3,n14__47_carry_n_4,n14__47_carry_n_5,n14__47_carry_n_6,n14__47_carry_n_7}),
        .DI({1'b0,n14__47_carry_i_1__1_n_0,n14__47_carry_i_2__1_n_0,n14__47_carry_i_3__0_n_0,n14__47_carry_i_4__0_n_0,1'b1,1'b0,1'b1}),
        .O({n14__47_carry_n_8,n14__47_carry_n_9,n14__47_carry_n_10,n14__47_carry_n_11,n14__47_carry_n_12,n14__47_carry_n_13,n14__47_carry_n_14,n14__47_carry_n_15}),
        .S({n14__47_carry_i_5__0_n_0,n14__47_carry_i_6__1_n_0,n14__47_carry_i_7__0_n_0,n14__47_carry_i_8__0_n_0,n14__47_carry_i_9__0_n_0,n14__47_carry_i_10__0_n_0,n14__47_carry_i_11__0_n_0,n14__47_carry_i_12__0_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n14__47_carry_i_10__0
       (.I0(B),
        .I1(n22__3_n_0),
        .O(n14__47_carry_i_10__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__47_carry_i_11__0
       (.I0(B),
        .I1(n22__4_n_0),
        .O(n14__47_carry_i_11__0_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n14__47_carry_i_12__0
       (.I0(n22__5_n_0),
        .I1(B),
        .O(n14__47_carry_i_12__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__47_carry_i_1__1
       (.I0(B),
        .I1(n22__0_n_0),
        .O(n14__47_carry_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__47_carry_i_2__1
       (.I0(B),
        .I1(n22__1_n_0),
        .O(n14__47_carry_i_2__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__47_carry_i_3__0
       (.I0(B),
        .I1(n22__2_n_0),
        .O(n14__47_carry_i_3__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__47_carry_i_4__0
       (.I0(B),
        .I1(n22__3_n_0),
        .O(n14__47_carry_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n14__47_carry_i_5__0
       (.I0(n22_n_0),
        .I1(B),
        .O(n14__47_carry_i_5__0_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n14__47_carry_i_6__1
       (.I0(n22__0_n_0),
        .I1(B),
        .I2(n22_n_0),
        .O(n14__47_carry_i_6__1_n_0));
  LUT3 #(
    .INIT(8'hB7)) 
    n14__47_carry_i_7__0
       (.I0(n22__1_n_0),
        .I1(B),
        .I2(n22__0_n_0),
        .O(n14__47_carry_i_7__0_n_0));
  LUT3 #(
    .INIT(8'hB7)) 
    n14__47_carry_i_8__0
       (.I0(n22__2_n_0),
        .I1(B),
        .I2(n22__1_n_0),
        .O(n14__47_carry_i_8__0_n_0));
  LUT3 #(
    .INIT(8'hB7)) 
    n14__47_carry_i_9__0
       (.I0(n22__3_n_0),
        .I1(B),
        .I2(n22__2_n_0),
        .O(n14__47_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__67_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14__67_carry_n_0,n14__67_carry_n_1,n14__67_carry_n_2,n14__67_carry_n_3,n14__67_carry_n_4,n14__67_carry_n_5,n14__67_carry_n_6,n14__67_carry_n_7}),
        .DI({n14__67_carry_i_1__1_n_0,n14__67_carry_i_2__1_n_0,n14__67_carry_i_3__1_n_0,n14__67_carry_i_4__1_n_0,n14__67_carry_i_5__1_n_0,n14__67_carry_i_6__1_n_0,n14__67_carry_i_7__1_n_0,1'b0}),
        .O({n15[3:0],NLW_n14__67_carry_O_UNCONNECTED[3:0]}),
        .S({n14__67_carry_i_8__1_n_0,n14__67_carry_i_9__1_n_0,n14__67_carry_i_10__1_n_0,n14__67_carry_i_11__1_n_0,n14__67_carry_i_12__1_n_0,n14__67_carry_i_13__1_n_0,n14__67_carry_i_14__1_n_0,n14__67_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14__67_carry__0
       (.CI(n14__67_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14__67_carry__0_CO_UNCONNECTED[7:3],n14__67_carry__0_n_5,n14__67_carry__0_n_6,n14__67_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n14__67_carry__0_i_1__1_n_0,n14__67_carry__0_i_2__1_n_0,n14__67_carry__0_i_3__1_n_0}),
        .O({NLW_n14__67_carry__0_O_UNCONNECTED[7:4],n15[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n14__67_carry__0_i_4__1_n_0,n14__67_carry__0_i_5__1_n_0,n14__67_carry__0_i_6__1_n_0,n14__67_carry__0_i_7__1_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry__0_i_1__1
       (.I0(n14__21_carry__0_n_14),
        .I1(n14__47_carry_n_10),
        .O(n14__67_carry__0_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry__0_i_2__1
       (.I0(n14__21_carry__0_n_15),
        .I1(n14__47_carry_n_11),
        .O(n14__67_carry__0_i_2__1_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n14__67_carry__0_i_3__1
       (.I0(n14__47_carry_n_12),
        .I1(n14__21_carry_n_8),
        .I2(n14_carry__0_n_5),
        .O(n14__67_carry__0_i_3__1_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n14__67_carry__0_i_4__1
       (.I0(n14__21_carry__0_n_5),
        .I1(n14__47_carry_n_9),
        .I2(n14__47_carry_n_8),
        .O(n14__67_carry__0_i_4__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__67_carry__0_i_5__1
       (.I0(n14__21_carry__0_n_14),
        .I1(n14__47_carry_n_10),
        .I2(n14__47_carry_n_9),
        .I3(n14__21_carry__0_n_5),
        .O(n14__67_carry__0_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__67_carry__0_i_6__1
       (.I0(n14__21_carry__0_n_15),
        .I1(n14__47_carry_n_11),
        .I2(n14__47_carry_n_10),
        .I3(n14__21_carry__0_n_14),
        .O(n14__67_carry__0_i_6__1_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n14__67_carry__0_i_7__1
       (.I0(n14_carry__0_n_5),
        .I1(n14__21_carry_n_8),
        .I2(n14__47_carry_n_12),
        .I3(n14__47_carry_n_11),
        .I4(n14__21_carry__0_n_15),
        .O(n14__67_carry__0_i_7__1_n_0));
  (* HLUTNM = "lutpair78" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__67_carry_i_10__1
       (.I0(n14__47_carry_n_14),
        .I1(n14__21_carry_n_10),
        .I2(n14_carry__0_n_15),
        .I3(n14__67_carry_i_3__1_n_0),
        .O(n14__67_carry_i_10__1_n_0));
  (* HLUTNM = "lutpair77" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__67_carry_i_11__1
       (.I0(n14__47_carry_n_15),
        .I1(n14__21_carry_n_11),
        .I2(n14_carry_n_8),
        .I3(n14__67_carry_i_4__1_n_0),
        .O(n14__67_carry_i_11__1_n_0));
  (* HLUTNM = "lutpair76" *) 
  LUT5 #(
    .INIT(32'h78878778)) 
    n14__67_carry_i_12__1
       (.I0(B),
        .I1(n22__6_n_0),
        .I2(n14__21_carry_n_12),
        .I3(n14_carry_n_9),
        .I4(n14__67_carry_i_5__1_n_0),
        .O(n14__67_carry_i_12__1_n_0));
  (* HLUTNM = "lutpair111" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n14__67_carry_i_13__1
       (.I0(n14__21_carry_n_13),
        .I1(n14_carry_n_10),
        .I2(n14_carry_n_11),
        .I3(n14__21_carry_n_14),
        .O(n14__67_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n14__67_carry_i_14__1
       (.I0(n14_carry_n_12),
        .I1(n14_carry_n_15),
        .I2(n14__21_carry_n_14),
        .I3(n14_carry_n_11),
        .O(n14__67_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n14__67_carry_i_15__1
       (.I0(n14_carry_n_12),
        .I1(n14_carry_n_15),
        .O(n14__67_carry_i_15__1_n_0));
  (* HLUTNM = "lutpair79" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__67_carry_i_1__1
       (.I0(n14__47_carry_n_13),
        .I1(n14__21_carry_n_9),
        .I2(n14_carry__0_n_14),
        .O(n14__67_carry_i_1__1_n_0));
  (* HLUTNM = "lutpair78" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__67_carry_i_2__1
       (.I0(n14__47_carry_n_14),
        .I1(n14__21_carry_n_10),
        .I2(n14_carry__0_n_15),
        .O(n14__67_carry_i_2__1_n_0));
  (* HLUTNM = "lutpair77" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n14__67_carry_i_3__1
       (.I0(n14__47_carry_n_15),
        .I1(n14__21_carry_n_11),
        .I2(n14_carry_n_8),
        .O(n14__67_carry_i_3__1_n_0));
  (* HLUTNM = "lutpair76" *) 
  LUT4 #(
    .INIT(16'hF880)) 
    n14__67_carry_i_4__1
       (.I0(B),
        .I1(n22__6_n_0),
        .I2(n14__21_carry_n_12),
        .I3(n14_carry_n_9),
        .O(n14__67_carry_i_4__1_n_0));
  (* HLUTNM = "lutpair111" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry_i_5__1
       (.I0(n14__21_carry_n_13),
        .I1(n14_carry_n_10),
        .O(n14__67_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry_i_6__1
       (.I0(n14_carry_n_11),
        .I1(n14__21_carry_n_14),
        .O(n14__67_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14__67_carry_i_7__1
       (.I0(n14_carry_n_12),
        .I1(n14_carry_n_15),
        .O(n14__67_carry_i_7__1_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n14__67_carry_i_8__1
       (.I0(n14__67_carry_i_1__1_n_0),
        .I1(n14__21_carry_n_8),
        .I2(n14__47_carry_n_12),
        .I3(n14_carry__0_n_5),
        .O(n14__67_carry_i_8__1_n_0));
  (* HLUTNM = "lutpair79" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n14__67_carry_i_9__1
       (.I0(n14__47_carry_n_13),
        .I1(n14__21_carry_n_9),
        .I2(n14_carry__0_n_14),
        .I3(n14__67_carry_i_2__1_n_0),
        .O(n14__67_carry_i_9__1_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n14_carry_n_0,n14_carry_n_1,n14_carry_n_2,n14_carry_n_3,n14_carry_n_4,n14_carry_n_5,n14_carry_n_6,n14_carry_n_7}),
        .DI({n14_carry_i_1__1_n_0,n14_carry_i_2__1_n_0,n14_carry_i_3__1_n_0,n14_carry_i_4__1_n_0,n14_carry_i_5__1_n_0,n14_carry_i_6__1_n_0,n14_carry_i_7__0_n_0,1'b0}),
        .O({n14_carry_n_8,n14_carry_n_9,n14_carry_n_10,n14_carry_n_11,n14_carry_n_12,NLW_n14_carry_O_UNCONNECTED[2:1],n14_carry_n_15}),
        .S({n14_carry_i_8__0_n_0,n14_carry_i_9__1_n_0,n14_carry_i_10__1_n_0,n14_carry_i_11__1_n_0,n14_carry_i_12__1_n_0,n14_carry_i_13__0_n_0,n14_carry_i_14__0_n_0,n14_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n14_carry__0
       (.CI(n14_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n14_carry__0_CO_UNCONNECTED[7:3],n14_carry__0_n_5,NLW_n14_carry__0_CO_UNCONNECTED[1],n14_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n14_carry__0_i_1__1_n_0,n14_carry__0_i_2__1_n_0}),
        .O({NLW_n14_carry__0_O_UNCONNECTED[7:2],n14_carry__0_n_14,n14_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n14_carry__0_i_3__0_n_0,n14_carry__0_i_4__1_n_0}));
  LUT3 #(
    .INIT(8'h40)) 
    n14_carry__0_i_1__1
       (.I0(n22_n_0),
        .I1(B),
        .I2(n22__0_n_0),
        .O(n14_carry__0_i_1__1_n_0));
  LUT4 #(
    .INIT(16'h80C8)) 
    n14_carry__0_i_2__1
       (.I0(n22__1_n_0),
        .I1(B),
        .I2(n22__0_n_0),
        .I3(n22_n_0),
        .O(n14_carry__0_i_2__1_n_0));
  LUT3 #(
    .INIT(8'h37)) 
    n14_carry__0_i_3__0
       (.I0(n22__0_n_0),
        .I1(B),
        .I2(n22_n_0),
        .O(n14_carry__0_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h4FDF)) 
    n14_carry__0_i_4__1
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(B),
        .I3(n22_n_0),
        .O(n14_carry__0_i_4__1_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n14_carry_i_10__1
       (.I0(n22__4_n_0),
        .I1(n22__2_n_0),
        .I2(B),
        .I3(n22__3_n_0),
        .I4(n22__1_n_0),
        .O(n14_carry_i_10__1_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n14_carry_i_11__1
       (.I0(n22__5_n_0),
        .I1(n22__3_n_0),
        .I2(B),
        .I3(n22__4_n_0),
        .I4(n22__2_n_0),
        .O(n14_carry_i_11__1_n_0));
  LUT5 #(
    .INIT(32'h66009600)) 
    n14_carry_i_12__1
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__5_n_0),
        .I3(B),
        .I4(n22__6_n_0),
        .O(n14_carry_i_12__1_n_0));
  LUT4 #(
    .INIT(16'h9060)) 
    n14_carry_i_13__0
       (.I0(n22__6_n_0),
        .I1(n22__5_n_0),
        .I2(B),
        .I3(n22__4_n_0),
        .O(n14_carry_i_13__0_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n14_carry_i_14__0
       (.I0(n22__5_n_0),
        .I1(B),
        .I2(n22__6_n_0),
        .O(n14_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14_carry_i_15__0
       (.I0(B),
        .I1(n22__6_n_0),
        .O(n14_carry_i_15__0_n_0));
  (* HLUTNM = "lutpair110" *) 
  LUT4 #(
    .INIT(16'hC880)) 
    n14_carry_i_1__1
       (.I0(n22__2_n_0),
        .I1(B),
        .I2(n22__1_n_0),
        .I3(n22__0_n_0),
        .O(n14_carry_i_1__1_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n14_carry_i_2__1
       (.I0(n22__3_n_0),
        .I1(B),
        .I2(n22__2_n_0),
        .I3(n22__1_n_0),
        .O(n14_carry_i_2__1_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n14_carry_i_3__1
       (.I0(n22__4_n_0),
        .I1(B),
        .I2(n22__3_n_0),
        .I3(n22__2_n_0),
        .O(n14_carry_i_3__1_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n14_carry_i_4__1
       (.I0(n22__5_n_0),
        .I1(B),
        .I2(n22__4_n_0),
        .I3(n22__3_n_0),
        .O(n14_carry_i_4__1_n_0));
  LUT4 #(
    .INIT(16'h8448)) 
    n14_carry_i_5__1
       (.I0(n22__4_n_0),
        .I1(B),
        .I2(n22__5_n_0),
        .I3(n22__3_n_0),
        .O(n14_carry_i_5__1_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n14_carry_i_6__1
       (.I0(n22__5_n_0),
        .I1(B),
        .I2(n22__6_n_0),
        .O(n14_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n14_carry_i_7__0
       (.I0(B),
        .I1(n22__5_n_0),
        .O(n14_carry_i_7__0_n_0));
  LUT5 #(
    .INIT(32'h95656595)) 
    n14_carry_i_8__0
       (.I0(n14_carry_i_1__1_n_0),
        .I1(n22__0_n_0),
        .I2(B),
        .I3(n22__1_n_0),
        .I4(n22_n_0),
        .O(n14_carry_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n14_carry_i_9__1
       (.I0(n22__3_n_0),
        .I1(n22__1_n_0),
        .I2(B),
        .I3(n22__2_n_0),
        .I4(n22__0_n_0),
        .O(n14_carry_i_9__1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[0]),
        .Q(\n16_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[1]),
        .Q(\n16_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[2]),
        .Q(\n16_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[3]),
        .Q(\n16_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[4]),
        .Q(\n16_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[5]),
        .Q(\n16_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[6]),
        .Q(\n16_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[7]),
        .Q(\n16_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [0]),
        .Q(\n1_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [10]),
        .Q(n2_2[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [11]),
        .Q(n2_2[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [12]),
        .Q(n2_2[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [13]),
        .Q(n2_2[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [14]),
        .Q(n2_2[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [15]),
        .Q(n2_2[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [1]),
        .Q(\n1_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [2]),
        .Q(\n1_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [3]),
        .Q(\n1_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [4]),
        .Q(\n1_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [5]),
        .Q(\n1_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [6]),
        .Q(\n1_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [7]),
        .Q(\n1_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [8]),
        .Q(n2_2[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg[15]_0 [9]),
        .Q(n2_2[1]),
        .R(rst_i));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_2 
       (.I0(\n16_reg_n_0_[7] ),
        .O(\n21[7]_i_2_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_3 
       (.I0(\n16_reg_n_0_[6] ),
        .O(\n21[7]_i_3_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_4 
       (.I0(\n16_reg_n_0_[5] ),
        .O(\n21[7]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_5 
       (.I0(\n16_reg_n_0_[4] ),
        .O(\n21[7]_i_5_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_6 
       (.I0(\n16_reg_n_0_[3] ),
        .O(\n21[7]_i_6_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_7 
       (.I0(\n16_reg_n_0_[2] ),
        .O(\n21[7]_i_7_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_8 
       (.I0(\n16_reg_n_0_[1] ),
        .O(\n21[7]_i_8_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_9 
       (.I0(\n16_reg_n_0_[0] ),
        .O(\n21[7]_i_9_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[0]),
        .Q(n21[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[1]),
        .Q(n21[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[2]),
        .Q(n21[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[3]),
        .Q(n21[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[4]),
        .Q(n21[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[5]),
        .Q(n21[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[6]),
        .Q(n21[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[7]),
        .Q(n21[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n21_reg[7]_i_1__3 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\NLW_n21_reg[7]_i_1__3_CO_UNCONNECTED [7],\n21_reg[7]_i_1__3_n_1 ,\n21_reg[7]_i_1__3_n_2 ,\n21_reg[7]_i_1__3_n_3 ,\n21_reg[7]_i_1__3_n_4 ,\n21_reg[7]_i_1__3_n_5 ,\n21_reg[7]_i_1__3_n_6 ,\n21_reg[7]_i_1__3_n_7 }),
        .DI({1'b0,\n16_reg_n_0_[6] ,\n16_reg_n_0_[5] ,\n16_reg_n_0_[4] ,\n16_reg_n_0_[3] ,\n16_reg_n_0_[2] ,\n16_reg_n_0_[1] ,\n16_reg_n_0_[0] }),
        .O(n202_out),
        .S({\n21[7]_i_2_n_0 ,\n21[7]_i_3_n_0 ,\n21[7]_i_4_n_0 ,\n21[7]_i_5_n_0 ,\n21[7]_i_6_n_0 ,\n21[7]_i_7_n_0 ,\n21[7]_i_8_n_0 ,\n21[7]_i_9_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    n22
       (.C(clk_i),
        .CE(enable_i),
        .D(n22_0[7]),
        .Q(n22_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__0
       (.C(clk_i),
        .CE(enable_i),
        .D(n22_0[6]),
        .Q(n22__0_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__1
       (.C(clk_i),
        .CE(enable_i),
        .D(n22_0[5]),
        .Q(n22__1_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__2
       (.C(clk_i),
        .CE(enable_i),
        .D(n22_0[4]),
        .Q(n22__2_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__3
       (.C(clk_i),
        .CE(enable_i),
        .D(n22_0[3]),
        .Q(n22__3_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__4
       (.C(clk_i),
        .CE(enable_i),
        .D(n22_0[2]),
        .Q(n22__4_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__5
       (.C(clk_i),
        .CE(enable_i),
        .D(n22_0[1]),
        .Q(n22__5_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__6
       (.C(clk_i),
        .CE(enable_i),
        .D(n22_0[0]),
        .Q(n22__6_n_0),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__17_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__17_carry_n_0,n25__17_carry_n_1,n25__17_carry_n_2,n25__17_carry_n_3,n25__17_carry_n_4,n25__17_carry_n_5,n25__17_carry_n_6,n25__17_carry_n_7}),
        .DI({n25_carry_i_1__1_n_0,n25__17_carry_i_1__1_n_0,n25__17_carry_i_2__1_n_0,n25__17_carry_i_3__1_n_0,n25__17_carry_i_4__1_n_0,n25__17_carry_i_5__1_n_0,n25__17_carry_i_6__0_n_0,1'b0}),
        .O({n25__17_carry_n_8,n25__17_carry_n_9,n25__17_carry_n_10,n25__17_carry_n_11,n25__17_carry_n_12,n25__17_carry_n_13,n25__17_carry_n_14,NLW_n25__17_carry_O_UNCONNECTED[0]}),
        .S({n25__17_carry_i_7__0_n_0,n25__17_carry_i_8__1_n_0,n25__17_carry_i_9__0_n_0,n25__17_carry_i_10__1_n_0,n25__17_carry_i_11__0_n_0,n25__17_carry_i_12__0_n_0,n25__17_carry_i_13__0_n_0,n25__17_carry_i_14__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__17_carry__0
       (.CI(n25__17_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__17_carry__0_CO_UNCONNECTED[7:3],n25__17_carry__0_n_5,NLW_n25__17_carry__0_CO_UNCONNECTED[1],n25__17_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25__17_carry__0_i_1__0_n_0,n25__17_carry__0_i_2__1_n_0}),
        .O({NLW_n25__17_carry__0_O_UNCONNECTED[7:2],n25__17_carry__0_n_14,n25__17_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n25__17_carry__0_i_3__0_n_0,n25__17_carry__0_i_4__1_n_0}));
  LUT3 #(
    .INIT(8'h40)) 
    n25__17_carry__0_i_1__0
       (.I0(\n4_reg_n_0_[7] ),
        .I1(B),
        .I2(\n4_reg_n_0_[6] ),
        .O(n25__17_carry__0_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h80C8)) 
    n25__17_carry__0_i_2__1
       (.I0(\n4_reg_n_0_[5] ),
        .I1(B),
        .I2(\n4_reg_n_0_[6] ),
        .I3(\n4_reg_n_0_[7] ),
        .O(n25__17_carry__0_i_2__1_n_0));
  LUT3 #(
    .INIT(8'h37)) 
    n25__17_carry__0_i_3__0
       (.I0(\n4_reg_n_0_[6] ),
        .I1(B),
        .I2(\n4_reg_n_0_[7] ),
        .O(n25__17_carry__0_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h4FDF)) 
    n25__17_carry__0_i_4__1
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(B),
        .I3(\n4_reg_n_0_[7] ),
        .O(n25__17_carry__0_i_4__1_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n25__17_carry_i_10__1
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(B),
        .I3(\n4_reg_n_0_[2] ),
        .I4(\n4_reg_n_0_[4] ),
        .O(n25__17_carry_i_10__1_n_0));
  LUT5 #(
    .INIT(32'h66009600)) 
    n25__17_carry_i_11__0
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[1] ),
        .I3(B),
        .I4(\n4_reg_n_0_[0] ),
        .O(n25__17_carry_i_11__0_n_0));
  LUT4 #(
    .INIT(16'h9060)) 
    n25__17_carry_i_12__0
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(B),
        .I3(\n4_reg_n_0_[2] ),
        .O(n25__17_carry_i_12__0_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n25__17_carry_i_13__0
       (.I0(\n4_reg_n_0_[1] ),
        .I1(B),
        .I2(\n4_reg_n_0_[0] ),
        .O(n25__17_carry_i_13__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__17_carry_i_14__0
       (.I0(B),
        .I1(\n4_reg_n_0_[0] ),
        .O(n25__17_carry_i_14__0_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n25__17_carry_i_1__1
       (.I0(\n4_reg_n_0_[3] ),
        .I1(B),
        .I2(\n4_reg_n_0_[4] ),
        .I3(\n4_reg_n_0_[5] ),
        .O(n25__17_carry_i_1__1_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n25__17_carry_i_2__1
       (.I0(\n4_reg_n_0_[2] ),
        .I1(B),
        .I2(\n4_reg_n_0_[3] ),
        .I3(\n4_reg_n_0_[4] ),
        .O(n25__17_carry_i_2__1_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n25__17_carry_i_3__1
       (.I0(\n4_reg_n_0_[1] ),
        .I1(B),
        .I2(\n4_reg_n_0_[2] ),
        .I3(\n4_reg_n_0_[3] ),
        .O(n25__17_carry_i_3__1_n_0));
  LUT4 #(
    .INIT(16'h8448)) 
    n25__17_carry_i_4__1
       (.I0(\n4_reg_n_0_[2] ),
        .I1(B),
        .I2(\n4_reg_n_0_[1] ),
        .I3(\n4_reg_n_0_[3] ),
        .O(n25__17_carry_i_4__1_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n25__17_carry_i_5__1
       (.I0(\n4_reg_n_0_[1] ),
        .I1(B),
        .I2(\n4_reg_n_0_[0] ),
        .O(n25__17_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__17_carry_i_6__0
       (.I0(B),
        .I1(\n4_reg_n_0_[1] ),
        .O(n25__17_carry_i_6__0_n_0));
  LUT5 #(
    .INIT(32'h95656595)) 
    n25__17_carry_i_7__0
       (.I0(n25_carry_i_1__1_n_0),
        .I1(\n4_reg_n_0_[6] ),
        .I2(B),
        .I3(\n4_reg_n_0_[5] ),
        .I4(\n4_reg_n_0_[7] ),
        .O(n25__17_carry_i_7__0_n_0));
  (* HLUTNM = "lutpair108" *) 
  LUT5 #(
    .INIT(32'h4C8004C8)) 
    n25__17_carry_i_8__1
       (.I0(\n4_reg_n_0_[4] ),
        .I1(B),
        .I2(\n4_reg_n_0_[5] ),
        .I3(\n4_reg_n_0_[6] ),
        .I4(\n4_reg_n_0_[3] ),
        .O(n25__17_carry_i_8__1_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n25__17_carry_i_9__0
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(B),
        .I3(\n4_reg_n_0_[3] ),
        .I4(\n4_reg_n_0_[5] ),
        .O(n25__17_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__47_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__47_carry_CO_UNCONNECTED[7],n25__47_carry_n_1,n25__47_carry_n_2,n25__47_carry_n_3,n25__47_carry_n_4,n25__47_carry_n_5,n25__47_carry_n_6,n25__47_carry_n_7}),
        .DI({1'b0,n25__47_carry_i_1__1_n_0,n25__47_carry_i_2__1_n_0,n25__47_carry_i_3__0_n_0,n25__47_carry_i_4__0_n_0,1'b1,1'b0,1'b1}),
        .O({n25__47_carry_n_8,n25__47_carry_n_9,n25__47_carry_n_10,n25__47_carry_n_11,n25__47_carry_n_12,n25__47_carry_n_13,n25__47_carry_n_14,n25__47_carry_n_15}),
        .S({n25__47_carry_i_5__0_n_0,n25__47_carry_i_6__1_n_0,n25__47_carry_i_7__0_n_0,n25__47_carry_i_8__0_n_0,n25__47_carry_i_9__0_n_0,n25__47_carry_i_10__0_n_0,n25__47_carry_i_11__0_n_0,n25__47_carry_i_12__0_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n25__47_carry_i_10__0
       (.I0(B),
        .I1(\n4_reg_n_0_[3] ),
        .O(n25__47_carry_i_10__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__47_carry_i_11__0
       (.I0(B),
        .I1(\n4_reg_n_0_[2] ),
        .O(n25__47_carry_i_11__0_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n25__47_carry_i_12__0
       (.I0(\n4_reg_n_0_[1] ),
        .I1(B),
        .O(n25__47_carry_i_12__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__47_carry_i_1__1
       (.I0(B),
        .I1(\n4_reg_n_0_[6] ),
        .O(n25__47_carry_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__47_carry_i_2__1
       (.I0(B),
        .I1(\n4_reg_n_0_[5] ),
        .O(n25__47_carry_i_2__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__47_carry_i_3__0
       (.I0(B),
        .I1(\n4_reg_n_0_[4] ),
        .O(n25__47_carry_i_3__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__47_carry_i_4__0
       (.I0(B),
        .I1(\n4_reg_n_0_[3] ),
        .O(n25__47_carry_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    n25__47_carry_i_5__0
       (.I0(\n4_reg_n_0_[7] ),
        .I1(B),
        .O(n25__47_carry_i_5__0_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n25__47_carry_i_6__1
       (.I0(\n4_reg_n_0_[6] ),
        .I1(B),
        .I2(\n4_reg_n_0_[7] ),
        .O(n25__47_carry_i_6__1_n_0));
  LUT3 #(
    .INIT(8'hB7)) 
    n25__47_carry_i_7__0
       (.I0(\n4_reg_n_0_[5] ),
        .I1(B),
        .I2(\n4_reg_n_0_[6] ),
        .O(n25__47_carry_i_7__0_n_0));
  LUT3 #(
    .INIT(8'hB7)) 
    n25__47_carry_i_8__0
       (.I0(\n4_reg_n_0_[4] ),
        .I1(B),
        .I2(\n4_reg_n_0_[5] ),
        .O(n25__47_carry_i_8__0_n_0));
  LUT3 #(
    .INIT(8'hB7)) 
    n25__47_carry_i_9__0
       (.I0(\n4_reg_n_0_[3] ),
        .I1(B),
        .I2(\n4_reg_n_0_[4] ),
        .O(n25__47_carry_i_9__0_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__67_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25__67_carry_n_0,n25__67_carry_n_1,n25__67_carry_n_2,n25__67_carry_n_3,n25__67_carry_n_4,n25__67_carry_n_5,n25__67_carry_n_6,n25__67_carry_n_7}),
        .DI({n25__67_carry_i_1__1_n_0,n25__67_carry_i_2__1_n_0,n25__67_carry_i_3__1_n_0,n25__67_carry_i_4__1_n_0,n25__67_carry_i_5__1_n_0,n25__67_carry_i_6__1_n_0,n25__67_carry_i_7__1_n_0,1'b0}),
        .O({n26[3:0],NLW_n25__67_carry_O_UNCONNECTED[3:0]}),
        .S({n25__67_carry_i_8__1_n_0,n25__67_carry_i_9__1_n_0,n25__67_carry_i_10__1_n_0,n25__67_carry_i_11__1_n_0,n25__67_carry_i_12__1_n_0,n25__67_carry_i_13__1_n_0,n25__67_carry_i_14__1_n_0,n25__67_carry_i_15__1_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25__67_carry__0
       (.CI(n25__67_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25__67_carry__0_CO_UNCONNECTED[7:3],n25__67_carry__0_n_5,n25__67_carry__0_n_6,n25__67_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,n25__67_carry__0_i_1__1_n_0,n25__67_carry__0_i_2__1_n_0,n25__67_carry__0_i_3__1_n_0}),
        .O({NLW_n25__67_carry__0_O_UNCONNECTED[7:4],n26[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,n25__67_carry__0_i_4__1_n_0,n25__67_carry__0_i_5__1_n_0,n25__67_carry__0_i_6__1_n_0,n25__67_carry__0_i_7__1_n_0}));
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry__0_i_1__1
       (.I0(n25__17_carry__0_n_14),
        .I1(n25__47_carry_n_10),
        .O(n25__67_carry__0_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry__0_i_2__1
       (.I0(n25__17_carry__0_n_15),
        .I1(n25__47_carry_n_11),
        .O(n25__67_carry__0_i_2__1_n_0));
  LUT3 #(
    .INIT(8'hE8)) 
    n25__67_carry__0_i_3__1
       (.I0(n25__47_carry_n_12),
        .I1(n25__17_carry_n_8),
        .I2(n25_carry__0_n_5),
        .O(n25__67_carry__0_i_3__1_n_0));
  LUT3 #(
    .INIT(8'h78)) 
    n25__67_carry__0_i_4__1
       (.I0(n25__17_carry__0_n_5),
        .I1(n25__47_carry_n_9),
        .I2(n25__47_carry_n_8),
        .O(n25__67_carry__0_i_4__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__67_carry__0_i_5__1
       (.I0(n25__17_carry__0_n_14),
        .I1(n25__47_carry_n_10),
        .I2(n25__47_carry_n_9),
        .I3(n25__17_carry__0_n_5),
        .O(n25__67_carry__0_i_5__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__67_carry__0_i_6__1
       (.I0(n25__17_carry__0_n_15),
        .I1(n25__47_carry_n_11),
        .I2(n25__47_carry_n_10),
        .I3(n25__17_carry__0_n_14),
        .O(n25__67_carry__0_i_6__1_n_0));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    n25__67_carry__0_i_7__1
       (.I0(n25_carry__0_n_5),
        .I1(n25__17_carry_n_8),
        .I2(n25__47_carry_n_12),
        .I3(n25__47_carry_n_11),
        .I4(n25__17_carry__0_n_15),
        .O(n25__67_carry__0_i_7__1_n_0));
  (* HLUTNM = "lutpair74" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__67_carry_i_10__1
       (.I0(n25__47_carry_n_14),
        .I1(n25__17_carry_n_10),
        .I2(n25_carry__0_n_15),
        .I3(n25__67_carry_i_3__1_n_0),
        .O(n25__67_carry_i_10__1_n_0));
  (* HLUTNM = "lutpair73" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__67_carry_i_11__1
       (.I0(n25__47_carry_n_15),
        .I1(n25__17_carry_n_11),
        .I2(n25_carry_n_8),
        .I3(n25__67_carry_i_4__1_n_0),
        .O(n25__67_carry_i_11__1_n_0));
  (* HLUTNM = "lutpair72" *) 
  LUT5 #(
    .INIT(32'h78878778)) 
    n25__67_carry_i_12__1
       (.I0(B),
        .I1(\n4_reg_n_0_[0] ),
        .I2(n25__17_carry_n_12),
        .I3(n25_carry_n_9),
        .I4(n25__67_carry_i_5__1_n_0),
        .O(n25__67_carry_i_12__1_n_0));
  (* HLUTNM = "lutpair109" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    n25__67_carry_i_13__1
       (.I0(n25__17_carry_n_13),
        .I1(n25_carry_n_10),
        .I2(n25_carry_n_11),
        .I3(n25__17_carry_n_14),
        .O(n25__67_carry_i_13__1_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    n25__67_carry_i_14__1
       (.I0(n25_carry_n_12),
        .I1(n25_carry_n_15),
        .I2(n25__17_carry_n_14),
        .I3(n25_carry_n_11),
        .O(n25__67_carry_i_14__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    n25__67_carry_i_15__1
       (.I0(n25_carry_n_12),
        .I1(n25_carry_n_15),
        .O(n25__67_carry_i_15__1_n_0));
  (* HLUTNM = "lutpair75" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__67_carry_i_1__1
       (.I0(n25__47_carry_n_13),
        .I1(n25__17_carry_n_9),
        .I2(n25_carry__0_n_14),
        .O(n25__67_carry_i_1__1_n_0));
  (* HLUTNM = "lutpair74" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__67_carry_i_2__1
       (.I0(n25__47_carry_n_14),
        .I1(n25__17_carry_n_10),
        .I2(n25_carry__0_n_15),
        .O(n25__67_carry_i_2__1_n_0));
  (* HLUTNM = "lutpair73" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    n25__67_carry_i_3__1
       (.I0(n25__47_carry_n_15),
        .I1(n25__17_carry_n_11),
        .I2(n25_carry_n_8),
        .O(n25__67_carry_i_3__1_n_0));
  (* HLUTNM = "lutpair72" *) 
  LUT4 #(
    .INIT(16'hF880)) 
    n25__67_carry_i_4__1
       (.I0(B),
        .I1(\n4_reg_n_0_[0] ),
        .I2(n25__17_carry_n_12),
        .I3(n25_carry_n_9),
        .O(n25__67_carry_i_4__1_n_0));
  (* HLUTNM = "lutpair109" *) 
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry_i_5__1
       (.I0(n25__17_carry_n_13),
        .I1(n25_carry_n_10),
        .O(n25__67_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry_i_6__1
       (.I0(n25_carry_n_11),
        .I1(n25__17_carry_n_14),
        .O(n25__67_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25__67_carry_i_7__1
       (.I0(n25_carry_n_12),
        .I1(n25_carry_n_15),
        .O(n25__67_carry_i_7__1_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    n25__67_carry_i_8__1
       (.I0(n25__67_carry_i_1__1_n_0),
        .I1(n25__17_carry_n_8),
        .I2(n25__47_carry_n_12),
        .I3(n25_carry__0_n_5),
        .O(n25__67_carry_i_8__1_n_0));
  (* HLUTNM = "lutpair75" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    n25__67_carry_i_9__1
       (.I0(n25__47_carry_n_13),
        .I1(n25__17_carry_n_9),
        .I2(n25_carry__0_n_14),
        .I3(n25__67_carry_i_2__1_n_0),
        .O(n25__67_carry_i_9__1_n_0));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25_carry
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({n25_carry_n_0,n25_carry_n_1,n25_carry_n_2,n25_carry_n_3,n25_carry_n_4,n25_carry_n_5,n25_carry_n_6,n25_carry_n_7}),
        .DI({n25_carry_i_1__1_n_0,n25_carry_i_2__1_n_0,n25_carry_i_3__1_n_0,n25_carry_i_4__1_n_0,n25_carry_i_5__1_n_0,n25_carry_i_6__1_n_0,n25_carry_i_7__0_n_0,1'b0}),
        .O({n25_carry_n_8,n25_carry_n_9,n25_carry_n_10,n25_carry_n_11,n25_carry_n_12,NLW_n25_carry_O_UNCONNECTED[2:1],n25_carry_n_15}),
        .S({n25_carry_i_8__0_n_0,n25_carry_i_9__1_n_0,n25_carry_i_10__1_n_0,n25_carry_i_11__1_n_0,n25_carry_i_12__1_n_0,n25_carry_i_13__0_n_0,n25_carry_i_14__0_n_0,n25_carry_i_15__0_n_0}));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    n25_carry__0
       (.CI(n25_carry_n_0),
        .CI_TOP(1'b0),
        .CO({NLW_n25_carry__0_CO_UNCONNECTED[7:3],n25_carry__0_n_5,NLW_n25_carry__0_CO_UNCONNECTED[1],n25_carry__0_n_7}),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,n25_carry__0_i_1__1_n_0,n25_carry__0_i_2__1_n_0}),
        .O({NLW_n25_carry__0_O_UNCONNECTED[7:2],n25_carry__0_n_14,n25_carry__0_n_15}),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,n25_carry__0_i_3__0_n_0,n25_carry__0_i_4__1_n_0}));
  LUT3 #(
    .INIT(8'h40)) 
    n25_carry__0_i_1__1
       (.I0(\n4_reg_n_0_[7] ),
        .I1(B),
        .I2(\n4_reg_n_0_[6] ),
        .O(n25_carry__0_i_1__1_n_0));
  LUT4 #(
    .INIT(16'h80C8)) 
    n25_carry__0_i_2__1
       (.I0(\n4_reg_n_0_[5] ),
        .I1(B),
        .I2(\n4_reg_n_0_[6] ),
        .I3(\n4_reg_n_0_[7] ),
        .O(n25_carry__0_i_2__1_n_0));
  LUT3 #(
    .INIT(8'h37)) 
    n25_carry__0_i_3__0
       (.I0(\n4_reg_n_0_[6] ),
        .I1(B),
        .I2(\n4_reg_n_0_[7] ),
        .O(n25_carry__0_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h4FDF)) 
    n25_carry__0_i_4__1
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(B),
        .I3(\n4_reg_n_0_[7] ),
        .O(n25_carry__0_i_4__1_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n25_carry_i_10__1
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(B),
        .I3(\n4_reg_n_0_[3] ),
        .I4(\n4_reg_n_0_[5] ),
        .O(n25_carry_i_10__1_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n25_carry_i_11__1
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(B),
        .I3(\n4_reg_n_0_[2] ),
        .I4(\n4_reg_n_0_[4] ),
        .O(n25_carry_i_11__1_n_0));
  LUT5 #(
    .INIT(32'h66009600)) 
    n25_carry_i_12__1
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[1] ),
        .I3(B),
        .I4(\n4_reg_n_0_[0] ),
        .O(n25_carry_i_12__1_n_0));
  LUT4 #(
    .INIT(16'h9060)) 
    n25_carry_i_13__0
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(B),
        .I3(\n4_reg_n_0_[2] ),
        .O(n25_carry_i_13__0_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n25_carry_i_14__0
       (.I0(\n4_reg_n_0_[1] ),
        .I1(B),
        .I2(\n4_reg_n_0_[0] ),
        .O(n25_carry_i_14__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25_carry_i_15__0
       (.I0(B),
        .I1(\n4_reg_n_0_[0] ),
        .O(n25_carry_i_15__0_n_0));
  (* HLUTNM = "lutpair108" *) 
  LUT4 #(
    .INIT(16'hC880)) 
    n25_carry_i_1__1
       (.I0(\n4_reg_n_0_[4] ),
        .I1(B),
        .I2(\n4_reg_n_0_[5] ),
        .I3(\n4_reg_n_0_[6] ),
        .O(n25_carry_i_1__1_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n25_carry_i_2__1
       (.I0(\n4_reg_n_0_[3] ),
        .I1(B),
        .I2(\n4_reg_n_0_[4] ),
        .I3(\n4_reg_n_0_[5] ),
        .O(n25_carry_i_2__1_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n25_carry_i_3__1
       (.I0(\n4_reg_n_0_[2] ),
        .I1(B),
        .I2(\n4_reg_n_0_[3] ),
        .I3(\n4_reg_n_0_[4] ),
        .O(n25_carry_i_3__1_n_0));
  LUT4 #(
    .INIT(16'hC880)) 
    n25_carry_i_4__1
       (.I0(\n4_reg_n_0_[1] ),
        .I1(B),
        .I2(\n4_reg_n_0_[2] ),
        .I3(\n4_reg_n_0_[3] ),
        .O(n25_carry_i_4__1_n_0));
  LUT4 #(
    .INIT(16'h8448)) 
    n25_carry_i_5__1
       (.I0(\n4_reg_n_0_[2] ),
        .I1(B),
        .I2(\n4_reg_n_0_[1] ),
        .I3(\n4_reg_n_0_[3] ),
        .O(n25_carry_i_5__1_n_0));
  LUT3 #(
    .INIT(8'h48)) 
    n25_carry_i_6__1
       (.I0(\n4_reg_n_0_[1] ),
        .I1(B),
        .I2(\n4_reg_n_0_[0] ),
        .O(n25_carry_i_6__1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    n25_carry_i_7__0
       (.I0(B),
        .I1(\n4_reg_n_0_[1] ),
        .O(n25_carry_i_7__0_n_0));
  LUT5 #(
    .INIT(32'h95656595)) 
    n25_carry_i_8__0
       (.I0(n25_carry_i_1__1_n_0),
        .I1(\n4_reg_n_0_[6] ),
        .I2(B),
        .I3(\n4_reg_n_0_[5] ),
        .I4(\n4_reg_n_0_[7] ),
        .O(n25_carry_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h20B0D040)) 
    n25_carry_i_9__1
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[5] ),
        .I2(B),
        .I3(\n4_reg_n_0_[4] ),
        .I4(\n4_reg_n_0_[6] ),
        .O(n25_carry_i_9__1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[0]),
        .Q(n27[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[1]),
        .Q(n27[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[2]),
        .Q(n27[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[3]),
        .Q(n27[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[4]),
        .Q(n27[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[5]),
        .Q(n27[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[6]),
        .Q(n27[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[7]),
        .Q(n27[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[0]),
        .Q(n29[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[1]),
        .Q(n29[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[2]),
        .Q(n29[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[3]),
        .Q(n29[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[4]),
        .Q(n29[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[5]),
        .Q(n29[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[6]),
        .Q(n29[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[7]),
        .Q(n29[7]),
        .R(rst_i));
  LUT2 #(
    .INIT(4'h6)) 
    \n33[0]_i_1__7 
       (.I0(n29[0]),
        .I1(n10[0]),
        .O(n31[0]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[10]_i_1__7 
       (.I0(n21[2]),
        .I1(\n8_reg_n_0_[2] ),
        .I2(\n8_reg_n_0_[1] ),
        .I3(n21[1]),
        .I4(\n8_reg_n_0_[0] ),
        .I5(n21[0]),
        .O(\n33[10]_i_1__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[11]_i_1__7 
       (.I0(n21[3]),
        .I1(\n8_reg_n_0_[3] ),
        .I2(\n33[12]_i_2__7_n_0 ),
        .O(\n33[11]_i_1__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[12]_i_1__7 
       (.I0(n21[4]),
        .I1(\n8_reg_n_0_[4] ),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[3]),
        .I4(\n33[12]_i_2__7_n_0 ),
        .O(\n33[12]_i_1__7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[12]_i_2__7 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n33[12]_i_2__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[13]_i_1__7 
       (.I0(n21[5]),
        .I1(\n8_reg_n_0_[5] ),
        .I2(\n33[14]_i_2__7_n_0 ),
        .O(\n33[13]_i_1__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[14]_i_1__7 
       (.I0(n21[6]),
        .I1(\n8_reg_n_0_[6] ),
        .I2(\n8_reg_n_0_[5] ),
        .I3(n21[5]),
        .I4(\n33[14]_i_2__7_n_0 ),
        .O(\n33[14]_i_1__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[14]_i_2__7 
       (.I0(\n33[12]_i_2__7_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n33[14]_i_2__7_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[15]_i_1__7 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n33[15]_i_2__7_n_0 ),
        .O(n30));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[15]_i_2__7 
       (.I0(\n33[14]_i_2__7_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n33[15]_i_2__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[1]_i_1__7 
       (.I0(n29[1]),
        .I1(n10[1]),
        .I2(n10[0]),
        .I3(n29[0]),
        .O(n31[1]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[2]_i_1__7 
       (.I0(n29[2]),
        .I1(n10[2]),
        .I2(n10[1]),
        .I3(n29[1]),
        .I4(n10[0]),
        .I5(n29[0]),
        .O(\n33[2]_i_1__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[3]_i_1__7 
       (.I0(n29[3]),
        .I1(n10[3]),
        .I2(\n33[4]_i_2__7_n_0 ),
        .O(\n33[3]_i_1__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[4]_i_1__7 
       (.I0(n29[4]),
        .I1(n10[4]),
        .I2(n10[3]),
        .I3(n29[3]),
        .I4(\n33[4]_i_2__7_n_0 ),
        .O(\n33[4]_i_1__7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[4]_i_2__7 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n33[4]_i_2__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[5]_i_1__7 
       (.I0(n29[5]),
        .I1(n10[5]),
        .I2(\n33[6]_i_2__7_n_0 ),
        .O(\n33[5]_i_1__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[6]_i_1__7 
       (.I0(n29[6]),
        .I1(n10[6]),
        .I2(n10[5]),
        .I3(n29[5]),
        .I4(\n33[6]_i_2__7_n_0 ),
        .O(\n33[6]_i_1__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[6]_i_2__7 
       (.I0(\n33[4]_i_2__7_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n33[6]_i_2__7_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[7]_i_1__7 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n33[7]_i_2__7_n_0 ),
        .O(n31[7]));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[7]_i_2__7 
       (.I0(\n33[6]_i_2__7_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n33[7]_i_2__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[9]_i_1__7 
       (.I0(n21[1]),
        .I1(\n8_reg_n_0_[1] ),
        .I2(\n8_reg_n_0_[0] ),
        .I3(n21[0]),
        .O(\n33[9]_i_1__7_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[0]),
        .Q(i1[15]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[10]_i_1__7_n_0 ),
        .Q(i1[24]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[11]_i_1__7_n_0 ),
        .Q(i1[25]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[12]_i_1__7_n_0 ),
        .Q(i1[26]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[13]_i_1__7_n_0 ),
        .Q(i1[27]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[14]_i_1__7_n_0 ),
        .Q(i1[28]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n30),
        .Q(i1[29]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[1]),
        .Q(i1[16]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[2]_i_1__7_n_0 ),
        .Q(i1[17]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[3]_i_1__7_n_0 ),
        .Q(i1[18]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[4]_i_1__7_n_0 ),
        .Q(i1[19]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[5]_i_1__7_n_0 ),
        .Q(i1[20]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[6]_i_1__7_n_0 ),
        .Q(i1[21]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[7]),
        .Q(i1[22]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[9]_i_1__7_n_0 ),
        .Q(i1[23]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[10]_i_1__7 
       (.I0(\n8_reg_n_0_[1] ),
        .I1(n21[1]),
        .I2(n21[0]),
        .I3(\n8_reg_n_0_[0] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(n341_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[11]_i_1__7 
       (.I0(\n37[12]_i_2__7_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .O(n341_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[12]_i_1__7 
       (.I0(\n8_reg_n_0_[3] ),
        .I1(n21[3]),
        .I2(\n37[12]_i_2__7_n_0 ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(n341_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[12]_i_2__7 
       (.I0(\n8_reg_n_0_[0] ),
        .I1(n21[0]),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n37[12]_i_2__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[13]_i_1__7 
       (.I0(\n37[14]_i_2__7_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(n341_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[14]_i_1__7 
       (.I0(\n8_reg_n_0_[5] ),
        .I1(n21[5]),
        .I2(\n37[14]_i_2__7_n_0 ),
        .I3(n21[6]),
        .I4(\n8_reg_n_0_[6] ),
        .O(n341_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[14]_i_2__7 
       (.I0(\n37[12]_i_2__7_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n37[14]_i_2__7_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[15]_i_1__7 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n37[15]_i_2__7_n_0 ),
        .O(n341_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[15]_i_2__7 
       (.I0(\n37[14]_i_2__7_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n37[15]_i_2__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[1]_i_1__7 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .O(n350_out[1]));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[2]_i_1__7 
       (.I0(n10[1]),
        .I1(n29[1]),
        .I2(n29[0]),
        .I3(n10[0]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(n350_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[3]_i_1__7 
       (.I0(\n37[4]_i_2__7_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .O(n350_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[4]_i_1__7 
       (.I0(n10[3]),
        .I1(n29[3]),
        .I2(\n37[4]_i_2__7_n_0 ),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(n350_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[4]_i_2__7 
       (.I0(n10[0]),
        .I1(n29[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n37[4]_i_2__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[5]_i_1__7 
       (.I0(\n37[6]_i_2__7_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(n350_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[6]_i_1__7 
       (.I0(n10[5]),
        .I1(n29[5]),
        .I2(\n37[6]_i_2__7_n_0 ),
        .I3(n29[6]),
        .I4(n10[6]),
        .O(n350_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[6]_i_2__7 
       (.I0(\n37[4]_i_2__7_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n37[6]_i_2__7_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[7]_i_1__7 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n37[7]_i_2__7_n_0 ),
        .O(n350_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[7]_i_2__7 
       (.I0(\n37[6]_i_2__7_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n37[7]_i_2__7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n37[8]_i_1__4 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .O(n341_out[0]));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[9]_i_1__7 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .O(n341_out[1]));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[2]),
        .Q(i1[9]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[3]),
        .Q(i1[10]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[4]),
        .Q(i1[11]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[5]),
        .Q(i1[12]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[6]),
        .Q(i1[13]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[7]),
        .Q(i1[14]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[1]),
        .Q(i1[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[2]),
        .Q(i1[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[3]),
        .Q(i1[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[4]),
        .Q(i1[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[5]),
        .Q(i1[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[6]),
        .Q(i1[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[7]),
        .Q(i1[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[0]),
        .Q(i1[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[1]),
        .Q(i1[8]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n4_reg[7]_0 [0]),
        .Q(\n4_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n4_reg[7]_0 [1]),
        .Q(\n4_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n4_reg[7]_0 [2]),
        .Q(\n4_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n4_reg[7]_0 [3]),
        .Q(\n4_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n4_reg[7]_0 [4]),
        .Q(\n4_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n4_reg[7]_0 [5]),
        .Q(\n4_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n4_reg[7]_0 [6]),
        .Q(\n4_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n4_reg[7]_0 [7]),
        .Q(\n4_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2_2[0]),
        .Q(\n7_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2_2[1]),
        .Q(\n7_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2_2[2]),
        .Q(\n7_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2_2[3]),
        .Q(\n7_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2_2[4]),
        .Q(\n7_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2_2[5]),
        .Q(\n7_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2_2[6]),
        .Q(\n7_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2_2[7]),
        .Q(\n7_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[0] ),
        .Q(\n8_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[1] ),
        .Q(\n8_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[2] ),
        .Q(\n8_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[3] ),
        .Q(\n8_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[4] ),
        .Q(\n8_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[5] ),
        .Q(\n8_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[6] ),
        .Q(\n8_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[7] ),
        .Q(\n8_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[0] ),
        .Q(\n9_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[1] ),
        .Q(\n9_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[2] ),
        .Q(\n9_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[3] ),
        .Q(\n9_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[4] ),
        .Q(\n9_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[5] ),
        .Q(\n9_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[6] ),
        .Q(\n9_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[7] ),
        .Q(\n9_reg_n_0_[7] ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_4" *) 
module switch_elements_cf_fft_512_8_4
   (\n5_reg[0] ,
    \n5_reg[0]_0 ,
    clk_i,
    i2,
    i8,
    n22,
    enable_i,
    rst_i);
  output [7:0]\n5_reg[0] ;
  output [7:0]\n5_reg[0]_0 ;
  input clk_i;
  input [31:0]i2;
  input [0:0]i8;
  input n22;
  input [0:0]enable_i;
  input rst_i;

  wire clk_i;
  wire [0:0]enable_i;
  wire [31:0]i2;
  wire [0:0]i8;
  wire n22;
  wire [5:0]n2__0;
  wire [5:0]n3_reg;
  wire [7:0]\n5_reg[0] ;
  wire [7:0]\n5_reg[0]_0 ;
  wire \n6a_reg_n_0_[0] ;
  wire \n6a_reg_n_0_[1] ;
  wire \n6a_reg_n_0_[2] ;
  wire \n6a_reg_n_0_[3] ;
  wire \n6a_reg_n_0_[4] ;
  wire \n6a_reg_n_0_[5] ;
  wire n6m_reg_0_63_0_6_n_0;
  wire n6m_reg_0_63_0_6_n_1;
  wire n6m_reg_0_63_0_6_n_2;
  wire n6m_reg_0_63_0_6_n_3;
  wire n6m_reg_0_63_0_6_n_4;
  wire n6m_reg_0_63_0_6_n_5;
  wire n6m_reg_0_63_0_6_n_6;
  wire n6m_reg_0_63_14_20_n_0;
  wire n6m_reg_0_63_14_20_n_1;
  wire n6m_reg_0_63_14_20_n_2;
  wire n6m_reg_0_63_14_20_n_3;
  wire n6m_reg_0_63_14_20_n_4;
  wire n6m_reg_0_63_14_20_n_5;
  wire n6m_reg_0_63_14_20_n_6;
  wire n6m_reg_0_63_21_27_n_0;
  wire n6m_reg_0_63_21_27_n_1;
  wire n6m_reg_0_63_21_27_n_2;
  wire n6m_reg_0_63_21_27_n_3;
  wire n6m_reg_0_63_21_27_n_4;
  wire n6m_reg_0_63_21_27_n_5;
  wire n6m_reg_0_63_21_27_n_6;
  wire n6m_reg_0_63_28_31_n_0;
  wire n6m_reg_0_63_28_31_n_1;
  wire n6m_reg_0_63_28_31_n_2;
  wire n6m_reg_0_63_28_31_n_3;
  wire n6m_reg_0_63_7_13_n_0;
  wire n6m_reg_0_63_7_13_n_1;
  wire n6m_reg_0_63_7_13_n_2;
  wire n6m_reg_0_63_7_13_n_3;
  wire n6m_reg_0_63_7_13_n_4;
  wire n6m_reg_0_63_7_13_n_5;
  wire n6m_reg_0_63_7_13_n_6;
  wire [31:0]n8;
  wire [5:0]n8a_0;
  wire rst_i;
  wire NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED;
  wire NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED;
  wire NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED;

  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    n22__0_i_1__6
       (.I0(n8[14]),
        .I1(n6m_reg_0_63_14_20_n_0),
        .I2(i8),
        .I3(n8[30]),
        .I4(n22),
        .I5(n6m_reg_0_63_28_31_n_2),
        .O(\n5_reg[0]_0 [6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    n22__1_i_1__6
       (.I0(n8[13]),
        .I1(n6m_reg_0_63_7_13_n_6),
        .I2(i8),
        .I3(n8[29]),
        .I4(n22),
        .I5(n6m_reg_0_63_28_31_n_1),
        .O(\n5_reg[0]_0 [5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    n22__2_i_1__6
       (.I0(n8[12]),
        .I1(n6m_reg_0_63_7_13_n_5),
        .I2(i8),
        .I3(n8[28]),
        .I4(n22),
        .I5(n6m_reg_0_63_28_31_n_0),
        .O(\n5_reg[0]_0 [4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    n22__3_i_1__6
       (.I0(n8[11]),
        .I1(n6m_reg_0_63_7_13_n_4),
        .I2(i8),
        .I3(n8[27]),
        .I4(n22),
        .I5(n6m_reg_0_63_21_27_n_6),
        .O(\n5_reg[0]_0 [3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    n22__4_i_1__6
       (.I0(n8[10]),
        .I1(n6m_reg_0_63_7_13_n_3),
        .I2(i8),
        .I3(n8[26]),
        .I4(n22),
        .I5(n6m_reg_0_63_21_27_n_5),
        .O(\n5_reg[0]_0 [2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    n22__5_i_1__6
       (.I0(n8[9]),
        .I1(n6m_reg_0_63_7_13_n_2),
        .I2(i8),
        .I3(n8[25]),
        .I4(n22),
        .I5(n6m_reg_0_63_21_27_n_4),
        .O(\n5_reg[0]_0 [1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    n22__6_i_1__6
       (.I0(n8[8]),
        .I1(n6m_reg_0_63_7_13_n_1),
        .I2(i8),
        .I3(n8[24]),
        .I4(n22),
        .I5(n6m_reg_0_63_21_27_n_3),
        .O(\n5_reg[0]_0 [0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    n22_i_1__6
       (.I0(n8[15]),
        .I1(n6m_reg_0_63_14_20_n_1),
        .I2(i8),
        .I3(n8[31]),
        .I4(n22),
        .I5(n6m_reg_0_63_28_31_n_3),
        .O(\n5_reg[0]_0 [7]));
  LUT1 #(
    .INIT(2'h1)) 
    \n3[0]_i_1__16 
       (.I0(n3_reg[0]),
        .O(n2__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n3[1]_i_1__16 
       (.I0(n3_reg[0]),
        .I1(n3_reg[1]),
        .O(n2__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \n3[2]_i_1__16 
       (.I0(n3_reg[1]),
        .I1(n3_reg[0]),
        .I2(n3_reg[2]),
        .O(n2__0[2]));
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT4 #(
    .INIT(16'h7F80)) 
    \n3[3]_i_1__16 
       (.I0(n3_reg[2]),
        .I1(n3_reg[0]),
        .I2(n3_reg[1]),
        .I3(n3_reg[3]),
        .O(n2__0[3]));
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \n3[4]_i_1__16 
       (.I0(n3_reg[3]),
        .I1(n3_reg[1]),
        .I2(n3_reg[0]),
        .I3(n3_reg[2]),
        .I4(n3_reg[4]),
        .O(n2__0[4]));
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \n3[5]_i_1__16 
       (.I0(n3_reg[4]),
        .I1(n3_reg[2]),
        .I2(n3_reg[0]),
        .I3(n3_reg[1]),
        .I4(n3_reg[3]),
        .I5(n3_reg[5]),
        .O(n2__0[5]));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[0]),
        .Q(n3_reg[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[1]),
        .Q(n3_reg[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[2]),
        .Q(n3_reg[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[3]),
        .Q(n3_reg[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[4]),
        .Q(n3_reg[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n3_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2__0[5]),
        .Q(n3_reg[5]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \n4[0]_i_1__6 
       (.I0(n8[0]),
        .I1(n6m_reg_0_63_0_6_n_0),
        .I2(i8),
        .I3(n8[16]),
        .I4(n22),
        .I5(n6m_reg_0_63_14_20_n_2),
        .O(\n5_reg[0] [0]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \n4[1]_i_1__6 
       (.I0(n8[1]),
        .I1(n6m_reg_0_63_0_6_n_1),
        .I2(i8),
        .I3(n8[17]),
        .I4(n22),
        .I5(n6m_reg_0_63_14_20_n_3),
        .O(\n5_reg[0] [1]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \n4[2]_i_1__6 
       (.I0(n8[2]),
        .I1(n6m_reg_0_63_0_6_n_2),
        .I2(i8),
        .I3(n8[18]),
        .I4(n22),
        .I5(n6m_reg_0_63_14_20_n_4),
        .O(\n5_reg[0] [2]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \n4[3]_i_1__6 
       (.I0(n8[3]),
        .I1(n6m_reg_0_63_0_6_n_3),
        .I2(i8),
        .I3(n8[19]),
        .I4(n22),
        .I5(n6m_reg_0_63_14_20_n_5),
        .O(\n5_reg[0] [3]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \n4[4]_i_1__6 
       (.I0(n8[4]),
        .I1(n6m_reg_0_63_0_6_n_4),
        .I2(i8),
        .I3(n8[20]),
        .I4(n22),
        .I5(n6m_reg_0_63_14_20_n_6),
        .O(\n5_reg[0] [4]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \n4[5]_i_1__6 
       (.I0(n8[5]),
        .I1(n6m_reg_0_63_0_6_n_5),
        .I2(i8),
        .I3(n8[21]),
        .I4(n22),
        .I5(n6m_reg_0_63_21_27_n_0),
        .O(\n5_reg[0] [5]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \n4[6]_i_1__6 
       (.I0(n8[6]),
        .I1(n6m_reg_0_63_0_6_n_6),
        .I2(i8),
        .I3(n8[22]),
        .I4(n22),
        .I5(n6m_reg_0_63_21_27_n_1),
        .O(\n5_reg[0] [6]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \n4[7]_i_1__6 
       (.I0(n8[7]),
        .I1(n6m_reg_0_63_7_13_n_0),
        .I2(i8),
        .I3(n8[23]),
        .I4(n22),
        .I5(n6m_reg_0_63_21_27_n_2),
        .O(\n5_reg[0] [7]));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(\n6a_reg_n_0_[0] ),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(\n6a_reg_n_0_[1] ),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(\n6a_reg_n_0_[2] ),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(\n6a_reg_n_0_[3] ),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(\n6a_reg_n_0_[4] ),
        .R(1'b0));
  (* equivalent_register_removal = "no" *) 
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(\n6a_reg_n_0_[5] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[0]),
        .Q(n8a_0[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[1]),
        .Q(n8a_0[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[2]),
        .Q(n8a_0[2]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[3]),
        .Q(n8a_0[3]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[4]),
        .Q(n8a_0[4]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \n6a_reg_rep[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n3_reg[5]),
        .Q(n8a_0[5]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s14/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39908 n6m_reg_0_63_0_6
       (.ADDRA(n8a_0),
        .ADDRB(n8a_0),
        .ADDRC(n8a_0),
        .ADDRD(n8a_0),
        .ADDRE(n8a_0),
        .ADDRF(n8a_0),
        .ADDRG(n8a_0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[0]),
        .DIB(i2[1]),
        .DIC(i2[2]),
        .DID(i2[3]),
        .DIE(i2[4]),
        .DIF(i2[5]),
        .DIG(i2[6]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_0_6_n_0),
        .DOB(n6m_reg_0_63_0_6_n_1),
        .DOC(n6m_reg_0_63_0_6_n_2),
        .DOD(n6m_reg_0_63_0_6_n_3),
        .DOE(n6m_reg_0_63_0_6_n_4),
        .DOF(n6m_reg_0_63_0_6_n_5),
        .DOG(n6m_reg_0_63_0_6_n_6),
        .DOH(NLW_n6m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s14/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39909 n6m_reg_0_63_14_20
       (.ADDRA(n8a_0),
        .ADDRB(n8a_0),
        .ADDRC(n8a_0),
        .ADDRD(n8a_0),
        .ADDRE(n8a_0),
        .ADDRF(n8a_0),
        .ADDRG(n8a_0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[14]),
        .DIB(i2[15]),
        .DIC(i2[16]),
        .DID(i2[17]),
        .DIE(i2[18]),
        .DIF(i2[19]),
        .DIG(i2[20]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_14_20_n_0),
        .DOB(n6m_reg_0_63_14_20_n_1),
        .DOC(n6m_reg_0_63_14_20_n_2),
        .DOD(n6m_reg_0_63_14_20_n_3),
        .DOE(n6m_reg_0_63_14_20_n_4),
        .DOF(n6m_reg_0_63_14_20_n_5),
        .DOG(n6m_reg_0_63_14_20_n_6),
        .DOH(NLW_n6m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s14/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39910 n6m_reg_0_63_21_27
       (.ADDRA(n8a_0),
        .ADDRB(n8a_0),
        .ADDRC(n8a_0),
        .ADDRD(n8a_0),
        .ADDRE(n8a_0),
        .ADDRF(n8a_0),
        .ADDRG(n8a_0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[21]),
        .DIB(i2[22]),
        .DIC(i2[23]),
        .DID(i2[24]),
        .DIE(i2[25]),
        .DIF(i2[26]),
        .DIG(i2[27]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_21_27_n_0),
        .DOB(n6m_reg_0_63_21_27_n_1),
        .DOC(n6m_reg_0_63_21_27_n_2),
        .DOD(n6m_reg_0_63_21_27_n_3),
        .DOE(n6m_reg_0_63_21_27_n_4),
        .DOF(n6m_reg_0_63_21_27_n_5),
        .DOG(n6m_reg_0_63_21_27_n_6),
        .DOH(NLW_n6m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s14/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39911 n6m_reg_0_63_28_31
       (.ADDRA(n8a_0),
        .ADDRB(n8a_0),
        .ADDRC(n8a_0),
        .ADDRD(n8a_0),
        .ADDRE(n8a_0),
        .ADDRF(n8a_0),
        .ADDRG(n8a_0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[28]),
        .DIB(i2[29]),
        .DIC(i2[30]),
        .DID(i2[31]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_28_31_n_0),
        .DOB(n6m_reg_0_63_28_31_n_1),
        .DOC(n6m_reg_0_63_28_31_n_2),
        .DOD(n6m_reg_0_63_28_31_n_3),
        .DOE(NLW_n6m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n6m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n6m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n6m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s14/n6m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39912 n6m_reg_0_63_7_13
       (.ADDRA(n8a_0),
        .ADDRB(n8a_0),
        .ADDRC(n8a_0),
        .ADDRD(n8a_0),
        .ADDRE(n8a_0),
        .ADDRF(n8a_0),
        .ADDRG(n8a_0),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[7]),
        .DIB(i2[8]),
        .DIC(i2[9]),
        .DID(i2[10]),
        .DIE(i2[11]),
        .DIF(i2[12]),
        .DIG(i2[13]),
        .DIH(1'b0),
        .DOA(n6m_reg_0_63_7_13_n_0),
        .DOB(n6m_reg_0_63_7_13_n_1),
        .DOC(n6m_reg_0_63_7_13_n_2),
        .DOD(n6m_reg_0_63_7_13_n_3),
        .DOE(n6m_reg_0_63_7_13_n_4),
        .DOF(n6m_reg_0_63_7_13_n_5),
        .DOG(n6m_reg_0_63_7_13_n_6),
        .DOH(NLW_n6m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s14/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "6" *) 
  RAM64M8_HD39913 n8m_reg_0_63_0_6
       (.ADDRA({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRB({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRC({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRD({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRE({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRF({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRG({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[0]),
        .DIB(i2[1]),
        .DIC(i2[2]),
        .DID(i2[3]),
        .DIE(i2[4]),
        .DIF(i2[5]),
        .DIG(i2[6]),
        .DIH(1'b0),
        .DOA(n8[0]),
        .DOB(n8[1]),
        .DOC(n8[2]),
        .DOD(n8[3]),
        .DOE(n8[4]),
        .DOF(n8[5]),
        .DOG(n8[6]),
        .DOH(NLW_n8m_reg_0_63_0_6_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s14/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "14" *) 
  (* ram_slice_end = "20" *) 
  RAM64M8_HD39914 n8m_reg_0_63_14_20
       (.ADDRA({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRB({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRC({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRD({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRE({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRF({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRG({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[14]),
        .DIB(i2[15]),
        .DIC(i2[16]),
        .DID(i2[17]),
        .DIE(i2[18]),
        .DIF(i2[19]),
        .DIG(i2[20]),
        .DIH(1'b0),
        .DOA(n8[14]),
        .DOB(n8[15]),
        .DOC(n8[16]),
        .DOD(n8[17]),
        .DOE(n8[18]),
        .DOF(n8[19]),
        .DOG(n8[20]),
        .DOH(NLW_n8m_reg_0_63_14_20_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s14/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "21" *) 
  (* ram_slice_end = "27" *) 
  RAM64M8_HD39915 n8m_reg_0_63_21_27
       (.ADDRA({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRB({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRC({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRD({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRE({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRF({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRG({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[21]),
        .DIB(i2[22]),
        .DIC(i2[23]),
        .DID(i2[24]),
        .DIE(i2[25]),
        .DIF(i2[26]),
        .DIG(i2[27]),
        .DIH(1'b0),
        .DOA(n8[21]),
        .DOB(n8[22]),
        .DOC(n8[23]),
        .DOD(n8[24]),
        .DOE(n8[25]),
        .DOF(n8[26]),
        .DOG(n8[27]),
        .DOH(NLW_n8m_reg_0_63_21_27_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s14/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "28" *) 
  (* ram_slice_end = "31" *) 
  RAM64M8_HD39916 n8m_reg_0_63_28_31
       (.ADDRA({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRB({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRC({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRD({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRE({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRF({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRG({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[28]),
        .DIB(i2[29]),
        .DIC(i2[30]),
        .DID(i2[31]),
        .DIE(1'b0),
        .DIF(1'b0),
        .DIG(1'b0),
        .DIH(1'b0),
        .DOA(n8[28]),
        .DOB(n8[29]),
        .DOC(n8[30]),
        .DOD(n8[31]),
        .DOE(NLW_n8m_reg_0_63_28_31_DOE_UNCONNECTED),
        .DOF(NLW_n8m_reg_0_63_28_31_DOF_UNCONNECTED),
        .DOG(NLW_n8m_reg_0_63_28_31_DOG_UNCONNECTED),
        .DOH(NLW_n8m_reg_0_63_28_31_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
  (* INIT_A = "64'h0000000000000000" *) 
  (* INIT_B = "64'h0000000000000000" *) 
  (* INIT_C = "64'h0000000000000000" *) 
  (* INIT_D = "64'h0000000000000000" *) 
  (* INIT_E = "64'h0000000000000000" *) 
  (* INIT_F = "64'h0000000000000000" *) 
  (* INIT_G = "64'h0000000000000000" *) 
  (* INIT_H = "64'h0000000000000000" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  (* RTL_RAM_BITS = "4096" *) 
  (* RTL_RAM_NAME = "activity_blocks[0].switch3/s1/s3/s14/n8m" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "63" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "7" *) 
  (* ram_slice_end = "13" *) 
  RAM64M8_HD39917 n8m_reg_0_63_7_13
       (.ADDRA({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRB({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRC({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRD({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRE({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRF({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRG({\n6a_reg_n_0_[5] ,\n6a_reg_n_0_[4] ,\n6a_reg_n_0_[3] ,\n6a_reg_n_0_[2] ,\n6a_reg_n_0_[1] ,\n6a_reg_n_0_[0] }),
        .ADDRH({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .DIA(i2[7]),
        .DIB(i2[8]),
        .DIC(i2[9]),
        .DID(i2[10]),
        .DIE(i2[11]),
        .DIF(i2[12]),
        .DIG(i2[13]),
        .DIH(1'b0),
        .DOA(n8[7]),
        .DOB(n8[8]),
        .DOC(n8[9]),
        .DOD(n8[10]),
        .DOE(n8[11]),
        .DOF(n8[12]),
        .DOG(n8[13]),
        .DOH(NLW_n8m_reg_0_63_7_13_DOH_UNCONNECTED),
        .WCLK(clk_i),
        .WE(1'b0));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_5" *) 
module switch_elements_cf_fft_512_8_5
   (p_6_out,
    inf4_s,
    rst_i,
    enable_i,
    clk_i,
    enable_s,
    DOUTADOUT,
    n14__56_carry,
    i3,
    i2);
  output [31:0]p_6_out;
  output [31:0]inf4_s;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [31:0]enable_s;
  input [15:0]DOUTADOUT;
  input [15:0]n14__56_carry;
  input [15:0]i3;
  input [15:0]i2;

  wire [15:0]DOUTADOUT;
  wire clk_i;
  wire [0:0]enable_i;
  wire [31:0]enable_s;
  wire [15:0]i2;
  wire [15:0]i3;
  wire [31:0]inf4_s;
  wire [15:0]n14__56_carry;
  wire [31:0]p_6_out;
  wire rst_i;
  wire [15:0]s2_2;
  wire [15:0]s2_3;
  wire [15:0]s3_2;
  wire [15:0]s3_3;
  wire [15:0]s4_2;
  wire [15:0]s4_3;
  wire [15:0]s5_2;
  wire [15:0]s5_3;
  wire [15:0]s6_2;
  wire [15:0]s6_3;
  wire [15:0]s7_2;
  wire [15:0]s7_3;
  wire [15:0]s8_2;
  wire [15:0]s8_3;

  switch_elements_cf_fft_512_8_19 s1
       (.D(s2_2),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .enable_s(enable_s),
        .inf4_s(inf4_s),
        .p_6_out(p_6_out),
        .rst_i(rst_i),
        .s2_3(s2_3));
  switch_elements_cf_fft_512_8_17 s2
       (.D(s3_2),
        .DOUTADOUT(DOUTADOUT),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .\n9_reg[0] (s2_2),
        .rst_i(rst_i),
        .s2_3(s2_3),
        .s3_3(s3_3));
  switch_elements_cf_fft_512_8_15 s3
       (.D(s4_2),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .n14__56_carry(n14__56_carry),
        .\n9_reg[0] (s3_2),
        .rst_i(rst_i),
        .s3_3(s3_3),
        .s4_3(s4_3));
  switch_elements_cf_fft_512_8_13 s4
       (.D(s5_2),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .\n9_reg[0] (s4_2),
        .rst_i(rst_i),
        .s4_3(s4_3),
        .s5_3(s5_3));
  switch_elements_cf_fft_512_8_11 s5
       (.D(s6_2),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .\n9_reg[0] (s5_2),
        .rst_i(rst_i),
        .s5_3(s5_3),
        .s6_3(s6_3));
  switch_elements_cf_fft_512_8_9 s6
       (.D(s7_2),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .\n9_reg[0] (s6_2),
        .rst_i(rst_i),
        .s6_3(s6_3),
        .s7_3(s7_3));
  switch_elements_cf_fft_512_8_7 s7
       (.D(s8_2),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .\n9_reg[0] (s7_2),
        .rst_i(rst_i),
        .s7_3(s7_3),
        .s8_3(s8_3));
  switch_elements_cf_fft_512_8_6 s8
       (.D(s8_2),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .i2(i2),
        .i3(i3),
        .rst_i(rst_i),
        .s8_3(s8_3));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_6" *) 
module switch_elements_cf_fft_512_8_6
   (D,
    s8_3,
    rst_i,
    enable_i,
    clk_i,
    i3,
    i2);
  output [15:0]D;
  output [15:0]s8_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]i3;
  input [15:0]i2;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [15:0]i2;
  wire [15:0]i3;
  wire [0:0]i8;
  wire [15:0]n33;
  wire [15:1]n37;
  wire n4;
  wire rst_i;
  wire s28_n_0;
  wire [15:0]s8_3;

  switch_elements_cf_fft_512_8_37 s25
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .i2(i2),
        .i3(i3),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_31_0 s26
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i8(i8),
        .n4(n4),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_26 s27
       (.D(D),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .i8(i8),
        .\n1_reg[0] (s28_n_0),
        .n4(n4),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_27 s28
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .i8(i8),
        .\n9_reg[0]_0 (s28_n_0),
        .rst_i(rst_i),
        .s8_3(s8_3));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_7" *) 
module switch_elements_cf_fft_512_8_7
   (\n9_reg[0] ,
    s7_3,
    rst_i,
    enable_i,
    clk_i,
    s8_3,
    D);
  output [15:0]\n9_reg[0] ;
  output [15:0]s7_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]s8_3;
  input [15:0]D;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire [15:0]n33;
  wire [15:1]n37;
  wire n4;
  wire [15:0]\n9_reg[0] ;
  wire rst_i;
  wire s29_n_0;
  wire [15:0]s7_3;
  wire [15:0]s8_3;

  switch_elements_cf_fft_512_8_31_1 s25
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i8(i8),
        .n4(n4),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_8 s26
       (.D(D),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .rst_i(rst_i),
        .s8_3(s8_3));
  switch_elements_cf_fft_512_8_26_2 s28
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .i8(i8),
        .\n1_reg[0] (s29_n_0),
        .n4(n4),
        .\n9_reg[0] (\n9_reg[0] ),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_27_3 s29
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .i8(i8),
        .\n9_reg[0]_0 (s29_n_0),
        .rst_i(rst_i),
        .s7_3(s7_3));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_8" *) 
module switch_elements_cf_fft_512_8_8
   (i1,
    rst_i,
    enable_i,
    clk_i,
    s8_3,
    D);
  output [29:0]i1;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]s8_3;
  input [15:0]D;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [29:0]i1;
  wire [7:0]n10;
  wire [7:0]n15;
  wire \n16[3]_i_10_n_0 ;
  wire \n16[3]_i_11_n_0 ;
  wire \n16[3]_i_12_n_0 ;
  wire \n16[3]_i_13_n_0 ;
  wire \n16[3]_i_14__1_n_0 ;
  wire \n16[3]_i_15__1_n_0 ;
  wire \n16[3]_i_16_n_0 ;
  wire \n16[3]_i_18_n_0 ;
  wire \n16[3]_i_19_n_0 ;
  wire \n16[3]_i_20_n_0 ;
  wire \n16[3]_i_21_n_0 ;
  wire \n16[3]_i_22_n_0 ;
  wire \n16[3]_i_23__1_n_0 ;
  wire \n16[3]_i_24__1_n_0 ;
  wire \n16[3]_i_25__1_n_0 ;
  wire \n16[3]_i_26__1_n_0 ;
  wire \n16[3]_i_27_n_0 ;
  wire \n16[3]_i_28__1_n_0 ;
  wire \n16[3]_i_2_n_0 ;
  wire \n16[3]_i_3_n_0 ;
  wire \n16[3]_i_4_n_0 ;
  wire \n16[3]_i_5_n_0 ;
  wire \n16[3]_i_6__1_n_0 ;
  wire \n16[3]_i_7_n_0 ;
  wire \n16[3]_i_8_n_0 ;
  wire \n16[3]_i_9_n_0 ;
  wire \n16[7]_i_13__1_n_0 ;
  wire \n16[7]_i_14_n_0 ;
  wire \n16[7]_i_15__1_n_0 ;
  wire \n16[7]_i_16__1_n_0 ;
  wire \n16[7]_i_17_n_0 ;
  wire \n16[7]_i_18_n_0 ;
  wire \n16[7]_i_19__1_n_0 ;
  wire \n16[7]_i_20__1_n_0 ;
  wire \n16[7]_i_21__1_n_0 ;
  wire \n16[7]_i_22_n_0 ;
  wire \n16[7]_i_23__1_n_0 ;
  wire \n16[7]_i_24_n_0 ;
  wire \n16[7]_i_25_n_0 ;
  wire \n16[7]_i_26_n_0 ;
  wire \n16[7]_i_27_n_0 ;
  wire \n16[7]_i_28_n_0 ;
  wire \n16[7]_i_29__1_n_0 ;
  wire \n16[7]_i_2_n_0 ;
  wire \n16[7]_i_30__1_n_0 ;
  wire \n16[7]_i_31__1_n_0 ;
  wire \n16[7]_i_32__1_n_0 ;
  wire \n16[7]_i_33_n_0 ;
  wire \n16[7]_i_34__1_n_0 ;
  wire \n16[7]_i_35__1_n_0 ;
  wire \n16[7]_i_36_n_0 ;
  wire \n16[7]_i_37__1_n_0 ;
  wire \n16[7]_i_38__1_n_0 ;
  wire \n16[7]_i_3_n_0 ;
  wire \n16[7]_i_4_n_0 ;
  wire \n16[7]_i_5__1_n_0 ;
  wire \n16[7]_i_6__1_n_0 ;
  wire \n16[7]_i_7__1_n_0 ;
  wire \n16[7]_i_8_n_0 ;
  wire \n16_reg[3]_i_17_n_0 ;
  wire \n16_reg[3]_i_17_n_1 ;
  wire \n16_reg[3]_i_17_n_10 ;
  wire \n16_reg[3]_i_17_n_11 ;
  wire \n16_reg[3]_i_17_n_12 ;
  wire \n16_reg[3]_i_17_n_15 ;
  wire \n16_reg[3]_i_17_n_2 ;
  wire \n16_reg[3]_i_17_n_3 ;
  wire \n16_reg[3]_i_17_n_4 ;
  wire \n16_reg[3]_i_17_n_5 ;
  wire \n16_reg[3]_i_17_n_6 ;
  wire \n16_reg[3]_i_17_n_7 ;
  wire \n16_reg[3]_i_17_n_8 ;
  wire \n16_reg[3]_i_17_n_9 ;
  wire \n16_reg[3]_i_1_n_0 ;
  wire \n16_reg[3]_i_1_n_1 ;
  wire \n16_reg[3]_i_1_n_2 ;
  wire \n16_reg[3]_i_1_n_3 ;
  wire \n16_reg[3]_i_1_n_4 ;
  wire \n16_reg[3]_i_1_n_5 ;
  wire \n16_reg[3]_i_1_n_6 ;
  wire \n16_reg[3]_i_1_n_7 ;
  wire \n16_reg[7]_i_10_n_1 ;
  wire \n16_reg[7]_i_10_n_10 ;
  wire \n16_reg[7]_i_10_n_11 ;
  wire \n16_reg[7]_i_10_n_12 ;
  wire \n16_reg[7]_i_10_n_13 ;
  wire \n16_reg[7]_i_10_n_14 ;
  wire \n16_reg[7]_i_10_n_15 ;
  wire \n16_reg[7]_i_10_n_2 ;
  wire \n16_reg[7]_i_10_n_3 ;
  wire \n16_reg[7]_i_10_n_4 ;
  wire \n16_reg[7]_i_10_n_5 ;
  wire \n16_reg[7]_i_10_n_6 ;
  wire \n16_reg[7]_i_10_n_7 ;
  wire \n16_reg[7]_i_10_n_8 ;
  wire \n16_reg[7]_i_10_n_9 ;
  wire \n16_reg[7]_i_11_n_0 ;
  wire \n16_reg[7]_i_11_n_1 ;
  wire \n16_reg[7]_i_11_n_10 ;
  wire \n16_reg[7]_i_11_n_11 ;
  wire \n16_reg[7]_i_11_n_12 ;
  wire \n16_reg[7]_i_11_n_13 ;
  wire \n16_reg[7]_i_11_n_14 ;
  wire \n16_reg[7]_i_11_n_2 ;
  wire \n16_reg[7]_i_11_n_3 ;
  wire \n16_reg[7]_i_11_n_4 ;
  wire \n16_reg[7]_i_11_n_5 ;
  wire \n16_reg[7]_i_11_n_6 ;
  wire \n16_reg[7]_i_11_n_7 ;
  wire \n16_reg[7]_i_11_n_8 ;
  wire \n16_reg[7]_i_11_n_9 ;
  wire \n16_reg[7]_i_12_n_14 ;
  wire \n16_reg[7]_i_12_n_15 ;
  wire \n16_reg[7]_i_12_n_5 ;
  wire \n16_reg[7]_i_12_n_7 ;
  wire \n16_reg[7]_i_1_n_5 ;
  wire \n16_reg[7]_i_1_n_6 ;
  wire \n16_reg[7]_i_1_n_7 ;
  wire \n16_reg[7]_i_9_n_14 ;
  wire \n16_reg[7]_i_9_n_15 ;
  wire \n16_reg[7]_i_9_n_5 ;
  wire \n16_reg[7]_i_9_n_7 ;
  wire \n16_reg_n_0_[0] ;
  wire \n16_reg_n_0_[1] ;
  wire \n16_reg_n_0_[2] ;
  wire \n16_reg_n_0_[3] ;
  wire \n16_reg_n_0_[4] ;
  wire \n16_reg_n_0_[5] ;
  wire \n16_reg_n_0_[6] ;
  wire \n16_reg_n_0_[7] ;
  wire \n1_reg_n_0_[0] ;
  wire \n1_reg_n_0_[1] ;
  wire \n1_reg_n_0_[2] ;
  wire \n1_reg_n_0_[3] ;
  wire \n1_reg_n_0_[4] ;
  wire \n1_reg_n_0_[5] ;
  wire \n1_reg_n_0_[6] ;
  wire \n1_reg_n_0_[7] ;
  wire [7:0]n2;
  wire [7:0]n202_out;
  wire [7:0]n21;
  wire \n21[7]_i_2__1_n_0 ;
  wire \n21[7]_i_3__1_n_0 ;
  wire \n21[7]_i_4__1_n_0 ;
  wire \n21[7]_i_5__1_n_0 ;
  wire \n21[7]_i_6__1_n_0 ;
  wire \n21[7]_i_7__1_n_0 ;
  wire \n21[7]_i_8__1_n_0 ;
  wire \n21[7]_i_9__1_n_0 ;
  wire \n21_reg[7]_i_1__1_n_1 ;
  wire \n21_reg[7]_i_1__1_n_2 ;
  wire \n21_reg[7]_i_1__1_n_3 ;
  wire \n21_reg[7]_i_1__1_n_4 ;
  wire \n21_reg[7]_i_1__1_n_5 ;
  wire \n21_reg[7]_i_1__1_n_6 ;
  wire \n21_reg[7]_i_1__1_n_7 ;
  wire n22__0_n_0;
  wire n22__1_n_0;
  wire n22__2_n_0;
  wire n22__3_n_0;
  wire n22__4_n_0;
  wire n22__5_n_0;
  wire n22__6_n_0;
  wire n22_n_0;
  wire [7:0]n26;
  wire [7:0]n27;
  wire \n27[3]_i_10_n_0 ;
  wire \n27[3]_i_11_n_0 ;
  wire \n27[3]_i_12_n_0 ;
  wire \n27[3]_i_13_n_0 ;
  wire \n27[3]_i_14__1_n_0 ;
  wire \n27[3]_i_15__1_n_0 ;
  wire \n27[3]_i_16_n_0 ;
  wire \n27[3]_i_18_n_0 ;
  wire \n27[3]_i_19_n_0 ;
  wire \n27[3]_i_20_n_0 ;
  wire \n27[3]_i_21_n_0 ;
  wire \n27[3]_i_22_n_0 ;
  wire \n27[3]_i_23__1_n_0 ;
  wire \n27[3]_i_24__1_n_0 ;
  wire \n27[3]_i_25__1_n_0 ;
  wire \n27[3]_i_26__1_n_0 ;
  wire \n27[3]_i_27_n_0 ;
  wire \n27[3]_i_28__1_n_0 ;
  wire \n27[3]_i_2_n_0 ;
  wire \n27[3]_i_3_n_0 ;
  wire \n27[3]_i_4_n_0 ;
  wire \n27[3]_i_5_n_0 ;
  wire \n27[3]_i_6__1_n_0 ;
  wire \n27[3]_i_7_n_0 ;
  wire \n27[3]_i_8_n_0 ;
  wire \n27[3]_i_9_n_0 ;
  wire \n27[7]_i_13__1_n_0 ;
  wire \n27[7]_i_14_n_0 ;
  wire \n27[7]_i_15__1_n_0 ;
  wire \n27[7]_i_16__1_n_0 ;
  wire \n27[7]_i_17_n_0 ;
  wire \n27[7]_i_18_n_0 ;
  wire \n27[7]_i_19__1_n_0 ;
  wire \n27[7]_i_20__1_n_0 ;
  wire \n27[7]_i_21__1_n_0 ;
  wire \n27[7]_i_22_n_0 ;
  wire \n27[7]_i_23__1_n_0 ;
  wire \n27[7]_i_24_n_0 ;
  wire \n27[7]_i_25_n_0 ;
  wire \n27[7]_i_26_n_0 ;
  wire \n27[7]_i_27_n_0 ;
  wire \n27[7]_i_28_n_0 ;
  wire \n27[7]_i_29__1_n_0 ;
  wire \n27[7]_i_2_n_0 ;
  wire \n27[7]_i_30__1_n_0 ;
  wire \n27[7]_i_31__1_n_0 ;
  wire \n27[7]_i_32__1_n_0 ;
  wire \n27[7]_i_33_n_0 ;
  wire \n27[7]_i_34__1_n_0 ;
  wire \n27[7]_i_35__1_n_0 ;
  wire \n27[7]_i_36_n_0 ;
  wire \n27[7]_i_37__1_n_0 ;
  wire \n27[7]_i_38__1_n_0 ;
  wire \n27[7]_i_3_n_0 ;
  wire \n27[7]_i_4_n_0 ;
  wire \n27[7]_i_5__1_n_0 ;
  wire \n27[7]_i_6__1_n_0 ;
  wire \n27[7]_i_7__1_n_0 ;
  wire \n27[7]_i_8_n_0 ;
  wire \n27_reg[3]_i_17_n_0 ;
  wire \n27_reg[3]_i_17_n_1 ;
  wire \n27_reg[3]_i_17_n_10 ;
  wire \n27_reg[3]_i_17_n_11 ;
  wire \n27_reg[3]_i_17_n_12 ;
  wire \n27_reg[3]_i_17_n_15 ;
  wire \n27_reg[3]_i_17_n_2 ;
  wire \n27_reg[3]_i_17_n_3 ;
  wire \n27_reg[3]_i_17_n_4 ;
  wire \n27_reg[3]_i_17_n_5 ;
  wire \n27_reg[3]_i_17_n_6 ;
  wire \n27_reg[3]_i_17_n_7 ;
  wire \n27_reg[3]_i_17_n_8 ;
  wire \n27_reg[3]_i_17_n_9 ;
  wire \n27_reg[3]_i_1_n_0 ;
  wire \n27_reg[3]_i_1_n_1 ;
  wire \n27_reg[3]_i_1_n_2 ;
  wire \n27_reg[3]_i_1_n_3 ;
  wire \n27_reg[3]_i_1_n_4 ;
  wire \n27_reg[3]_i_1_n_5 ;
  wire \n27_reg[3]_i_1_n_6 ;
  wire \n27_reg[3]_i_1_n_7 ;
  wire \n27_reg[7]_i_10_n_1 ;
  wire \n27_reg[7]_i_10_n_10 ;
  wire \n27_reg[7]_i_10_n_11 ;
  wire \n27_reg[7]_i_10_n_12 ;
  wire \n27_reg[7]_i_10_n_13 ;
  wire \n27_reg[7]_i_10_n_14 ;
  wire \n27_reg[7]_i_10_n_15 ;
  wire \n27_reg[7]_i_10_n_2 ;
  wire \n27_reg[7]_i_10_n_3 ;
  wire \n27_reg[7]_i_10_n_4 ;
  wire \n27_reg[7]_i_10_n_5 ;
  wire \n27_reg[7]_i_10_n_6 ;
  wire \n27_reg[7]_i_10_n_7 ;
  wire \n27_reg[7]_i_10_n_8 ;
  wire \n27_reg[7]_i_10_n_9 ;
  wire \n27_reg[7]_i_11_n_0 ;
  wire \n27_reg[7]_i_11_n_1 ;
  wire \n27_reg[7]_i_11_n_10 ;
  wire \n27_reg[7]_i_11_n_11 ;
  wire \n27_reg[7]_i_11_n_12 ;
  wire \n27_reg[7]_i_11_n_13 ;
  wire \n27_reg[7]_i_11_n_14 ;
  wire \n27_reg[7]_i_11_n_2 ;
  wire \n27_reg[7]_i_11_n_3 ;
  wire \n27_reg[7]_i_11_n_4 ;
  wire \n27_reg[7]_i_11_n_5 ;
  wire \n27_reg[7]_i_11_n_6 ;
  wire \n27_reg[7]_i_11_n_7 ;
  wire \n27_reg[7]_i_11_n_8 ;
  wire \n27_reg[7]_i_11_n_9 ;
  wire \n27_reg[7]_i_12_n_14 ;
  wire \n27_reg[7]_i_12_n_15 ;
  wire \n27_reg[7]_i_12_n_5 ;
  wire \n27_reg[7]_i_12_n_7 ;
  wire \n27_reg[7]_i_1_n_5 ;
  wire \n27_reg[7]_i_1_n_6 ;
  wire \n27_reg[7]_i_1_n_7 ;
  wire \n27_reg[7]_i_9_n_14 ;
  wire \n27_reg[7]_i_9_n_15 ;
  wire \n27_reg[7]_i_9_n_5 ;
  wire \n27_reg[7]_i_9_n_7 ;
  wire [7:0]n29;
  wire [7:7]n30;
  wire [7:0]n31;
  wire \n33[10]_i_1__5_n_0 ;
  wire \n33[11]_i_1__5_n_0 ;
  wire \n33[12]_i_1__5_n_0 ;
  wire \n33[12]_i_2__5_n_0 ;
  wire \n33[13]_i_1__5_n_0 ;
  wire \n33[14]_i_1__5_n_0 ;
  wire \n33[14]_i_2__5_n_0 ;
  wire \n33[15]_i_2__5_n_0 ;
  wire \n33[2]_i_1__5_n_0 ;
  wire \n33[3]_i_1__5_n_0 ;
  wire \n33[4]_i_1__5_n_0 ;
  wire \n33[4]_i_2__5_n_0 ;
  wire \n33[5]_i_1__5_n_0 ;
  wire \n33[6]_i_1__5_n_0 ;
  wire \n33[6]_i_2__5_n_0 ;
  wire \n33[7]_i_2__5_n_0 ;
  wire \n33[9]_i_1__5_n_0 ;
  wire [7:0]n341_out;
  wire [7:1]n350_out;
  wire \n37[12]_i_2__5_n_0 ;
  wire \n37[14]_i_2__5_n_0 ;
  wire \n37[15]_i_2__5_n_0 ;
  wire \n37[4]_i_2__5_n_0 ;
  wire \n37[6]_i_2__5_n_0 ;
  wire \n37[7]_i_2__5_n_0 ;
  wire \n4_reg_n_0_[0] ;
  wire \n4_reg_n_0_[1] ;
  wire \n4_reg_n_0_[2] ;
  wire \n4_reg_n_0_[3] ;
  wire \n4_reg_n_0_[4] ;
  wire \n4_reg_n_0_[5] ;
  wire \n4_reg_n_0_[6] ;
  wire \n4_reg_n_0_[7] ;
  wire \n7_reg_n_0_[0] ;
  wire \n7_reg_n_0_[1] ;
  wire \n7_reg_n_0_[2] ;
  wire \n7_reg_n_0_[3] ;
  wire \n7_reg_n_0_[4] ;
  wire \n7_reg_n_0_[5] ;
  wire \n7_reg_n_0_[6] ;
  wire \n7_reg_n_0_[7] ;
  wire \n8_reg_n_0_[0] ;
  wire \n8_reg_n_0_[1] ;
  wire \n8_reg_n_0_[2] ;
  wire \n8_reg_n_0_[3] ;
  wire \n8_reg_n_0_[4] ;
  wire \n8_reg_n_0_[5] ;
  wire \n8_reg_n_0_[6] ;
  wire \n8_reg_n_0_[7] ;
  wire \n9_reg_n_0_[0] ;
  wire \n9_reg_n_0_[1] ;
  wire \n9_reg_n_0_[2] ;
  wire \n9_reg_n_0_[3] ;
  wire \n9_reg_n_0_[4] ;
  wire \n9_reg_n_0_[5] ;
  wire \n9_reg_n_0_[6] ;
  wire \n9_reg_n_0_[7] ;
  wire rst_i;
  wire [15:0]s8_3;
  wire [3:0]\NLW_n16_reg[3]_i_1_O_UNCONNECTED ;
  wire [2:1]\NLW_n16_reg[3]_i_17_O_UNCONNECTED ;
  wire [7:3]\NLW_n16_reg[7]_i_1_CO_UNCONNECTED ;
  wire [7:4]\NLW_n16_reg[7]_i_1_O_UNCONNECTED ;
  wire [7:7]\NLW_n16_reg[7]_i_10_CO_UNCONNECTED ;
  wire [0:0]\NLW_n16_reg[7]_i_11_O_UNCONNECTED ;
  wire [7:1]\NLW_n16_reg[7]_i_12_CO_UNCONNECTED ;
  wire [7:2]\NLW_n16_reg[7]_i_12_O_UNCONNECTED ;
  wire [7:1]\NLW_n16_reg[7]_i_9_CO_UNCONNECTED ;
  wire [7:2]\NLW_n16_reg[7]_i_9_O_UNCONNECTED ;
  wire [7:7]\NLW_n21_reg[7]_i_1__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_n27_reg[3]_i_1_O_UNCONNECTED ;
  wire [2:1]\NLW_n27_reg[3]_i_17_O_UNCONNECTED ;
  wire [7:3]\NLW_n27_reg[7]_i_1_CO_UNCONNECTED ;
  wire [7:4]\NLW_n27_reg[7]_i_1_O_UNCONNECTED ;
  wire [7:7]\NLW_n27_reg[7]_i_10_CO_UNCONNECTED ;
  wire [0:0]\NLW_n27_reg[7]_i_11_O_UNCONNECTED ;
  wire [7:1]\NLW_n27_reg[7]_i_12_CO_UNCONNECTED ;
  wire [7:2]\NLW_n27_reg[7]_i_12_O_UNCONNECTED ;
  wire [7:1]\NLW_n27_reg[7]_i_9_CO_UNCONNECTED ;
  wire [7:2]\NLW_n27_reg[7]_i_9_O_UNCONNECTED ;

  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[0] ),
        .Q(n10[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[1] ),
        .Q(n10[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[2] ),
        .Q(n10[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[3] ),
        .Q(n10[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[4] ),
        .Q(n10[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[5] ),
        .Q(n10[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[6] ),
        .Q(n10[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n10_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n9_reg_n_0_[7] ),
        .Q(n10[7]),
        .R(rst_i));
  (* HLUTNM = "lutpair63" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_10 
       (.I0(\n16_reg[7]_i_10_n_13 ),
        .I1(\n16_reg[7]_i_11_n_9 ),
        .I2(\n16_reg[7]_i_12_n_14 ),
        .I3(\n16[3]_i_3_n_0 ),
        .O(\n16[3]_i_10_n_0 ));
  (* HLUTNM = "lutpair62" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_11 
       (.I0(\n16_reg[7]_i_10_n_14 ),
        .I1(\n16_reg[7]_i_11_n_10 ),
        .I2(\n16_reg[7]_i_12_n_15 ),
        .I3(\n16[3]_i_4_n_0 ),
        .O(\n16[3]_i_11_n_0 ));
  (* HLUTNM = "lutpair61" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_12 
       (.I0(\n16_reg[7]_i_10_n_15 ),
        .I1(\n16_reg[7]_i_11_n_11 ),
        .I2(\n16_reg[3]_i_17_n_8 ),
        .I3(\n16[3]_i_5_n_0 ),
        .O(\n16[3]_i_12_n_0 ));
  (* HLUTNM = "lutpair60" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_13 
       (.I0(\n16_reg[3]_i_17_n_15 ),
        .I1(\n16_reg[7]_i_11_n_12 ),
        .I2(\n16_reg[3]_i_17_n_9 ),
        .I3(\n16[3]_i_6__1_n_0 ),
        .O(\n16[3]_i_13_n_0 ));
  (* HLUTNM = "lutpair103" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n16[3]_i_14__1 
       (.I0(\n16_reg[7]_i_11_n_13 ),
        .I1(\n16_reg[3]_i_17_n_10 ),
        .I2(\n16_reg[3]_i_17_n_11 ),
        .I3(\n16_reg[7]_i_11_n_14 ),
        .O(\n16[3]_i_14__1_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n16[3]_i_15__1 
       (.I0(\n16_reg[3]_i_17_n_12 ),
        .I1(n22__6_n_0),
        .I2(\n16_reg[7]_i_11_n_14 ),
        .I3(\n16_reg[3]_i_17_n_11 ),
        .O(\n16[3]_i_15__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n16[3]_i_16 
       (.I0(\n16_reg[3]_i_17_n_12 ),
        .I1(n22__6_n_0),
        .O(\n16[3]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_18 
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(n22__1_n_0),
        .O(\n16[3]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_19 
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__2_n_0),
        .O(\n16[3]_i_19_n_0 ));
  (* HLUTNM = "lutpair63" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_2 
       (.I0(\n16_reg[7]_i_10_n_13 ),
        .I1(\n16_reg[7]_i_11_n_9 ),
        .I2(\n16_reg[7]_i_12_n_14 ),
        .O(\n16[3]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_20 
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(n22__3_n_0),
        .O(\n16[3]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n16[3]_i_21 
       (.I0(n22__4_n_0),
        .I1(n22__5_n_0),
        .I2(n22__3_n_0),
        .O(\n16[3]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h9669)) 
    \n16[3]_i_22 
       (.I0(\n16[7]_i_23__1_n_0 ),
        .I1(n22__0_n_0),
        .I2(n22__1_n_0),
        .I3(n22_n_0),
        .O(\n16[3]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[3]_i_23__1 
       (.I0(n22__3_n_0),
        .I1(n22__1_n_0),
        .I2(n22__2_n_0),
        .I3(n22__0_n_0),
        .O(\n16[3]_i_23__1_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[3]_i_24__1 
       (.I0(n22__4_n_0),
        .I1(n22__2_n_0),
        .I2(n22__3_n_0),
        .I3(n22__1_n_0),
        .O(\n16[3]_i_24__1_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[3]_i_25__1 
       (.I0(n22__5_n_0),
        .I1(n22__3_n_0),
        .I2(n22__4_n_0),
        .I3(n22__2_n_0),
        .O(\n16[3]_i_25__1_n_0 ));
  LUT4 #(
    .INIT(16'h6696)) 
    \n16[3]_i_26__1 
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__5_n_0),
        .I3(n22__6_n_0),
        .O(\n16[3]_i_26__1_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n16[3]_i_27 
       (.I0(n22__6_n_0),
        .I1(n22__5_n_0),
        .I2(n22__4_n_0),
        .O(\n16[3]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n16[3]_i_28__1 
       (.I0(n22__5_n_0),
        .I1(n22__6_n_0),
        .O(\n16[3]_i_28__1_n_0 ));
  (* HLUTNM = "lutpair62" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_3 
       (.I0(\n16_reg[7]_i_10_n_14 ),
        .I1(\n16_reg[7]_i_11_n_10 ),
        .I2(\n16_reg[7]_i_12_n_15 ),
        .O(\n16[3]_i_3_n_0 ));
  (* HLUTNM = "lutpair61" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_4 
       (.I0(\n16_reg[7]_i_10_n_15 ),
        .I1(\n16_reg[7]_i_11_n_11 ),
        .I2(\n16_reg[3]_i_17_n_8 ),
        .O(\n16[3]_i_4_n_0 ));
  (* HLUTNM = "lutpair60" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[3]_i_5 
       (.I0(\n16_reg[3]_i_17_n_15 ),
        .I1(\n16_reg[7]_i_11_n_12 ),
        .I2(\n16_reg[3]_i_17_n_9 ),
        .O(\n16[3]_i_5_n_0 ));
  (* HLUTNM = "lutpair103" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \n16[3]_i_6__1 
       (.I0(\n16_reg[7]_i_11_n_13 ),
        .I1(\n16_reg[3]_i_17_n_10 ),
        .O(\n16[3]_i_6__1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n16[3]_i_7 
       (.I0(\n16_reg[3]_i_17_n_11 ),
        .I1(\n16_reg[7]_i_11_n_14 ),
        .O(\n16[3]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n16[3]_i_8 
       (.I0(\n16_reg[3]_i_17_n_12 ),
        .I1(n22__6_n_0),
        .O(\n16[3]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \n16[3]_i_9 
       (.I0(\n16[3]_i_2_n_0 ),
        .I1(\n16_reg[7]_i_11_n_8 ),
        .I2(\n16_reg[7]_i_10_n_12 ),
        .I3(\n16_reg[7]_i_12_n_5 ),
        .O(\n16[3]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \n16[7]_i_13__1 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_13__1_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \n16[7]_i_14 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(\n16[7]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \n16[7]_i_15__1 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_15__1_n_0 ));
  LUT3 #(
    .INIT(8'h4D)) 
    \n16[7]_i_16__1 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(\n16[7]_i_16__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n16[7]_i_17 
       (.I0(n22_n_0),
        .O(\n16[7]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n16[7]_i_18 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n16[7]_i_19__1 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .O(\n16[7]_i_19__1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n16[7]_i_2 
       (.I0(\n16_reg[7]_i_9_n_14 ),
        .I1(\n16_reg[7]_i_10_n_10 ),
        .O(\n16[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n16[7]_i_20__1 
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .O(\n16[7]_i_20__1_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n16[7]_i_21__1 
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .O(\n16[7]_i_21__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n16[7]_i_22 
       (.I0(n22__5_n_0),
        .O(\n16[7]_i_22_n_0 ));
  (* HLUTNM = "lutpair102" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_23__1 
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .O(\n16[7]_i_23__1_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_24 
       (.I0(n22__3_n_0),
        .I1(n22__2_n_0),
        .I2(n22__1_n_0),
        .O(\n16[7]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_25 
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__2_n_0),
        .O(\n16[7]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_26 
       (.I0(n22__5_n_0),
        .I1(n22__4_n_0),
        .I2(n22__3_n_0),
        .O(\n16[7]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n16[7]_i_27 
       (.I0(n22__4_n_0),
        .I1(n22__5_n_0),
        .I2(n22__3_n_0),
        .O(\n16[7]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h9669)) 
    \n16[7]_i_28 
       (.I0(\n16[7]_i_23__1_n_0 ),
        .I1(n22__0_n_0),
        .I2(n22__1_n_0),
        .I3(n22_n_0),
        .O(\n16[7]_i_28_n_0 ));
  (* HLUTNM = "lutpair102" *) 
  LUT4 #(
    .INIT(16'h781E)) 
    \n16[7]_i_29__1 
       (.I0(n22__2_n_0),
        .I1(n22__1_n_0),
        .I2(n22__0_n_0),
        .I3(n22__3_n_0),
        .O(\n16[7]_i_29__1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n16[7]_i_3 
       (.I0(\n16_reg[7]_i_9_n_15 ),
        .I1(\n16_reg[7]_i_10_n_11 ),
        .O(\n16[7]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[7]_i_30__1 
       (.I0(n22__4_n_0),
        .I1(n22__2_n_0),
        .I2(n22__3_n_0),
        .I3(n22__1_n_0),
        .O(\n16[7]_i_30__1_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n16[7]_i_31__1 
       (.I0(n22__5_n_0),
        .I1(n22__3_n_0),
        .I2(n22__4_n_0),
        .I3(n22__2_n_0),
        .O(\n16[7]_i_31__1_n_0 ));
  LUT4 #(
    .INIT(16'h6696)) 
    \n16[7]_i_32__1 
       (.I0(n22__4_n_0),
        .I1(n22__3_n_0),
        .I2(n22__5_n_0),
        .I3(n22__6_n_0),
        .O(\n16[7]_i_32__1_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n16[7]_i_33 
       (.I0(n22__6_n_0),
        .I1(n22__5_n_0),
        .I2(n22__4_n_0),
        .O(\n16[7]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n16[7]_i_34__1 
       (.I0(n22__5_n_0),
        .I1(n22__6_n_0),
        .O(\n16[7]_i_34__1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \n16[7]_i_35__1 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_35__1_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \n16[7]_i_36 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(\n16[7]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \n16[7]_i_37__1 
       (.I0(n22__0_n_0),
        .I1(n22_n_0),
        .O(\n16[7]_i_37__1_n_0 ));
  LUT3 #(
    .INIT(8'h4D)) 
    \n16[7]_i_38__1 
       (.I0(n22__1_n_0),
        .I1(n22__0_n_0),
        .I2(n22_n_0),
        .O(\n16[7]_i_38__1_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n16[7]_i_4 
       (.I0(\n16_reg[7]_i_10_n_12 ),
        .I1(\n16_reg[7]_i_11_n_8 ),
        .I2(\n16_reg[7]_i_12_n_5 ),
        .O(\n16[7]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \n16[7]_i_5__1 
       (.I0(\n16_reg[7]_i_9_n_5 ),
        .I1(\n16_reg[7]_i_10_n_9 ),
        .I2(\n16_reg[7]_i_10_n_8 ),
        .O(\n16[7]_i_5__1_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n16[7]_i_6__1 
       (.I0(\n16_reg[7]_i_9_n_14 ),
        .I1(\n16_reg[7]_i_10_n_10 ),
        .I2(\n16_reg[7]_i_10_n_9 ),
        .I3(\n16_reg[7]_i_9_n_5 ),
        .O(\n16[7]_i_6__1_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n16[7]_i_7__1 
       (.I0(\n16_reg[7]_i_9_n_15 ),
        .I1(\n16_reg[7]_i_10_n_11 ),
        .I2(\n16_reg[7]_i_10_n_10 ),
        .I3(\n16_reg[7]_i_9_n_14 ),
        .O(\n16[7]_i_7__1_n_0 ));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    \n16[7]_i_8 
       (.I0(\n16_reg[7]_i_12_n_5 ),
        .I1(\n16_reg[7]_i_11_n_8 ),
        .I2(\n16_reg[7]_i_10_n_12 ),
        .I3(\n16_reg[7]_i_10_n_11 ),
        .I4(\n16_reg[7]_i_9_n_15 ),
        .O(\n16[7]_i_8_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[0]),
        .Q(\n16_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[1]),
        .Q(\n16_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[2]),
        .Q(\n16_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[3]),
        .Q(\n16_reg_n_0_[3] ),
        .R(rst_i));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[3]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n16_reg[3]_i_1_n_0 ,\n16_reg[3]_i_1_n_1 ,\n16_reg[3]_i_1_n_2 ,\n16_reg[3]_i_1_n_3 ,\n16_reg[3]_i_1_n_4 ,\n16_reg[3]_i_1_n_5 ,\n16_reg[3]_i_1_n_6 ,\n16_reg[3]_i_1_n_7 }),
        .DI({\n16[3]_i_2_n_0 ,\n16[3]_i_3_n_0 ,\n16[3]_i_4_n_0 ,\n16[3]_i_5_n_0 ,\n16[3]_i_6__1_n_0 ,\n16[3]_i_7_n_0 ,\n16[3]_i_8_n_0 ,1'b0}),
        .O({n15[3:0],\NLW_n16_reg[3]_i_1_O_UNCONNECTED [3:0]}),
        .S({\n16[3]_i_9_n_0 ,\n16[3]_i_10_n_0 ,\n16[3]_i_11_n_0 ,\n16[3]_i_12_n_0 ,\n16[3]_i_13_n_0 ,\n16[3]_i_14__1_n_0 ,\n16[3]_i_15__1_n_0 ,\n16[3]_i_16_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[3]_i_17 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n16_reg[3]_i_17_n_0 ,\n16_reg[3]_i_17_n_1 ,\n16_reg[3]_i_17_n_2 ,\n16_reg[3]_i_17_n_3 ,\n16_reg[3]_i_17_n_4 ,\n16_reg[3]_i_17_n_5 ,\n16_reg[3]_i_17_n_6 ,\n16_reg[3]_i_17_n_7 }),
        .DI({\n16[7]_i_23__1_n_0 ,\n16[3]_i_18_n_0 ,\n16[3]_i_19_n_0 ,\n16[3]_i_20_n_0 ,\n16[3]_i_21_n_0 ,n22__4_n_0,n22__5_n_0,1'b0}),
        .O({\n16_reg[3]_i_17_n_8 ,\n16_reg[3]_i_17_n_9 ,\n16_reg[3]_i_17_n_10 ,\n16_reg[3]_i_17_n_11 ,\n16_reg[3]_i_17_n_12 ,\NLW_n16_reg[3]_i_17_O_UNCONNECTED [2:1],\n16_reg[3]_i_17_n_15 }),
        .S({\n16[3]_i_22_n_0 ,\n16[3]_i_23__1_n_0 ,\n16[3]_i_24__1_n_0 ,\n16[3]_i_25__1_n_0 ,\n16[3]_i_26__1_n_0 ,\n16[3]_i_27_n_0 ,\n16[3]_i_28__1_n_0 ,n22__6_n_0}));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[4]),
        .Q(\n16_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[5]),
        .Q(\n16_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[6]),
        .Q(\n16_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n16_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n15[7]),
        .Q(\n16_reg_n_0_[7] ),
        .R(rst_i));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_1 
       (.CI(\n16_reg[3]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n16_reg[7]_i_1_CO_UNCONNECTED [7:3],\n16_reg[7]_i_1_n_5 ,\n16_reg[7]_i_1_n_6 ,\n16_reg[7]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,\n16[7]_i_2_n_0 ,\n16[7]_i_3_n_0 ,\n16[7]_i_4_n_0 }),
        .O({\NLW_n16_reg[7]_i_1_O_UNCONNECTED [7:4],n15[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,\n16[7]_i_5__1_n_0 ,\n16[7]_i_6__1_n_0 ,\n16[7]_i_7__1_n_0 ,\n16[7]_i_8_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_10 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\NLW_n16_reg[7]_i_10_CO_UNCONNECTED [7],\n16_reg[7]_i_10_n_1 ,\n16_reg[7]_i_10_n_2 ,\n16_reg[7]_i_10_n_3 ,\n16_reg[7]_i_10_n_4 ,\n16_reg[7]_i_10_n_5 ,\n16_reg[7]_i_10_n_6 ,\n16_reg[7]_i_10_n_7 }),
        .DI({1'b0,n22__0_n_0,n22__1_n_0,n22__2_n_0,n22__3_n_0,1'b1,1'b0,1'b1}),
        .O({\n16_reg[7]_i_10_n_8 ,\n16_reg[7]_i_10_n_9 ,\n16_reg[7]_i_10_n_10 ,\n16_reg[7]_i_10_n_11 ,\n16_reg[7]_i_10_n_12 ,\n16_reg[7]_i_10_n_13 ,\n16_reg[7]_i_10_n_14 ,\n16_reg[7]_i_10_n_15 }),
        .S({\n16[7]_i_17_n_0 ,\n16[7]_i_18_n_0 ,\n16[7]_i_19__1_n_0 ,\n16[7]_i_20__1_n_0 ,\n16[7]_i_21__1_n_0 ,n22__3_n_0,n22__4_n_0,\n16[7]_i_22_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_11 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n16_reg[7]_i_11_n_0 ,\n16_reg[7]_i_11_n_1 ,\n16_reg[7]_i_11_n_2 ,\n16_reg[7]_i_11_n_3 ,\n16_reg[7]_i_11_n_4 ,\n16_reg[7]_i_11_n_5 ,\n16_reg[7]_i_11_n_6 ,\n16_reg[7]_i_11_n_7 }),
        .DI({\n16[7]_i_23__1_n_0 ,\n16[7]_i_24_n_0 ,\n16[7]_i_25_n_0 ,\n16[7]_i_26_n_0 ,\n16[7]_i_27_n_0 ,n22__4_n_0,n22__5_n_0,1'b0}),
        .O({\n16_reg[7]_i_11_n_8 ,\n16_reg[7]_i_11_n_9 ,\n16_reg[7]_i_11_n_10 ,\n16_reg[7]_i_11_n_11 ,\n16_reg[7]_i_11_n_12 ,\n16_reg[7]_i_11_n_13 ,\n16_reg[7]_i_11_n_14 ,\NLW_n16_reg[7]_i_11_O_UNCONNECTED [0]}),
        .S({\n16[7]_i_28_n_0 ,\n16[7]_i_29__1_n_0 ,\n16[7]_i_30__1_n_0 ,\n16[7]_i_31__1_n_0 ,\n16[7]_i_32__1_n_0 ,\n16[7]_i_33_n_0 ,\n16[7]_i_34__1_n_0 ,n22__6_n_0}));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_12 
       (.CI(\n16_reg[3]_i_17_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n16_reg[7]_i_12_CO_UNCONNECTED [7:3],\n16_reg[7]_i_12_n_5 ,\NLW_n16_reg[7]_i_12_CO_UNCONNECTED [1],\n16_reg[7]_i_12_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\n16[7]_i_35__1_n_0 ,\n16[7]_i_36_n_0 }),
        .O({\NLW_n16_reg[7]_i_12_O_UNCONNECTED [7:2],\n16_reg[7]_i_12_n_14 ,\n16_reg[7]_i_12_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,\n16[7]_i_37__1_n_0 ,\n16[7]_i_38__1_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n16_reg[7]_i_9 
       (.CI(\n16_reg[7]_i_11_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n16_reg[7]_i_9_CO_UNCONNECTED [7:3],\n16_reg[7]_i_9_n_5 ,\NLW_n16_reg[7]_i_9_CO_UNCONNECTED [1],\n16_reg[7]_i_9_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\n16[7]_i_13__1_n_0 ,\n16[7]_i_14_n_0 }),
        .O({\NLW_n16_reg[7]_i_9_O_UNCONNECTED [7:2],\n16_reg[7]_i_9_n_14 ,\n16_reg[7]_i_9_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,\n16[7]_i_15__1_n_0 ,\n16[7]_i_16__1_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[0]),
        .Q(\n1_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[10]),
        .Q(n2[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[11]),
        .Q(n2[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[12]),
        .Q(n2[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[13]),
        .Q(n2[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[14]),
        .Q(n2[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[15]),
        .Q(n2[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[1]),
        .Q(\n1_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[2]),
        .Q(\n1_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[3]),
        .Q(\n1_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[4]),
        .Q(\n1_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[5]),
        .Q(\n1_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[6]),
        .Q(\n1_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[7]),
        .Q(\n1_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[8]),
        .Q(n2[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n1_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(D[9]),
        .Q(n2[1]),
        .R(rst_i));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_2__1 
       (.I0(\n16_reg_n_0_[7] ),
        .O(\n21[7]_i_2__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_3__1 
       (.I0(\n16_reg_n_0_[6] ),
        .O(\n21[7]_i_3__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_4__1 
       (.I0(\n16_reg_n_0_[5] ),
        .O(\n21[7]_i_4__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_5__1 
       (.I0(\n16_reg_n_0_[4] ),
        .O(\n21[7]_i_5__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_6__1 
       (.I0(\n16_reg_n_0_[3] ),
        .O(\n21[7]_i_6__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_7__1 
       (.I0(\n16_reg_n_0_[2] ),
        .O(\n21[7]_i_7__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_8__1 
       (.I0(\n16_reg_n_0_[1] ),
        .O(\n21[7]_i_8__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n21[7]_i_9__1 
       (.I0(\n16_reg_n_0_[0] ),
        .O(\n21[7]_i_9__1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[0]),
        .Q(n21[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[1]),
        .Q(n21[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[2]),
        .Q(n21[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[3]),
        .Q(n21[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[4]),
        .Q(n21[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[5]),
        .Q(n21[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[6]),
        .Q(n21[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n21_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n202_out[7]),
        .Q(n21[7]),
        .R(rst_i));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n21_reg[7]_i_1__1 
       (.CI(1'b1),
        .CI_TOP(1'b0),
        .CO({\NLW_n21_reg[7]_i_1__1_CO_UNCONNECTED [7],\n21_reg[7]_i_1__1_n_1 ,\n21_reg[7]_i_1__1_n_2 ,\n21_reg[7]_i_1__1_n_3 ,\n21_reg[7]_i_1__1_n_4 ,\n21_reg[7]_i_1__1_n_5 ,\n21_reg[7]_i_1__1_n_6 ,\n21_reg[7]_i_1__1_n_7 }),
        .DI({1'b0,\n16_reg_n_0_[6] ,\n16_reg_n_0_[5] ,\n16_reg_n_0_[4] ,\n16_reg_n_0_[3] ,\n16_reg_n_0_[2] ,\n16_reg_n_0_[1] ,\n16_reg_n_0_[0] }),
        .O(n202_out),
        .S({\n21[7]_i_2__1_n_0 ,\n21[7]_i_3__1_n_0 ,\n21[7]_i_4__1_n_0 ,\n21[7]_i_5__1_n_0 ,\n21[7]_i_6__1_n_0 ,\n21[7]_i_7__1_n_0 ,\n21[7]_i_8__1_n_0 ,\n21[7]_i_9__1_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    n22
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[15]),
        .Q(n22_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__0
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[14]),
        .Q(n22__0_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__1
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[13]),
        .Q(n22__1_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__2
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[12]),
        .Q(n22__2_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__3
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[11]),
        .Q(n22__3_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__4
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[10]),
        .Q(n22__4_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__5
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[9]),
        .Q(n22__5_n_0),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    n22__6
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[8]),
        .Q(n22__6_n_0),
        .R(rst_i));
  (* HLUTNM = "lutpair59" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_10 
       (.I0(\n27_reg[7]_i_10_n_13 ),
        .I1(\n27_reg[7]_i_11_n_9 ),
        .I2(\n27_reg[7]_i_12_n_14 ),
        .I3(\n27[3]_i_3_n_0 ),
        .O(\n27[3]_i_10_n_0 ));
  (* HLUTNM = "lutpair58" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_11 
       (.I0(\n27_reg[7]_i_10_n_14 ),
        .I1(\n27_reg[7]_i_11_n_10 ),
        .I2(\n27_reg[7]_i_12_n_15 ),
        .I3(\n27[3]_i_4_n_0 ),
        .O(\n27[3]_i_11_n_0 ));
  (* HLUTNM = "lutpair57" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_12 
       (.I0(\n27_reg[7]_i_10_n_15 ),
        .I1(\n27_reg[7]_i_11_n_11 ),
        .I2(\n27_reg[3]_i_17_n_8 ),
        .I3(\n27[3]_i_5_n_0 ),
        .O(\n27[3]_i_12_n_0 ));
  (* HLUTNM = "lutpair56" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_13 
       (.I0(\n27_reg[3]_i_17_n_15 ),
        .I1(\n27_reg[7]_i_11_n_12 ),
        .I2(\n27_reg[3]_i_17_n_9 ),
        .I3(\n27[3]_i_6__1_n_0 ),
        .O(\n27[3]_i_13_n_0 ));
  (* HLUTNM = "lutpair101" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n27[3]_i_14__1 
       (.I0(\n27_reg[7]_i_11_n_13 ),
        .I1(\n27_reg[3]_i_17_n_10 ),
        .I2(\n27_reg[3]_i_17_n_11 ),
        .I3(\n27_reg[7]_i_11_n_14 ),
        .O(\n27[3]_i_14__1_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n27[3]_i_15__1 
       (.I0(\n27_reg[3]_i_17_n_12 ),
        .I1(\n4_reg_n_0_[0] ),
        .I2(\n27_reg[7]_i_11_n_14 ),
        .I3(\n27_reg[3]_i_17_n_11 ),
        .O(\n27[3]_i_15__1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n27[3]_i_16 
       (.I0(\n27_reg[3]_i_17_n_12 ),
        .I1(\n4_reg_n_0_[0] ),
        .O(\n27[3]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_18 
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[5] ),
        .O(\n27[3]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_19 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[4] ),
        .O(\n27[3]_i_19_n_0 ));
  (* HLUTNM = "lutpair59" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_2 
       (.I0(\n27_reg[7]_i_10_n_13 ),
        .I1(\n27_reg[7]_i_11_n_9 ),
        .I2(\n27_reg[7]_i_12_n_14 ),
        .O(\n27[3]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_20 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[2] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(\n27[3]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n27[3]_i_21 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(\n27[3]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h9669)) 
    \n27[3]_i_22 
       (.I0(\n27[7]_i_23__1_n_0 ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[5] ),
        .I3(\n4_reg_n_0_[7] ),
        .O(\n27[3]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[3]_i_23__1 
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[5] ),
        .I2(\n4_reg_n_0_[4] ),
        .I3(\n4_reg_n_0_[6] ),
        .O(\n27[3]_i_23__1_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[3]_i_24__1 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[3] ),
        .I3(\n4_reg_n_0_[5] ),
        .O(\n27[3]_i_24__1_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[3]_i_25__1 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[2] ),
        .I3(\n4_reg_n_0_[4] ),
        .O(\n27[3]_i_25__1_n_0 ));
  LUT4 #(
    .INIT(16'h6696)) 
    \n27[3]_i_26__1 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[1] ),
        .I3(\n4_reg_n_0_[0] ),
        .O(\n27[3]_i_26__1_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n27[3]_i_27 
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[2] ),
        .O(\n27[3]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n27[3]_i_28__1 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[0] ),
        .O(\n27[3]_i_28__1_n_0 ));
  (* HLUTNM = "lutpair58" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_3 
       (.I0(\n27_reg[7]_i_10_n_14 ),
        .I1(\n27_reg[7]_i_11_n_10 ),
        .I2(\n27_reg[7]_i_12_n_15 ),
        .O(\n27[3]_i_3_n_0 ));
  (* HLUTNM = "lutpair57" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_4 
       (.I0(\n27_reg[7]_i_10_n_15 ),
        .I1(\n27_reg[7]_i_11_n_11 ),
        .I2(\n27_reg[3]_i_17_n_8 ),
        .O(\n27[3]_i_4_n_0 ));
  (* HLUTNM = "lutpair56" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[3]_i_5 
       (.I0(\n27_reg[3]_i_17_n_15 ),
        .I1(\n27_reg[7]_i_11_n_12 ),
        .I2(\n27_reg[3]_i_17_n_9 ),
        .O(\n27[3]_i_5_n_0 ));
  (* HLUTNM = "lutpair101" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \n27[3]_i_6__1 
       (.I0(\n27_reg[7]_i_11_n_13 ),
        .I1(\n27_reg[3]_i_17_n_10 ),
        .O(\n27[3]_i_6__1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n27[3]_i_7 
       (.I0(\n27_reg[3]_i_17_n_11 ),
        .I1(\n27_reg[7]_i_11_n_14 ),
        .O(\n27[3]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n27[3]_i_8 
       (.I0(\n27_reg[3]_i_17_n_12 ),
        .I1(\n4_reg_n_0_[0] ),
        .O(\n27[3]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \n27[3]_i_9 
       (.I0(\n27[3]_i_2_n_0 ),
        .I1(\n27_reg[7]_i_11_n_8 ),
        .I2(\n27_reg[7]_i_10_n_12 ),
        .I3(\n27_reg[7]_i_12_n_5 ),
        .O(\n27[3]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \n27[7]_i_13__1 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_13__1_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \n27[7]_i_14 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \n27[7]_i_15__1 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_15__1_n_0 ));
  LUT3 #(
    .INIT(8'h4D)) 
    \n27[7]_i_16__1 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_16__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n27[7]_i_17 
       (.I0(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n27[7]_i_18 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n27[7]_i_19__1 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .O(\n27[7]_i_19__1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n27[7]_i_2 
       (.I0(\n27_reg[7]_i_9_n_14 ),
        .I1(\n27_reg[7]_i_10_n_10 ),
        .O(\n27[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n27[7]_i_20__1 
       (.I0(\n4_reg_n_0_[4] ),
        .I1(\n4_reg_n_0_[5] ),
        .O(\n27[7]_i_20__1_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \n27[7]_i_21__1 
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[4] ),
        .O(\n27[7]_i_21__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \n27[7]_i_22 
       (.I0(\n4_reg_n_0_[1] ),
        .O(\n27[7]_i_22_n_0 ));
  (* HLUTNM = "lutpair100" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_23__1 
       (.I0(\n4_reg_n_0_[4] ),
        .I1(\n4_reg_n_0_[5] ),
        .I2(\n4_reg_n_0_[6] ),
        .O(\n27[7]_i_23__1_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_24 
       (.I0(\n4_reg_n_0_[3] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[5] ),
        .O(\n27[7]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_25 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[4] ),
        .O(\n27[7]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_26 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[2] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(\n27[7]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n27[7]_i_27 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[3] ),
        .O(\n27[7]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h9669)) 
    \n27[7]_i_28 
       (.I0(\n27[7]_i_23__1_n_0 ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[5] ),
        .I3(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_28_n_0 ));
  (* HLUTNM = "lutpair100" *) 
  LUT4 #(
    .INIT(16'h781E)) 
    \n27[7]_i_29__1 
       (.I0(\n4_reg_n_0_[4] ),
        .I1(\n4_reg_n_0_[5] ),
        .I2(\n4_reg_n_0_[6] ),
        .I3(\n4_reg_n_0_[3] ),
        .O(\n27[7]_i_29__1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \n27[7]_i_3 
       (.I0(\n27_reg[7]_i_9_n_15 ),
        .I1(\n27_reg[7]_i_10_n_11 ),
        .O(\n27[7]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[7]_i_30__1 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[4] ),
        .I2(\n4_reg_n_0_[3] ),
        .I3(\n4_reg_n_0_[5] ),
        .O(\n27[7]_i_30__1_n_0 ));
  LUT4 #(
    .INIT(16'h2BD4)) 
    \n27[7]_i_31__1 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[2] ),
        .I3(\n4_reg_n_0_[4] ),
        .O(\n27[7]_i_31__1_n_0 ));
  LUT4 #(
    .INIT(16'h6696)) 
    \n27[7]_i_32__1 
       (.I0(\n4_reg_n_0_[2] ),
        .I1(\n4_reg_n_0_[3] ),
        .I2(\n4_reg_n_0_[1] ),
        .I3(\n4_reg_n_0_[0] ),
        .O(\n27[7]_i_32__1_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \n27[7]_i_33 
       (.I0(\n4_reg_n_0_[0] ),
        .I1(\n4_reg_n_0_[1] ),
        .I2(\n4_reg_n_0_[2] ),
        .O(\n27[7]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n27[7]_i_34__1 
       (.I0(\n4_reg_n_0_[1] ),
        .I1(\n4_reg_n_0_[0] ),
        .O(\n27[7]_i_34__1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \n27[7]_i_35__1 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_35__1_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \n27[7]_i_36 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \n27[7]_i_37__1 
       (.I0(\n4_reg_n_0_[6] ),
        .I1(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_37__1_n_0 ));
  LUT3 #(
    .INIT(8'h4D)) 
    \n27[7]_i_38__1 
       (.I0(\n4_reg_n_0_[5] ),
        .I1(\n4_reg_n_0_[6] ),
        .I2(\n4_reg_n_0_[7] ),
        .O(\n27[7]_i_38__1_n_0 ));
  LUT3 #(
    .INIT(8'hE8)) 
    \n27[7]_i_4 
       (.I0(\n27_reg[7]_i_10_n_12 ),
        .I1(\n27_reg[7]_i_11_n_8 ),
        .I2(\n27_reg[7]_i_12_n_5 ),
        .O(\n27[7]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \n27[7]_i_5__1 
       (.I0(\n27_reg[7]_i_9_n_5 ),
        .I1(\n27_reg[7]_i_10_n_9 ),
        .I2(\n27_reg[7]_i_10_n_8 ),
        .O(\n27[7]_i_5__1_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n27[7]_i_6__1 
       (.I0(\n27_reg[7]_i_9_n_14 ),
        .I1(\n27_reg[7]_i_10_n_10 ),
        .I2(\n27_reg[7]_i_10_n_9 ),
        .I3(\n27_reg[7]_i_9_n_5 ),
        .O(\n27[7]_i_6__1_n_0 ));
  LUT4 #(
    .INIT(16'h8778)) 
    \n27[7]_i_7__1 
       (.I0(\n27_reg[7]_i_9_n_15 ),
        .I1(\n27_reg[7]_i_10_n_11 ),
        .I2(\n27_reg[7]_i_10_n_10 ),
        .I3(\n27_reg[7]_i_9_n_14 ),
        .O(\n27[7]_i_7__1_n_0 ));
  LUT5 #(
    .INIT(32'hE81717E8)) 
    \n27[7]_i_8 
       (.I0(\n27_reg[7]_i_12_n_5 ),
        .I1(\n27_reg[7]_i_11_n_8 ),
        .I2(\n27_reg[7]_i_10_n_12 ),
        .I3(\n27_reg[7]_i_10_n_11 ),
        .I4(\n27_reg[7]_i_9_n_15 ),
        .O(\n27[7]_i_8_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[0]),
        .Q(n27[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[1]),
        .Q(n27[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[2]),
        .Q(n27[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[3]),
        .Q(n27[3]),
        .R(rst_i));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[3]_i_1 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n27_reg[3]_i_1_n_0 ,\n27_reg[3]_i_1_n_1 ,\n27_reg[3]_i_1_n_2 ,\n27_reg[3]_i_1_n_3 ,\n27_reg[3]_i_1_n_4 ,\n27_reg[3]_i_1_n_5 ,\n27_reg[3]_i_1_n_6 ,\n27_reg[3]_i_1_n_7 }),
        .DI({\n27[3]_i_2_n_0 ,\n27[3]_i_3_n_0 ,\n27[3]_i_4_n_0 ,\n27[3]_i_5_n_0 ,\n27[3]_i_6__1_n_0 ,\n27[3]_i_7_n_0 ,\n27[3]_i_8_n_0 ,1'b0}),
        .O({n26[3:0],\NLW_n27_reg[3]_i_1_O_UNCONNECTED [3:0]}),
        .S({\n27[3]_i_9_n_0 ,\n27[3]_i_10_n_0 ,\n27[3]_i_11_n_0 ,\n27[3]_i_12_n_0 ,\n27[3]_i_13_n_0 ,\n27[3]_i_14__1_n_0 ,\n27[3]_i_15__1_n_0 ,\n27[3]_i_16_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[3]_i_17 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n27_reg[3]_i_17_n_0 ,\n27_reg[3]_i_17_n_1 ,\n27_reg[3]_i_17_n_2 ,\n27_reg[3]_i_17_n_3 ,\n27_reg[3]_i_17_n_4 ,\n27_reg[3]_i_17_n_5 ,\n27_reg[3]_i_17_n_6 ,\n27_reg[3]_i_17_n_7 }),
        .DI({\n27[7]_i_23__1_n_0 ,\n27[3]_i_18_n_0 ,\n27[3]_i_19_n_0 ,\n27[3]_i_20_n_0 ,\n27[3]_i_21_n_0 ,\n4_reg_n_0_[2] ,\n4_reg_n_0_[1] ,1'b0}),
        .O({\n27_reg[3]_i_17_n_8 ,\n27_reg[3]_i_17_n_9 ,\n27_reg[3]_i_17_n_10 ,\n27_reg[3]_i_17_n_11 ,\n27_reg[3]_i_17_n_12 ,\NLW_n27_reg[3]_i_17_O_UNCONNECTED [2:1],\n27_reg[3]_i_17_n_15 }),
        .S({\n27[3]_i_22_n_0 ,\n27[3]_i_23__1_n_0 ,\n27[3]_i_24__1_n_0 ,\n27[3]_i_25__1_n_0 ,\n27[3]_i_26__1_n_0 ,\n27[3]_i_27_n_0 ,\n27[3]_i_28__1_n_0 ,\n4_reg_n_0_[0] }));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[4]),
        .Q(n27[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[5]),
        .Q(n27[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[6]),
        .Q(n27[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n27_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n26[7]),
        .Q(n27[7]),
        .R(rst_i));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_1 
       (.CI(\n27_reg[3]_i_1_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n27_reg[7]_i_1_CO_UNCONNECTED [7:3],\n27_reg[7]_i_1_n_5 ,\n27_reg[7]_i_1_n_6 ,\n27_reg[7]_i_1_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,\n27[7]_i_2_n_0 ,\n27[7]_i_3_n_0 ,\n27[7]_i_4_n_0 }),
        .O({\NLW_n27_reg[7]_i_1_O_UNCONNECTED [7:4],n26[7:4]}),
        .S({1'b0,1'b0,1'b0,1'b0,\n27[7]_i_5__1_n_0 ,\n27[7]_i_6__1_n_0 ,\n27[7]_i_7__1_n_0 ,\n27[7]_i_8_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_10 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\NLW_n27_reg[7]_i_10_CO_UNCONNECTED [7],\n27_reg[7]_i_10_n_1 ,\n27_reg[7]_i_10_n_2 ,\n27_reg[7]_i_10_n_3 ,\n27_reg[7]_i_10_n_4 ,\n27_reg[7]_i_10_n_5 ,\n27_reg[7]_i_10_n_6 ,\n27_reg[7]_i_10_n_7 }),
        .DI({1'b0,\n4_reg_n_0_[6] ,\n4_reg_n_0_[5] ,\n4_reg_n_0_[4] ,\n4_reg_n_0_[3] ,1'b1,1'b0,1'b1}),
        .O({\n27_reg[7]_i_10_n_8 ,\n27_reg[7]_i_10_n_9 ,\n27_reg[7]_i_10_n_10 ,\n27_reg[7]_i_10_n_11 ,\n27_reg[7]_i_10_n_12 ,\n27_reg[7]_i_10_n_13 ,\n27_reg[7]_i_10_n_14 ,\n27_reg[7]_i_10_n_15 }),
        .S({\n27[7]_i_17_n_0 ,\n27[7]_i_18_n_0 ,\n27[7]_i_19__1_n_0 ,\n27[7]_i_20__1_n_0 ,\n27[7]_i_21__1_n_0 ,\n4_reg_n_0_[3] ,\n4_reg_n_0_[2] ,\n27[7]_i_22_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_11 
       (.CI(1'b0),
        .CI_TOP(1'b0),
        .CO({\n27_reg[7]_i_11_n_0 ,\n27_reg[7]_i_11_n_1 ,\n27_reg[7]_i_11_n_2 ,\n27_reg[7]_i_11_n_3 ,\n27_reg[7]_i_11_n_4 ,\n27_reg[7]_i_11_n_5 ,\n27_reg[7]_i_11_n_6 ,\n27_reg[7]_i_11_n_7 }),
        .DI({\n27[7]_i_23__1_n_0 ,\n27[7]_i_24_n_0 ,\n27[7]_i_25_n_0 ,\n27[7]_i_26_n_0 ,\n27[7]_i_27_n_0 ,\n4_reg_n_0_[2] ,\n4_reg_n_0_[1] ,1'b0}),
        .O({\n27_reg[7]_i_11_n_8 ,\n27_reg[7]_i_11_n_9 ,\n27_reg[7]_i_11_n_10 ,\n27_reg[7]_i_11_n_11 ,\n27_reg[7]_i_11_n_12 ,\n27_reg[7]_i_11_n_13 ,\n27_reg[7]_i_11_n_14 ,\NLW_n27_reg[7]_i_11_O_UNCONNECTED [0]}),
        .S({\n27[7]_i_28_n_0 ,\n27[7]_i_29__1_n_0 ,\n27[7]_i_30__1_n_0 ,\n27[7]_i_31__1_n_0 ,\n27[7]_i_32__1_n_0 ,\n27[7]_i_33_n_0 ,\n27[7]_i_34__1_n_0 ,\n4_reg_n_0_[0] }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_12 
       (.CI(\n27_reg[3]_i_17_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n27_reg[7]_i_12_CO_UNCONNECTED [7:3],\n27_reg[7]_i_12_n_5 ,\NLW_n27_reg[7]_i_12_CO_UNCONNECTED [1],\n27_reg[7]_i_12_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\n27[7]_i_35__1_n_0 ,\n27[7]_i_36_n_0 }),
        .O({\NLW_n27_reg[7]_i_12_O_UNCONNECTED [7:2],\n27_reg[7]_i_12_n_14 ,\n27_reg[7]_i_12_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,\n27[7]_i_37__1_n_0 ,\n27[7]_i_38__1_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-9 {cell *THIS*} {string 8x8}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \n27_reg[7]_i_9 
       (.CI(\n27_reg[7]_i_11_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_n27_reg[7]_i_9_CO_UNCONNECTED [7:3],\n27_reg[7]_i_9_n_5 ,\NLW_n27_reg[7]_i_9_CO_UNCONNECTED [1],\n27_reg[7]_i_9_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\n27[7]_i_13__1_n_0 ,\n27[7]_i_14_n_0 }),
        .O({\NLW_n27_reg[7]_i_9_O_UNCONNECTED [7:2],\n27_reg[7]_i_9_n_14 ,\n27_reg[7]_i_9_n_15 }),
        .S({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,\n27[7]_i_15__1_n_0 ,\n27[7]_i_16__1_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[0]),
        .Q(n29[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[1]),
        .Q(n29[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[2]),
        .Q(n29[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[3]),
        .Q(n29[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[4]),
        .Q(n29[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[5]),
        .Q(n29[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[6]),
        .Q(n29[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n29_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n27[7]),
        .Q(n29[7]),
        .R(rst_i));
  LUT2 #(
    .INIT(4'h6)) 
    \n33[0]_i_1__5 
       (.I0(n29[0]),
        .I1(n10[0]),
        .O(n31[0]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[10]_i_1__5 
       (.I0(n21[2]),
        .I1(\n8_reg_n_0_[2] ),
        .I2(\n8_reg_n_0_[1] ),
        .I3(n21[1]),
        .I4(\n8_reg_n_0_[0] ),
        .I5(n21[0]),
        .O(\n33[10]_i_1__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[11]_i_1__5 
       (.I0(n21[3]),
        .I1(\n8_reg_n_0_[3] ),
        .I2(\n33[12]_i_2__5_n_0 ),
        .O(\n33[11]_i_1__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[12]_i_1__5 
       (.I0(n21[4]),
        .I1(\n8_reg_n_0_[4] ),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[3]),
        .I4(\n33[12]_i_2__5_n_0 ),
        .O(\n33[12]_i_1__5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[12]_i_2__5 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n33[12]_i_2__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[13]_i_1__5 
       (.I0(n21[5]),
        .I1(\n8_reg_n_0_[5] ),
        .I2(\n33[14]_i_2__5_n_0 ),
        .O(\n33[13]_i_1__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[14]_i_1__5 
       (.I0(n21[6]),
        .I1(\n8_reg_n_0_[6] ),
        .I2(\n8_reg_n_0_[5] ),
        .I3(n21[5]),
        .I4(\n33[14]_i_2__5_n_0 ),
        .O(\n33[14]_i_1__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[14]_i_2__5 
       (.I0(\n33[12]_i_2__5_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n33[14]_i_2__5_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[15]_i_1__5 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n33[15]_i_2__5_n_0 ),
        .O(n30));
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[15]_i_2__5 
       (.I0(\n33[14]_i_2__5_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n33[15]_i_2__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[1]_i_1__5 
       (.I0(n29[1]),
        .I1(n10[1]),
        .I2(n10[0]),
        .I3(n29[0]),
        .O(n31[1]));
  LUT6 #(
    .INIT(64'h9996966696669666)) 
    \n33[2]_i_1__5 
       (.I0(n29[2]),
        .I1(n10[2]),
        .I2(n10[1]),
        .I3(n29[1]),
        .I4(n10[0]),
        .I5(n29[0]),
        .O(\n33[2]_i_1__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[3]_i_1__5 
       (.I0(n29[3]),
        .I1(n10[3]),
        .I2(\n33[4]_i_2__5_n_0 ),
        .O(\n33[3]_i_1__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[4]_i_1__5 
       (.I0(n29[4]),
        .I1(n10[4]),
        .I2(n10[3]),
        .I3(n29[3]),
        .I4(\n33[4]_i_2__5_n_0 ),
        .O(\n33[4]_i_1__5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF880F8800000)) 
    \n33[4]_i_2__5 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n33[4]_i_2__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \n33[5]_i_1__5 
       (.I0(n29[5]),
        .I1(n10[5]),
        .I2(\n33[6]_i_2__5_n_0 ),
        .O(\n33[5]_i_1__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[6]_i_1__5 
       (.I0(n29[6]),
        .I1(n10[6]),
        .I2(n10[5]),
        .I3(n29[5]),
        .I4(\n33[6]_i_2__5_n_0 ),
        .O(\n33[6]_i_1__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT5 #(
    .INIT(32'hFFE8E800)) 
    \n33[6]_i_2__5 
       (.I0(\n33[4]_i_2__5_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n33[6]_i_2__5_n_0 ));
  LUT5 #(
    .INIT(32'h99969666)) 
    \n33[7]_i_1__5 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n33[7]_i_2__5_n_0 ),
        .O(n31[7]));
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    \n33[7]_i_2__5 
       (.I0(\n33[6]_i_2__5_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n33[7]_i_2__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT4 #(
    .INIT(16'h9666)) 
    \n33[9]_i_1__5 
       (.I0(n21[1]),
        .I1(\n8_reg_n_0_[1] ),
        .I2(\n8_reg_n_0_[0] ),
        .I3(n21[0]),
        .O(\n33[9]_i_1__5_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[0]),
        .Q(i1[15]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[10]_i_1__5_n_0 ),
        .Q(i1[24]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[11]_i_1__5_n_0 ),
        .Q(i1[25]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[12]_i_1__5_n_0 ),
        .Q(i1[26]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[13]_i_1__5_n_0 ),
        .Q(i1[27]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[14]_i_1__5_n_0 ),
        .Q(i1[28]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n30),
        .Q(i1[29]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[1]),
        .Q(i1[16]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[2]_i_1__5_n_0 ),
        .Q(i1[17]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[3]_i_1__5_n_0 ),
        .Q(i1[18]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[4]_i_1__5_n_0 ),
        .Q(i1[19]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[5]_i_1__5_n_0 ),
        .Q(i1[20]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[6]_i_1__5_n_0 ),
        .Q(i1[21]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n31[7]),
        .Q(i1[22]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n33_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n33[9]_i_1__5_n_0 ),
        .Q(i1[23]),
        .R(rst_i));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[10]_i_1__5 
       (.I0(\n8_reg_n_0_[1] ),
        .I1(n21[1]),
        .I2(n21[0]),
        .I3(\n8_reg_n_0_[0] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(n341_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[11]_i_1__5 
       (.I0(\n37[12]_i_2__5_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .O(n341_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[12]_i_1__5 
       (.I0(\n8_reg_n_0_[3] ),
        .I1(n21[3]),
        .I2(\n37[12]_i_2__5_n_0 ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(n341_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[12]_i_2__5 
       (.I0(\n8_reg_n_0_[0] ),
        .I1(n21[0]),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .I4(n21[2]),
        .I5(\n8_reg_n_0_[2] ),
        .O(\n37[12]_i_2__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[13]_i_1__5 
       (.I0(\n37[14]_i_2__5_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(n341_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[14]_i_1__5 
       (.I0(\n8_reg_n_0_[5] ),
        .I1(n21[5]),
        .I2(\n37[14]_i_2__5_n_0 ),
        .I3(n21[6]),
        .I4(\n8_reg_n_0_[6] ),
        .O(n341_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[14]_i_2__5 
       (.I0(\n37[12]_i_2__5_n_0 ),
        .I1(n21[3]),
        .I2(\n8_reg_n_0_[3] ),
        .I3(n21[4]),
        .I4(\n8_reg_n_0_[4] ),
        .O(\n37[14]_i_2__5_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[15]_i_1__5 
       (.I0(\n8_reg_n_0_[7] ),
        .I1(n21[7]),
        .I2(\n8_reg_n_0_[6] ),
        .I3(n21[6]),
        .I4(\n37[15]_i_2__5_n_0 ),
        .O(n341_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[15]_i_2__5 
       (.I0(\n37[14]_i_2__5_n_0 ),
        .I1(n21[5]),
        .I2(\n8_reg_n_0_[5] ),
        .O(\n37[15]_i_2__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[1]_i_1__5 
       (.I0(n29[0]),
        .I1(n10[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .O(n350_out[1]));
  LUT6 #(
    .INIT(64'h44D4BB2BBB2B44D4)) 
    \n37[2]_i_1__5 
       (.I0(n10[1]),
        .I1(n29[1]),
        .I2(n29[0]),
        .I3(n10[0]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(n350_out[2]));
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[3]_i_1__5 
       (.I0(\n37[4]_i_2__5_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .O(n350_out[3]));
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[4]_i_1__5 
       (.I0(n10[3]),
        .I1(n29[3]),
        .I2(\n37[4]_i_2__5_n_0 ),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(n350_out[4]));
  LUT6 #(
    .INIT(64'hBF0BFFFF0000BF0B)) 
    \n37[4]_i_2__5 
       (.I0(n10[0]),
        .I1(n29[0]),
        .I2(n29[1]),
        .I3(n10[1]),
        .I4(n29[2]),
        .I5(n10[2]),
        .O(\n37[4]_i_2__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \n37[5]_i_1__5 
       (.I0(\n37[6]_i_2__5_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(n350_out[5]));
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT5 #(
    .INIT(32'h4DB2B24D)) 
    \n37[6]_i_1__5 
       (.I0(n10[5]),
        .I1(n29[5]),
        .I2(\n37[6]_i_2__5_n_0 ),
        .I3(n29[6]),
        .I4(n10[6]),
        .O(n350_out[6]));
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT5 #(
    .INIT(32'hB2FF00B2)) 
    \n37[6]_i_2__5 
       (.I0(\n37[4]_i_2__5_n_0 ),
        .I1(n29[3]),
        .I2(n10[3]),
        .I3(n29[4]),
        .I4(n10[4]),
        .O(\n37[6]_i_2__5_n_0 ));
  LUT5 #(
    .INIT(32'h69669969)) 
    \n37[7]_i_1__5 
       (.I0(n10[7]),
        .I1(n29[7]),
        .I2(n10[6]),
        .I3(n29[6]),
        .I4(\n37[7]_i_2__5_n_0 ),
        .O(n350_out[7]));
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \n37[7]_i_2__5 
       (.I0(\n37[6]_i_2__5_n_0 ),
        .I1(n29[5]),
        .I2(n10[5]),
        .O(\n37[7]_i_2__5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \n37[8]_i_1__2 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .O(n341_out[0]));
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    \n37[9]_i_1__5 
       (.I0(n21[0]),
        .I1(\n8_reg_n_0_[0] ),
        .I2(n21[1]),
        .I3(\n8_reg_n_0_[1] ),
        .O(n341_out[1]));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[10] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[2]),
        .Q(i1[9]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[11] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[3]),
        .Q(i1[10]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[12] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[4]),
        .Q(i1[11]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[13] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[5]),
        .Q(i1[12]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[14] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[6]),
        .Q(i1[13]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[15] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[7]),
        .Q(i1[14]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[1]),
        .Q(i1[0]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[2]),
        .Q(i1[1]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[3]),
        .Q(i1[2]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[4]),
        .Q(i1[3]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[5]),
        .Q(i1[4]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[6]),
        .Q(i1[5]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n350_out[7]),
        .Q(i1[6]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[8] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[0]),
        .Q(i1[7]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n37_reg[9] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n341_out[1]),
        .Q(i1[8]),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[0]),
        .Q(\n4_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[1]),
        .Q(\n4_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[2]),
        .Q(\n4_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[3]),
        .Q(\n4_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[4]),
        .Q(\n4_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[5]),
        .Q(\n4_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[6]),
        .Q(\n4_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n4_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(s8_3[7]),
        .Q(\n4_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[0]),
        .Q(\n7_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[1]),
        .Q(\n7_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[2]),
        .Q(\n7_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[3]),
        .Q(\n7_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[4]),
        .Q(\n7_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[5]),
        .Q(\n7_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[6]),
        .Q(\n7_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n7_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(n2[7]),
        .Q(\n7_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[0] ),
        .Q(\n8_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[1] ),
        .Q(\n8_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[2] ),
        .Q(\n8_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[3] ),
        .Q(\n8_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[4] ),
        .Q(\n8_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[5] ),
        .Q(\n8_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[6] ),
        .Q(\n8_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n8_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n7_reg_n_0_[7] ),
        .Q(\n8_reg_n_0_[7] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[0] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[0] ),
        .Q(\n9_reg_n_0_[0] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[1] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[1] ),
        .Q(\n9_reg_n_0_[1] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[2] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[2] ),
        .Q(\n9_reg_n_0_[2] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[3] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[3] ),
        .Q(\n9_reg_n_0_[3] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[4] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[4] ),
        .Q(\n9_reg_n_0_[4] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[5] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[5] ),
        .Q(\n9_reg_n_0_[5] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[6] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[6] ),
        .Q(\n9_reg_n_0_[6] ),
        .R(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \n9_reg[7] 
       (.C(clk_i),
        .CE(enable_i),
        .D(\n1_reg_n_0_[7] ),
        .Q(\n9_reg_n_0_[7] ),
        .R(rst_i));
endmodule

(* ORIG_REF_NAME = "cf_fft_512_8_9" *) 
module switch_elements_cf_fft_512_8_9
   (\n9_reg[0] ,
    s6_3,
    rst_i,
    enable_i,
    clk_i,
    s7_3,
    D);
  output [15:0]\n9_reg[0] ;
  output [15:0]s6_3;
  input rst_i;
  input [0:0]enable_i;
  input clk_i;
  input [15:0]s7_3;
  input [15:0]D;

  wire [15:0]D;
  wire clk_i;
  wire [0:0]enable_i;
  wire [0:0]i8;
  wire [15:0]n33;
  wire [15:1]n37;
  wire n4;
  wire [15:0]\n9_reg[0] ;
  wire rst_i;
  wire s29_n_0;
  wire [15:0]s6_3;
  wire [15:0]s7_3;

  switch_elements_cf_fft_512_8_31_4 s25
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i8(i8),
        .n4(n4),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_10 s26
       (.D(D),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .rst_i(rst_i),
        .s7_3(s7_3));
  switch_elements_cf_fft_512_8_26_5 s28
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .i8(i8),
        .\n1_reg[0] (s29_n_0),
        .n4(n4),
        .\n9_reg[0] (\n9_reg[0] ),
        .rst_i(rst_i));
  switch_elements_cf_fft_512_8_27_6 s29
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .i1({n33[15:9],n33[7:0],n37}),
        .i8(i8),
        .\n9_reg[0]_0 (s29_n_0),
        .rst_i(rst_i),
        .s6_3(s6_3));
endmodule

(* ORIG_REF_NAME = "switch_elements3" *) (* dont_touch = "true" *) 
module switch_elements_switch_elements3
   (enable_i,
    clk_i,
    rst_i,
    info_o);
  input [31:0]enable_i;
  input clk_i;
  input rst_i;
  output [31:0]info_o;

  wire \activity_blocks[0].switch3_n_3 ;
  wire clk_i;
  wire [31:0]enable_i;
  wire \enable_s_reg_n_0_[0] ;
  wire \enable_s_reg_n_0_[10] ;
  wire \enable_s_reg_n_0_[11] ;
  wire \enable_s_reg_n_0_[12] ;
  wire \enable_s_reg_n_0_[13] ;
  wire \enable_s_reg_n_0_[14] ;
  wire \enable_s_reg_n_0_[15] ;
  wire \enable_s_reg_n_0_[1] ;
  wire \enable_s_reg_n_0_[2] ;
  wire \enable_s_reg_n_0_[3] ;
  wire \enable_s_reg_n_0_[4] ;
  wire \enable_s_reg_n_0_[5] ;
  wire \enable_s_reg_n_0_[6] ;
  wire \enable_s_reg_n_0_[7] ;
  wire \enable_s_reg_n_0_[8] ;
  wire \enable_s_reg_n_0_[9] ;
  wire [31:0]info_o;
  wire n25__0_carry_i_16__0_n_40;
  wire n25__0_carry_i_16__0_n_41;
  wire n25__0_carry_i_16__0_n_42;
  wire n25__0_carry_i_16__0_n_43;
  wire n25__0_carry_i_16__0_n_44;
  wire n25__0_carry_i_16__0_n_45;
  wire n25__0_carry_i_16__0_n_46;
  wire n25__0_carry_i_16__0_n_47;
  wire n25__0_carry_i_16__1_n_40;
  wire n25__0_carry_i_16__1_n_41;
  wire n25__0_carry_i_16__1_n_42;
  wire n25__0_carry_i_16__1_n_43;
  wire n25__0_carry_i_16__1_n_44;
  wire n25__0_carry_i_16__1_n_45;
  wire n25__0_carry_i_16__1_n_46;
  wire n25__0_carry_i_16__1_n_47;
  wire [31:0]p_6_out;
  wire rst_i;
  wire [7:0]\s1/s2/s2/B ;
  wire [7:0]\s1/s2/s3/B ;
  wire [15:0]\vec32_ot[9] ;
  wire [15:0]NLW_n25__0_carry_i_16__0_CASDOUTA_UNCONNECTED;
  wire [15:0]NLW_n25__0_carry_i_16__0_CASDOUTB_UNCONNECTED;
  wire [1:0]NLW_n25__0_carry_i_16__0_CASDOUTPA_UNCONNECTED;
  wire [1:0]NLW_n25__0_carry_i_16__0_CASDOUTPB_UNCONNECTED;
  wire [15:0]NLW_n25__0_carry_i_16__0_DOUTBDOUT_UNCONNECTED;
  wire [1:0]NLW_n25__0_carry_i_16__0_DOUTPADOUTP_UNCONNECTED;
  wire [1:0]NLW_n25__0_carry_i_16__0_DOUTPBDOUTP_UNCONNECTED;
  wire [15:0]NLW_n25__0_carry_i_16__1_CASDOUTA_UNCONNECTED;
  wire [15:0]NLW_n25__0_carry_i_16__1_CASDOUTB_UNCONNECTED;
  wire [1:0]NLW_n25__0_carry_i_16__1_CASDOUTPA_UNCONNECTED;
  wire [1:0]NLW_n25__0_carry_i_16__1_CASDOUTPB_UNCONNECTED;
  wire [15:0]NLW_n25__0_carry_i_16__1_DOUTBDOUT_UNCONNECTED;
  wire [1:0]NLW_n25__0_carry_i_16__1_DOUTPADOUTP_UNCONNECTED;
  wire [1:0]NLW_n25__0_carry_i_16__1_DOUTPBDOUTP_UNCONNECTED;

  switch_elements_cf_fft_512_8 \activity_blocks[0].switch3 
       (.DOUTADOUT({\s1/s2/s2/B ,n25__0_carry_i_16__0_n_40,n25__0_carry_i_16__0_n_41,n25__0_carry_i_16__0_n_42,n25__0_carry_i_16__0_n_43,n25__0_carry_i_16__0_n_44,n25__0_carry_i_16__0_n_45,n25__0_carry_i_16__0_n_46,n25__0_carry_i_16__0_n_47}),
        .clk_i(clk_i),
        .enable_i(enable_i[3]),
        .enable_s({\vec32_ot[9] ,\enable_s_reg_n_0_[15] ,\enable_s_reg_n_0_[14] ,\enable_s_reg_n_0_[13] ,\enable_s_reg_n_0_[12] ,\enable_s_reg_n_0_[11] ,\enable_s_reg_n_0_[10] ,\enable_s_reg_n_0_[9] ,\enable_s_reg_n_0_[8] ,\enable_s_reg_n_0_[7] ,\enable_s_reg_n_0_[6] ,\enable_s_reg_n_0_[5] ,\enable_s_reg_n_0_[4] ,\enable_s_reg_n_0_[3] ,\enable_s_reg_n_0_[2] ,\enable_s_reg_n_0_[1] ,\enable_s_reg_n_0_[0] }),
        .n14__56_carry({\s1/s2/s3/B ,n25__0_carry_i_16__1_n_40,n25__0_carry_i_16__1_n_41,n25__0_carry_i_16__1_n_42,n25__0_carry_i_16__1_n_43,n25__0_carry_i_16__1_n_44,n25__0_carry_i_16__1_n_45,n25__0_carry_i_16__1_n_46,n25__0_carry_i_16__1_n_47}),
        .p_6_out({p_6_out[31:29],\activity_blocks[0].switch3_n_3 ,p_6_out[27:0]}),
        .rst_i(rst_i));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[0]),
        .Q(\enable_s_reg_n_0_[0] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[10]),
        .Q(\enable_s_reg_n_0_[10] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[11]),
        .Q(\enable_s_reg_n_0_[11] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[12]),
        .Q(\enable_s_reg_n_0_[12] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[13]),
        .Q(\enable_s_reg_n_0_[13] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[14]),
        .Q(\enable_s_reg_n_0_[14] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[15]),
        .Q(\enable_s_reg_n_0_[15] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[16]),
        .Q(\vec32_ot[9] [0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[17]),
        .Q(\vec32_ot[9] [1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[18]),
        .Q(\vec32_ot[9] [2]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[19]),
        .Q(\vec32_ot[9] [3]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[1]),
        .Q(\enable_s_reg_n_0_[1] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[20]),
        .Q(\vec32_ot[9] [4]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[21]),
        .Q(\vec32_ot[9] [5]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[22]),
        .Q(\vec32_ot[9] [6]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[23]),
        .Q(\vec32_ot[9] [7]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[24]),
        .Q(\vec32_ot[9] [8]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[25]),
        .Q(\vec32_ot[9] [9]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[26]),
        .Q(\vec32_ot[9] [10]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[27]),
        .Q(\vec32_ot[9] [11]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[28]),
        .Q(\vec32_ot[9] [12]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[29]),
        .Q(\vec32_ot[9] [13]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[2]),
        .Q(\enable_s_reg_n_0_[2] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[30]),
        .Q(\vec32_ot[9] [14]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[31]),
        .Q(\vec32_ot[9] [15]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[3]),
        .Q(\enable_s_reg_n_0_[3] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[4]),
        .Q(\enable_s_reg_n_0_[4] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[5]),
        .Q(\enable_s_reg_n_0_[5] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[6]),
        .Q(\enable_s_reg_n_0_[6] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[7]),
        .Q(\enable_s_reg_n_0_[7] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[8]),
        .Q(\enable_s_reg_n_0_[8] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \enable_s_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .D(enable_i[9]),
        .Q(\enable_s_reg_n_0_[9] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[0]),
        .Q(info_o[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[10]),
        .Q(info_o[10]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[11]),
        .Q(info_o[11]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[12]),
        .Q(info_o[12]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[13]),
        .Q(info_o[13]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[14]),
        .Q(info_o[14]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[15]),
        .Q(info_o[15]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[16]),
        .Q(info_o[16]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[17]),
        .Q(info_o[17]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[18]),
        .Q(info_o[18]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[19]),
        .Q(info_o[19]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[1]),
        .Q(info_o[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[20]),
        .Q(info_o[20]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[21]),
        .Q(info_o[21]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[22]),
        .Q(info_o[22]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[23]),
        .Q(info_o[23]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[24]),
        .Q(info_o[24]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[25]),
        .Q(info_o[25]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[26]),
        .Q(info_o[26]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[27]),
        .Q(info_o[27]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\activity_blocks[0].switch3_n_3 ),
        .Q(info_o[28]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[29]),
        .Q(info_o[29]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[2]),
        .Q(info_o[2]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[30]),
        .Q(info_o[30]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[31]),
        .Q(info_o[31]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[3]),
        .Q(info_o[3]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[4]),
        .Q(info_o[4]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[5]),
        .Q(info_o[5]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[6]),
        .Q(info_o[6]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[7]),
        .Q(info_o[7]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[8]),
        .Q(info_o[8]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \info_o_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_6_out[9]),
        .Q(info_o[9]),
        .R(1'b0));
  (* \MEM.PORTA.DATA_BIT_LAYOUT  = "p0_d16" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RDADDR_COLLISION_HWCONFIG = "PERFORMANCE" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "15" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "1023" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "15" *) 
  RAMB18E2 #(
    .CASCADE_ORDER_A("NONE"),
    .CASCADE_ORDER_B("NONE"),
    .CLOCK_DOMAINS("INDEPENDENT"),
    .DOA_REG(1),
    .DOB_REG(0),
    .ENADDRENA("FALSE"),
    .ENADDRENB("FALSE"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h77D178D479D77ADA7BDD7CE07CE37DE77EEA7EED7FF07FF37FF67FF97FFC7F00),
    .INIT_01(256'h5CA75EAA60AC62AE64B166B368B66AB86CBB6DBE6FC070C372C673C975CC76CF),
    .INIT_02(256'h338A368C398D3C8F3F9041924493479549974C994E9B519D539F55A158A35AA5),
    .INIT_03(256'h0380068009800C800F801281158118821C831F832284258528862B872E883089),
    .INIT_04(256'hD188D487D786DA85DD84E083E383E782EA81ED81F080F380F680F980FC800080),
    .INIT_05(256'hA7A3AAA1AC9FAE9DB19BB399B697B895BB93BE92C090C38FC68DC98CCC8ACF89),
    .INIT_06(256'h8ACC8CC98DC68FC390C092BE93BB95B897B699B39BB19DAE9FACA1AAA3A7A5A5),
    .INIT_07(256'h80FC80F980F680F380F081ED81EA82E783E383E084DD85DA86D787D488D189CF),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .RDADDRCHANGEA("FALSE"),
    .RDADDRCHANGEB("FALSE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(0),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SLEEP_ASYNC("FALSE"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    n25__0_carry_i_16__0
       (.ADDRARDADDR({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .ADDRBWRADDR({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .ADDRENA(1'b0),
        .ADDRENB(1'b0),
        .CASDIMUXA(1'b0),
        .CASDIMUXB(1'b0),
        .CASDINA({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .CASDINB({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .CASDINPA({1'b0,1'b0}),
        .CASDINPB({1'b0,1'b0}),
        .CASDOMUXA(1'b0),
        .CASDOMUXB(1'b0),
        .CASDOMUXEN_A(1'b1),
        .CASDOMUXEN_B(1'b1),
        .CASDOUTA(NLW_n25__0_carry_i_16__0_CASDOUTA_UNCONNECTED[15:0]),
        .CASDOUTB(NLW_n25__0_carry_i_16__0_CASDOUTB_UNCONNECTED[15:0]),
        .CASDOUTPA(NLW_n25__0_carry_i_16__0_CASDOUTPA_UNCONNECTED[1:0]),
        .CASDOUTPB(NLW_n25__0_carry_i_16__0_CASDOUTPB_UNCONNECTED[1:0]),
        .CASOREGIMUXA(1'b0),
        .CASOREGIMUXB(1'b0),
        .CASOREGIMUXEN_A(1'b1),
        .CASOREGIMUXEN_B(1'b1),
        .CLKARDCLK(clk_i),
        .CLKBWRCLK(1'b0),
        .DINADIN({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DINBDIN({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DINPADINP({1'b0,1'b0}),
        .DINPBDINP({1'b1,1'b1}),
        .DOUTADOUT({\s1/s2/s2/B ,n25__0_carry_i_16__0_n_40,n25__0_carry_i_16__0_n_41,n25__0_carry_i_16__0_n_42,n25__0_carry_i_16__0_n_43,n25__0_carry_i_16__0_n_44,n25__0_carry_i_16__0_n_45,n25__0_carry_i_16__0_n_46,n25__0_carry_i_16__0_n_47}),
        .DOUTBDOUT(NLW_n25__0_carry_i_16__0_DOUTBDOUT_UNCONNECTED[15:0]),
        .DOUTPADOUTP(NLW_n25__0_carry_i_16__0_DOUTPADOUTP_UNCONNECTED[1:0]),
        .DOUTPBDOUTP(NLW_n25__0_carry_i_16__0_DOUTPBDOUTP_UNCONNECTED[1:0]),
        .ENARDEN(rst_i),
        .ENBWREN(1'b0),
        .REGCEAREGCE(enable_i[3]),
        .REGCEB(1'b1),
        .RSTRAMARSTRAM(1'b0),
        .RSTRAMB(1'b0),
        .RSTREGARSTREG(1'b0),
        .RSTREGB(1'b0),
        .SLEEP(1'b0),
        .WEA({1'b0,1'b0}),
        .WEBWE({1'b0,1'b0,1'b0,1'b0}));
  (* \MEM.PORTA.DATA_BIT_LAYOUT  = "p0_d16" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RDADDR_COLLISION_HWCONFIG = "PERFORMANCE" *) 
  (* RTL_RAM_BITS = "1024" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "15" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "1023" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "15" *) 
  RAMB18E2 #(
    .CASCADE_ORDER_A("NONE"),
    .CASCADE_ORDER_B("NONE"),
    .CLOCK_DOMAINS("INDEPENDENT"),
    .DOA_REG(1),
    .DOB_REG(0),
    .ENADDRENA("FALSE"),
    .ENADDRENB("FALSE"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h5EAA62AE66B36AB86DBE70C373C976CF78D47ADA7CE07DE77EED7FF37FF97F00),
    .INIT_01(256'h06800C80128118821F8325852B873089368C3C8F419247954C99519D55A15AA5),
    .INIT_02(256'hAAA1AE9DB399B895BE92C38FC98CCF89D487DA85E083E782ED81F380F9800080),
    .INIT_03(256'h80F980F381ED82E783E085DA87D489CF8CC98FC392BE95B899B39DAEA1AAA5A5),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .RDADDRCHANGEA("FALSE"),
    .RDADDRCHANGEB("FALSE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(0),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SLEEP_ASYNC("FALSE"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    n25__0_carry_i_16__1
       (.ADDRARDADDR({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .ADDRBWRADDR({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .ADDRENA(1'b0),
        .ADDRENB(1'b0),
        .CASDIMUXA(1'b0),
        .CASDIMUXB(1'b0),
        .CASDINA({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .CASDINB({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .CASDINPA({1'b0,1'b0}),
        .CASDINPB({1'b0,1'b0}),
        .CASDOMUXA(1'b0),
        .CASDOMUXB(1'b0),
        .CASDOMUXEN_A(1'b1),
        .CASDOMUXEN_B(1'b1),
        .CASDOUTA(NLW_n25__0_carry_i_16__1_CASDOUTA_UNCONNECTED[15:0]),
        .CASDOUTB(NLW_n25__0_carry_i_16__1_CASDOUTB_UNCONNECTED[15:0]),
        .CASDOUTPA(NLW_n25__0_carry_i_16__1_CASDOUTPA_UNCONNECTED[1:0]),
        .CASDOUTPB(NLW_n25__0_carry_i_16__1_CASDOUTPB_UNCONNECTED[1:0]),
        .CASOREGIMUXA(1'b0),
        .CASOREGIMUXB(1'b0),
        .CASOREGIMUXEN_A(1'b1),
        .CASOREGIMUXEN_B(1'b1),
        .CLKARDCLK(clk_i),
        .CLKBWRCLK(1'b0),
        .DINADIN({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DINBDIN({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DINPADINP({1'b0,1'b0}),
        .DINPBDINP({1'b1,1'b1}),
        .DOUTADOUT({\s1/s2/s3/B ,n25__0_carry_i_16__1_n_40,n25__0_carry_i_16__1_n_41,n25__0_carry_i_16__1_n_42,n25__0_carry_i_16__1_n_43,n25__0_carry_i_16__1_n_44,n25__0_carry_i_16__1_n_45,n25__0_carry_i_16__1_n_46,n25__0_carry_i_16__1_n_47}),
        .DOUTBDOUT(NLW_n25__0_carry_i_16__1_DOUTBDOUT_UNCONNECTED[15:0]),
        .DOUTPADOUTP(NLW_n25__0_carry_i_16__1_DOUTPADOUTP_UNCONNECTED[1:0]),
        .DOUTPBDOUTP(NLW_n25__0_carry_i_16__1_DOUTPBDOUTP_UNCONNECTED[1:0]),
        .ENARDEN(rst_i),
        .ENBWREN(1'b0),
        .REGCEAREGCE(enable_i[3]),
        .REGCEB(1'b1),
        .RSTRAMARSTRAM(1'b0),
        .RSTRAMB(1'b0),
        .RSTREGARSTREG(1'b0),
        .RSTREGB(1'b0),
        .SLEEP(1'b0),
        .WEA({1'b0,1'b0}),
        .WEBWE({1'b0,1'b0,1'b0,1'b0}));
endmodule
`ifndef GLBL
`define GLBL
`timescale  1 ps / 1 ps

module glbl ();

    parameter ROC_WIDTH = 100000;
    parameter TOC_WIDTH = 0;

//--------   STARTUP Globals --------------
    wire GSR;
    wire GTS;
    wire GWE;
    wire PRLD;
    tri1 p_up_tmp;
    tri (weak1, strong0) PLL_LOCKG = p_up_tmp;

    wire PROGB_GLBL;
    wire CCLKO_GLBL;
    wire FCSBO_GLBL;
    wire [3:0] DO_GLBL;
    wire [3:0] DI_GLBL;
   
    reg GSR_int;
    reg GTS_int;
    reg PRLD_int;

//--------   JTAG Globals --------------
    wire JTAG_TDO_GLBL;
    wire JTAG_TCK_GLBL;
    wire JTAG_TDI_GLBL;
    wire JTAG_TMS_GLBL;
    wire JTAG_TRST_GLBL;

    reg JTAG_CAPTURE_GLBL;
    reg JTAG_RESET_GLBL;
    reg JTAG_SHIFT_GLBL;
    reg JTAG_UPDATE_GLBL;
    reg JTAG_RUNTEST_GLBL;

    reg JTAG_SEL1_GLBL = 0;
    reg JTAG_SEL2_GLBL = 0 ;
    reg JTAG_SEL3_GLBL = 0;
    reg JTAG_SEL4_GLBL = 0;

    reg JTAG_USER_TDO1_GLBL = 1'bz;
    reg JTAG_USER_TDO2_GLBL = 1'bz;
    reg JTAG_USER_TDO3_GLBL = 1'bz;
    reg JTAG_USER_TDO4_GLBL = 1'bz;

    assign (strong1, weak0) GSR = GSR_int;
    assign (strong1, weak0) GTS = GTS_int;
    assign (weak1, weak0) PRLD = PRLD_int;

    initial begin
	GSR_int = 1'b1;
	PRLD_int = 1'b1;
	#(ROC_WIDTH)
	GSR_int = 1'b0;
	PRLD_int = 1'b0;
    end

    initial begin
	GTS_int = 1'b1;
	#(TOC_WIDTH)
	GTS_int = 1'b0;
    end

endmodule
`endif
