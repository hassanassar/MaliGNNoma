`timescale 1 ps / 1 ps
`define XIL_TIMING

(* dont_touch = "true" *) 
(* NotValidForBitStream *)
module switch_elements
   (enable_i,
    clk_i,
    rst_i,
    info_o);
  input [31:0]enable_i;
  input clk_i;
  input rst_i;
  output [31:0]info_o;

  wire \<const0> ;
  wire clk_i;
  wire [31:0]enable_i;
  wire [31:0]\^info_o ;
  wire \info_o[0]_INST_0_i_8_n_0 ;
  wire \info_o[2]_INST_0_i_4_n_0 ;
  wire \info_o[3]_INST_0_i_2_n_0 ;
  wire rst_i;

  assign info_o[31:6] = \^info_o [31:6];
  assign info_o[5] = \<const0> ;
  assign info_o[4:0] = \^info_o [4:0];
  GND GND
       (.G(\<const0> ));
  (* SOFT_HLUTNM = "soft_lutpair313" *) 
  LUT4 #(
    .INIT(16'hEFFF)) 
    \info_o[0]_INST_0_i_8 
       (.I0(enable_i[3]),
        .I1(enable_i[4]),
        .I2(enable_i[6]),
        .I3(enable_i[0]),
        .O(\info_o[0]_INST_0_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair313" *) 
  LUT3 #(
    .INIT(8'hFD)) 
    \info_o[2]_INST_0_i_4 
       (.I0(enable_i[6]),
        .I1(enable_i[4]),
        .I2(enable_i[3]),
        .O(\info_o[2]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \info_o[3]_INST_0_i_2 
       (.I0(enable_i[0]),
        .I1(enable_i[1]),
        .I2(enable_i[2]),
        .I3(enable_i[3]),
        .I4(enable_i[4]),
        .I5(enable_i[6]),
        .O(\info_o[3]_INST_0_i_2_n_0 ));
  switch_elements_aes_ip switch
       (.clk_i(clk_i),
        .enable_i(enable_i),
        .info_o({\^info_o [31:6],\^info_o [4:0]}),
        .\info_o[0]_INST_0_i_4 (\info_o[0]_INST_0_i_8_n_0 ),
        .info_o_2_sp_1(\info_o[2]_INST_0_i_4_n_0 ),
        .info_o_3_sp_1(\info_o[3]_INST_0_i_2_n_0 ),
        .rst_i(rst_i));
endmodule

(* ORIG_REF_NAME = "aes_core" *) 
module switch_elements_aes_core
   (info_o,
    \KR[1].key_reg[2][12] ,
    enable_i_0_sp_1,
    \aes_cr_reg[2] ,
    ccf_reg,
    Q,
    \FSM_sequential_state_reg[2] ,
    \FSM_sequential_state_reg[3] ,
    \FSM_sequential_state_reg[2]_0 ,
    \FSM_sequential_state_reg[0] ,
    enable_i_6_sp_1,
    enable_i_3_sp_1,
    \enable_i[6]_0 ,
    \rd_count_reg[3] ,
    \rd_count_reg[2] ,
    \FSM_sequential_state_reg[2]_1 ,
    \aes_cr_reg[4] ,
    \FSM_sequential_state_reg[3]_0 ,
    \FSM_sequential_state_reg[3]_1 ,
    enable_i_2_sp_1,
    \FSM_sequential_state_reg[2]_2 ,
    bypass_rk,
    \CD[2].col_reg[1][31] ,
    last_round_pp2_reg,
    bus_swap,
    \FSM_sequential_state_reg[0]_0 ,
    data_in,
    iv_mux_out16_out,
    \col_en_cnt_unit_pp2_reg[3] ,
    \aes_cr_reg[5] ,
    \aes_cr_reg[5]_0 ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][31] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][31] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][31] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][31] ,
    clk_i,
    rst_i,
    rk_out_sel,
    \info_o[31] ,
    \info_o[31]_0 ,
    info_o_0_sp_1,
    \FSM_sequential_state_reg[3]_2 ,
    \info_o[0]_0 ,
    info_o_4_sp_1,
    info_o_6_sp_1,
    info_o_9_sp_1,
    info_o_10_sp_1,
    info_o_11_sp_1,
    info_o_12_sp_1,
    \FSM_sequential_state_reg[0]_1 ,
    \col_en_cnt_unit_pp1_reg[3] ,
    \FSM_sequential_state_reg[2]_3 ,
    enable_i,
    ccf,
    ccf_reg_0,
    \col_sel_pp1_reg[1] ,
    \info_o[0]_1 ,
    \key_en_pp1_reg[3] ,
    \FSM_sequential_state_reg[3]_3 ,
    \FSM_sequential_state_reg[3]_4 ,
    \FSM_sequential_state_reg[0]_2 ,
    \FSM_sequential_state_reg[0]_3 ,
    \sbox_pp2_reg[31] ,
    key_en,
    D,
    \IV_BKP_REGISTERS[3].bkp_reg[3][0] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][31] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][0] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][0] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][0] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][31] ,
    \CD[0].col[3][0]_i_2 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][1] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][1] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][1] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][1] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][2] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][2] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][2] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][2] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][3] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][3] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][3] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][3] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][4] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][4] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][4] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][4] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][5] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][5] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][5] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][5] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][6] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][6] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][6] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][6] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][7] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][7] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][7] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][7] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][8] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][8] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][9] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][9] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][10] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][10] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][11] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][11] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][12] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][12] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][13] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][13] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][14] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][14] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][15] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][15] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][16] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][16] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][16] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][16] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][17] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][17] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][17] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][17] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][18] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][18] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][18] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][18] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][19] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][19] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][19] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][19] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][20] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][20] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][20] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][20] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][21] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][21] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][21] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][21] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][22] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][22] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][22] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][22] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][23] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][23] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][23] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][23] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][24] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][24] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][25] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][25] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][26] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][26] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][27] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][27] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][28] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][28] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][29] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][29] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][30] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][30] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][31] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 ,
    \CD[0].col[3][5]_i_2 ,
    \CD[0].col[3][0]_i_2_0 ,
    \CD[0].col[3][10]_i_6 ,
    \CD[0].col[3][0]_i_4 ,
    first_block,
    col_en_host,
    \CD[0].col[3][31]_i_22 ,
    \CD[3].col_reg[0][31] ,
    \CD[3].col_reg[0][31]_0 ,
    \CD[0].col[3][10]_i_12 ,
    \KR[3].key_reg[0][31] ,
    key_sel_rd,
    key_derivation_en,
    \info_o[28]_INST_0_i_15 ,
    \info_o[28]_INST_0_i_15_0 ,
    \info_o[31]_INST_0_i_12 ,
    \FSM_sequential_state_reg[1] ,
    E,
    \KR[1].key_host_reg[2][0] ,
    \KR[2].key_host_reg[1][0] ,
    \KR[3].key_host_reg[0][0] ,
    \IV_BKP_REGISTERS[3].iv_reg[3][0] ,
    iv_en,
    \IV_BKP_REGISTERS[3].bkp_reg[3][0]_0 ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][31] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][15] ,
    enc_dec);
  output [27:0]info_o;
  output [5:0]\KR[1].key_reg[2][12] ;
  output enable_i_0_sp_1;
  output [2:0]\aes_cr_reg[2] ;
  output ccf_reg;
  output [3:0]Q;
  output \FSM_sequential_state_reg[2] ;
  output \FSM_sequential_state_reg[3] ;
  output \FSM_sequential_state_reg[2]_0 ;
  output \FSM_sequential_state_reg[0] ;
  output enable_i_6_sp_1;
  output enable_i_3_sp_1;
  output \enable_i[6]_0 ;
  output \rd_count_reg[3] ;
  output [0:0]\rd_count_reg[2] ;
  output [0:0]\FSM_sequential_state_reg[2]_1 ;
  output \aes_cr_reg[4] ;
  output \FSM_sequential_state_reg[3]_0 ;
  output \FSM_sequential_state_reg[3]_1 ;
  output enable_i_2_sp_1;
  output \FSM_sequential_state_reg[2]_2 ;
  output bypass_rk;
  output [31:0]\CD[2].col_reg[1][31] ;
  output [15:0]last_round_pp2_reg;
  output [31:0]bus_swap;
  output \FSM_sequential_state_reg[0]_0 ;
  output [15:0]data_in;
  output iv_mux_out16_out;
  output [3:0]\col_en_cnt_unit_pp2_reg[3] ;
  output \aes_cr_reg[5] ;
  output \aes_cr_reg[5]_0 ;
  output [31:0]\IV_BKP_REGISTERS[3].bkp_1_reg[3][31] ;
  output [31:0]\IV_BKP_REGISTERS[2].bkp_1_reg[2][31] ;
  output [31:0]\IV_BKP_REGISTERS[1].bkp_1_reg[1][31] ;
  output [31:0]\IV_BKP_REGISTERS[0].bkp_1_reg[0][31] ;
  input clk_i;
  input rst_i;
  input rk_out_sel;
  input \info_o[31] ;
  input \info_o[31]_0 ;
  input info_o_0_sp_1;
  input \FSM_sequential_state_reg[3]_2 ;
  input \info_o[0]_0 ;
  input info_o_4_sp_1;
  input info_o_6_sp_1;
  input info_o_9_sp_1;
  input info_o_10_sp_1;
  input info_o_11_sp_1;
  input info_o_12_sp_1;
  input \FSM_sequential_state_reg[0]_1 ;
  input \col_en_cnt_unit_pp1_reg[3] ;
  input \FSM_sequential_state_reg[2]_3 ;
  input [31:0]enable_i;
  input ccf;
  input ccf_reg_0;
  input \col_sel_pp1_reg[1] ;
  input [6:0]\info_o[0]_1 ;
  input \key_en_pp1_reg[3] ;
  input \FSM_sequential_state_reg[3]_3 ;
  input \FSM_sequential_state_reg[3]_4 ;
  input \FSM_sequential_state_reg[0]_2 ;
  input \FSM_sequential_state_reg[0]_3 ;
  input \sbox_pp2_reg[31] ;
  input [3:0]key_en;
  input [7:0]D;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][0] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][31] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][0] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][0] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][0] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][31] ;
  input \CD[0].col[3][0]_i_2 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][1] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][1] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][1] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][1] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][2] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][2] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][2] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][2] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][3] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][3] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][3] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][3] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][4] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][4] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][4] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][4] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][5] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][5] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][5] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][5] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][6] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][6] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][6] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][6] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][7] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][7] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][7] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][7] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][8] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][8] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][9] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][9] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][10] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][10] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][11] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][11] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][12] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][12] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][13] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][13] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][14] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][14] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][15] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][15] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][16] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][16] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][16] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][16] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][17] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][17] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][17] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][17] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][18] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][18] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][18] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][18] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][19] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][19] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][19] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][19] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][20] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][20] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][20] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][20] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][21] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][21] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][21] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][21] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][22] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][22] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][22] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][22] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][23] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][23] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][23] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][23] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][24] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][24] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][25] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][25] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][26] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][26] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][27] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][27] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][28] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][28] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][29] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][29] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][30] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][30] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][31] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 ;
  input \CD[0].col[3][5]_i_2 ;
  input \CD[0].col[3][0]_i_2_0 ;
  input \CD[0].col[3][10]_i_6 ;
  input \CD[0].col[3][0]_i_4 ;
  input first_block;
  input [3:0]col_en_host;
  input \CD[0].col[3][31]_i_22 ;
  input [1:0]\CD[3].col_reg[0][31] ;
  input \CD[3].col_reg[0][31]_0 ;
  input \CD[0].col[3][10]_i_12 ;
  input \KR[3].key_reg[0][31] ;
  input [0:0]key_sel_rd;
  input key_derivation_en;
  input \info_o[28]_INST_0_i_15 ;
  input \info_o[28]_INST_0_i_15_0 ;
  input \info_o[31]_INST_0_i_12 ;
  input [0:0]\FSM_sequential_state_reg[1] ;
  input [0:0]E;
  input [0:0]\KR[1].key_host_reg[2][0] ;
  input [0:0]\KR[2].key_host_reg[1][0] ;
  input [0:0]\KR[3].key_host_reg[0][0] ;
  input [0:0]\IV_BKP_REGISTERS[3].iv_reg[3][0] ;
  input [2:0]iv_en;
  input [0:0]\IV_BKP_REGISTERS[3].bkp_reg[3][0]_0 ;
  input [0:0]\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ;
  input [7:0]\IV_BKP_REGISTERS[2].bkp_reg[2][31] ;
  input [0:0]\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ;
  input [7:0]\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 ;
  input [0:0]\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ;
  input [7:0]\IV_BKP_REGISTERS[0].bkp_reg[0][15] ;
  input enc_dec;

  wire AES_CORE_CONTROL_UNIT_n_100;
  wire AES_CORE_CONTROL_UNIT_n_101;
  wire AES_CORE_CONTROL_UNIT_n_102;
  wire AES_CORE_CONTROL_UNIT_n_103;
  wire AES_CORE_CONTROL_UNIT_n_104;
  wire AES_CORE_CONTROL_UNIT_n_105;
  wire AES_CORE_CONTROL_UNIT_n_106;
  wire AES_CORE_CONTROL_UNIT_n_107;
  wire AES_CORE_CONTROL_UNIT_n_108;
  wire AES_CORE_CONTROL_UNIT_n_109;
  wire AES_CORE_CONTROL_UNIT_n_110;
  wire AES_CORE_CONTROL_UNIT_n_111;
  wire AES_CORE_CONTROL_UNIT_n_112;
  wire AES_CORE_CONTROL_UNIT_n_113;
  wire AES_CORE_CONTROL_UNIT_n_114;
  wire AES_CORE_CONTROL_UNIT_n_115;
  wire AES_CORE_CONTROL_UNIT_n_116;
  wire AES_CORE_CONTROL_UNIT_n_117;
  wire AES_CORE_CONTROL_UNIT_n_118;
  wire AES_CORE_CONTROL_UNIT_n_119;
  wire AES_CORE_CONTROL_UNIT_n_120;
  wire AES_CORE_CONTROL_UNIT_n_121;
  wire AES_CORE_CONTROL_UNIT_n_122;
  wire AES_CORE_CONTROL_UNIT_n_123;
  wire AES_CORE_CONTROL_UNIT_n_124;
  wire AES_CORE_CONTROL_UNIT_n_125;
  wire AES_CORE_CONTROL_UNIT_n_126;
  wire AES_CORE_CONTROL_UNIT_n_127;
  wire AES_CORE_CONTROL_UNIT_n_128;
  wire AES_CORE_CONTROL_UNIT_n_129;
  wire AES_CORE_CONTROL_UNIT_n_130;
  wire AES_CORE_CONTROL_UNIT_n_131;
  wire AES_CORE_CONTROL_UNIT_n_132;
  wire AES_CORE_CONTROL_UNIT_n_133;
  wire AES_CORE_CONTROL_UNIT_n_134;
  wire AES_CORE_CONTROL_UNIT_n_135;
  wire AES_CORE_CONTROL_UNIT_n_136;
  wire AES_CORE_CONTROL_UNIT_n_137;
  wire AES_CORE_CONTROL_UNIT_n_138;
  wire AES_CORE_CONTROL_UNIT_n_139;
  wire AES_CORE_CONTROL_UNIT_n_140;
  wire AES_CORE_CONTROL_UNIT_n_141;
  wire AES_CORE_CONTROL_UNIT_n_142;
  wire AES_CORE_CONTROL_UNIT_n_143;
  wire AES_CORE_CONTROL_UNIT_n_144;
  wire AES_CORE_CONTROL_UNIT_n_145;
  wire AES_CORE_CONTROL_UNIT_n_146;
  wire AES_CORE_CONTROL_UNIT_n_147;
  wire AES_CORE_CONTROL_UNIT_n_148;
  wire AES_CORE_CONTROL_UNIT_n_149;
  wire AES_CORE_CONTROL_UNIT_n_150;
  wire AES_CORE_CONTROL_UNIT_n_151;
  wire AES_CORE_CONTROL_UNIT_n_152;
  wire AES_CORE_CONTROL_UNIT_n_153;
  wire AES_CORE_CONTROL_UNIT_n_154;
  wire AES_CORE_CONTROL_UNIT_n_155;
  wire AES_CORE_CONTROL_UNIT_n_156;
  wire AES_CORE_CONTROL_UNIT_n_157;
  wire AES_CORE_CONTROL_UNIT_n_158;
  wire AES_CORE_CONTROL_UNIT_n_159;
  wire AES_CORE_CONTROL_UNIT_n_160;
  wire AES_CORE_CONTROL_UNIT_n_161;
  wire AES_CORE_CONTROL_UNIT_n_194;
  wire AES_CORE_CONTROL_UNIT_n_195;
  wire AES_CORE_CONTROL_UNIT_n_196;
  wire AES_CORE_CONTROL_UNIT_n_197;
  wire AES_CORE_CONTROL_UNIT_n_198;
  wire AES_CORE_CONTROL_UNIT_n_199;
  wire AES_CORE_CONTROL_UNIT_n_200;
  wire AES_CORE_CONTROL_UNIT_n_201;
  wire AES_CORE_CONTROL_UNIT_n_202;
  wire AES_CORE_CONTROL_UNIT_n_203;
  wire AES_CORE_CONTROL_UNIT_n_204;
  wire AES_CORE_CONTROL_UNIT_n_205;
  wire AES_CORE_CONTROL_UNIT_n_206;
  wire AES_CORE_CONTROL_UNIT_n_207;
  wire AES_CORE_CONTROL_UNIT_n_208;
  wire AES_CORE_CONTROL_UNIT_n_209;
  wire AES_CORE_CONTROL_UNIT_n_210;
  wire AES_CORE_CONTROL_UNIT_n_211;
  wire AES_CORE_CONTROL_UNIT_n_212;
  wire AES_CORE_CONTROL_UNIT_n_213;
  wire AES_CORE_CONTROL_UNIT_n_214;
  wire AES_CORE_CONTROL_UNIT_n_215;
  wire AES_CORE_CONTROL_UNIT_n_216;
  wire AES_CORE_CONTROL_UNIT_n_217;
  wire AES_CORE_CONTROL_UNIT_n_218;
  wire AES_CORE_CONTROL_UNIT_n_219;
  wire AES_CORE_CONTROL_UNIT_n_220;
  wire AES_CORE_CONTROL_UNIT_n_221;
  wire AES_CORE_CONTROL_UNIT_n_222;
  wire AES_CORE_CONTROL_UNIT_n_223;
  wire AES_CORE_CONTROL_UNIT_n_224;
  wire AES_CORE_CONTROL_UNIT_n_225;
  wire AES_CORE_CONTROL_UNIT_n_226;
  wire AES_CORE_CONTROL_UNIT_n_227;
  wire AES_CORE_CONTROL_UNIT_n_228;
  wire AES_CORE_CONTROL_UNIT_n_229;
  wire AES_CORE_CONTROL_UNIT_n_230;
  wire AES_CORE_CONTROL_UNIT_n_231;
  wire AES_CORE_CONTROL_UNIT_n_232;
  wire AES_CORE_CONTROL_UNIT_n_233;
  wire AES_CORE_CONTROL_UNIT_n_234;
  wire AES_CORE_CONTROL_UNIT_n_235;
  wire AES_CORE_CONTROL_UNIT_n_236;
  wire AES_CORE_CONTROL_UNIT_n_237;
  wire AES_CORE_CONTROL_UNIT_n_238;
  wire AES_CORE_CONTROL_UNIT_n_239;
  wire AES_CORE_CONTROL_UNIT_n_240;
  wire AES_CORE_CONTROL_UNIT_n_241;
  wire AES_CORE_CONTROL_UNIT_n_242;
  wire AES_CORE_CONTROL_UNIT_n_243;
  wire AES_CORE_CONTROL_UNIT_n_244;
  wire AES_CORE_CONTROL_UNIT_n_245;
  wire AES_CORE_CONTROL_UNIT_n_246;
  wire AES_CORE_CONTROL_UNIT_n_247;
  wire AES_CORE_CONTROL_UNIT_n_248;
  wire AES_CORE_CONTROL_UNIT_n_249;
  wire AES_CORE_CONTROL_UNIT_n_250;
  wire AES_CORE_CONTROL_UNIT_n_251;
  wire AES_CORE_CONTROL_UNIT_n_252;
  wire AES_CORE_CONTROL_UNIT_n_253;
  wire AES_CORE_CONTROL_UNIT_n_254;
  wire AES_CORE_CONTROL_UNIT_n_255;
  wire AES_CORE_CONTROL_UNIT_n_256;
  wire AES_CORE_CONTROL_UNIT_n_257;
  wire AES_CORE_CONTROL_UNIT_n_258;
  wire AES_CORE_CONTROL_UNIT_n_259;
  wire AES_CORE_CONTROL_UNIT_n_260;
  wire AES_CORE_CONTROL_UNIT_n_261;
  wire AES_CORE_CONTROL_UNIT_n_262;
  wire AES_CORE_CONTROL_UNIT_n_263;
  wire AES_CORE_CONTROL_UNIT_n_264;
  wire AES_CORE_CONTROL_UNIT_n_265;
  wire AES_CORE_CONTROL_UNIT_n_266;
  wire AES_CORE_CONTROL_UNIT_n_267;
  wire AES_CORE_CONTROL_UNIT_n_268;
  wire AES_CORE_CONTROL_UNIT_n_269;
  wire AES_CORE_CONTROL_UNIT_n_270;
  wire AES_CORE_CONTROL_UNIT_n_271;
  wire AES_CORE_CONTROL_UNIT_n_272;
  wire AES_CORE_CONTROL_UNIT_n_273;
  wire AES_CORE_CONTROL_UNIT_n_274;
  wire AES_CORE_CONTROL_UNIT_n_275;
  wire AES_CORE_CONTROL_UNIT_n_276;
  wire AES_CORE_CONTROL_UNIT_n_277;
  wire AES_CORE_CONTROL_UNIT_n_278;
  wire AES_CORE_CONTROL_UNIT_n_279;
  wire AES_CORE_CONTROL_UNIT_n_28;
  wire AES_CORE_CONTROL_UNIT_n_280;
  wire AES_CORE_CONTROL_UNIT_n_281;
  wire AES_CORE_CONTROL_UNIT_n_282;
  wire AES_CORE_CONTROL_UNIT_n_283;
  wire AES_CORE_CONTROL_UNIT_n_284;
  wire AES_CORE_CONTROL_UNIT_n_285;
  wire AES_CORE_CONTROL_UNIT_n_286;
  wire AES_CORE_CONTROL_UNIT_n_287;
  wire AES_CORE_CONTROL_UNIT_n_288;
  wire AES_CORE_CONTROL_UNIT_n_289;
  wire AES_CORE_CONTROL_UNIT_n_291;
  wire AES_CORE_CONTROL_UNIT_n_292;
  wire AES_CORE_CONTROL_UNIT_n_298;
  wire AES_CORE_CONTROL_UNIT_n_299;
  wire AES_CORE_CONTROL_UNIT_n_300;
  wire AES_CORE_CONTROL_UNIT_n_301;
  wire AES_CORE_CONTROL_UNIT_n_302;
  wire AES_CORE_CONTROL_UNIT_n_303;
  wire AES_CORE_CONTROL_UNIT_n_304;
  wire AES_CORE_CONTROL_UNIT_n_305;
  wire AES_CORE_CONTROL_UNIT_n_306;
  wire AES_CORE_CONTROL_UNIT_n_307;
  wire AES_CORE_CONTROL_UNIT_n_308;
  wire AES_CORE_CONTROL_UNIT_n_309;
  wire AES_CORE_CONTROL_UNIT_n_310;
  wire AES_CORE_CONTROL_UNIT_n_311;
  wire AES_CORE_CONTROL_UNIT_n_312;
  wire AES_CORE_CONTROL_UNIT_n_313;
  wire AES_CORE_CONTROL_UNIT_n_314;
  wire AES_CORE_CONTROL_UNIT_n_315;
  wire AES_CORE_CONTROL_UNIT_n_316;
  wire AES_CORE_CONTROL_UNIT_n_317;
  wire AES_CORE_CONTROL_UNIT_n_318;
  wire AES_CORE_CONTROL_UNIT_n_319;
  wire AES_CORE_CONTROL_UNIT_n_320;
  wire AES_CORE_CONTROL_UNIT_n_321;
  wire AES_CORE_CONTROL_UNIT_n_322;
  wire AES_CORE_CONTROL_UNIT_n_323;
  wire AES_CORE_CONTROL_UNIT_n_324;
  wire AES_CORE_CONTROL_UNIT_n_325;
  wire AES_CORE_CONTROL_UNIT_n_326;
  wire AES_CORE_CONTROL_UNIT_n_327;
  wire AES_CORE_CONTROL_UNIT_n_328;
  wire AES_CORE_CONTROL_UNIT_n_329;
  wire AES_CORE_CONTROL_UNIT_n_330;
  wire AES_CORE_CONTROL_UNIT_n_331;
  wire AES_CORE_CONTROL_UNIT_n_332;
  wire AES_CORE_CONTROL_UNIT_n_333;
  wire AES_CORE_CONTROL_UNIT_n_334;
  wire AES_CORE_CONTROL_UNIT_n_335;
  wire AES_CORE_CONTROL_UNIT_n_336;
  wire AES_CORE_CONTROL_UNIT_n_337;
  wire AES_CORE_CONTROL_UNIT_n_338;
  wire AES_CORE_CONTROL_UNIT_n_339;
  wire AES_CORE_CONTROL_UNIT_n_340;
  wire AES_CORE_CONTROL_UNIT_n_341;
  wire AES_CORE_CONTROL_UNIT_n_342;
  wire AES_CORE_CONTROL_UNIT_n_343;
  wire AES_CORE_CONTROL_UNIT_n_344;
  wire AES_CORE_CONTROL_UNIT_n_345;
  wire AES_CORE_CONTROL_UNIT_n_346;
  wire AES_CORE_CONTROL_UNIT_n_347;
  wire AES_CORE_CONTROL_UNIT_n_348;
  wire AES_CORE_CONTROL_UNIT_n_349;
  wire AES_CORE_CONTROL_UNIT_n_350;
  wire AES_CORE_CONTROL_UNIT_n_351;
  wire AES_CORE_CONTROL_UNIT_n_352;
  wire AES_CORE_CONTROL_UNIT_n_353;
  wire AES_CORE_CONTROL_UNIT_n_354;
  wire AES_CORE_CONTROL_UNIT_n_355;
  wire AES_CORE_CONTROL_UNIT_n_356;
  wire AES_CORE_CONTROL_UNIT_n_357;
  wire AES_CORE_CONTROL_UNIT_n_358;
  wire AES_CORE_CONTROL_UNIT_n_359;
  wire AES_CORE_CONTROL_UNIT_n_360;
  wire AES_CORE_CONTROL_UNIT_n_361;
  wire AES_CORE_CONTROL_UNIT_n_362;
  wire AES_CORE_CONTROL_UNIT_n_363;
  wire AES_CORE_CONTROL_UNIT_n_364;
  wire AES_CORE_CONTROL_UNIT_n_365;
  wire AES_CORE_CONTROL_UNIT_n_366;
  wire AES_CORE_CONTROL_UNIT_n_367;
  wire AES_CORE_CONTROL_UNIT_n_368;
  wire AES_CORE_CONTROL_UNIT_n_369;
  wire AES_CORE_CONTROL_UNIT_n_370;
  wire AES_CORE_CONTROL_UNIT_n_371;
  wire AES_CORE_CONTROL_UNIT_n_372;
  wire AES_CORE_CONTROL_UNIT_n_373;
  wire AES_CORE_CONTROL_UNIT_n_374;
  wire AES_CORE_CONTROL_UNIT_n_377;
  wire AES_CORE_CONTROL_UNIT_n_378;
  wire AES_CORE_CONTROL_UNIT_n_379;
  wire AES_CORE_CONTROL_UNIT_n_380;
  wire AES_CORE_CONTROL_UNIT_n_381;
  wire AES_CORE_CONTROL_UNIT_n_382;
  wire AES_CORE_CONTROL_UNIT_n_383;
  wire AES_CORE_CONTROL_UNIT_n_384;
  wire AES_CORE_CONTROL_UNIT_n_385;
  wire AES_CORE_CONTROL_UNIT_n_386;
  wire AES_CORE_CONTROL_UNIT_n_387;
  wire AES_CORE_CONTROL_UNIT_n_388;
  wire AES_CORE_CONTROL_UNIT_n_392;
  wire AES_CORE_CONTROL_UNIT_n_394;
  wire AES_CORE_CONTROL_UNIT_n_395;
  wire AES_CORE_CONTROL_UNIT_n_402;
  wire AES_CORE_CONTROL_UNIT_n_403;
  wire AES_CORE_CONTROL_UNIT_n_404;
  wire AES_CORE_CONTROL_UNIT_n_405;
  wire AES_CORE_CONTROL_UNIT_n_406;
  wire AES_CORE_CONTROL_UNIT_n_407;
  wire AES_CORE_CONTROL_UNIT_n_408;
  wire AES_CORE_CONTROL_UNIT_n_409;
  wire AES_CORE_CONTROL_UNIT_n_410;
  wire AES_CORE_CONTROL_UNIT_n_411;
  wire AES_CORE_CONTROL_UNIT_n_412;
  wire AES_CORE_CONTROL_UNIT_n_413;
  wire AES_CORE_CONTROL_UNIT_n_414;
  wire AES_CORE_CONTROL_UNIT_n_415;
  wire AES_CORE_CONTROL_UNIT_n_416;
  wire AES_CORE_CONTROL_UNIT_n_417;
  wire AES_CORE_CONTROL_UNIT_n_418;
  wire AES_CORE_CONTROL_UNIT_n_419;
  wire AES_CORE_CONTROL_UNIT_n_420;
  wire AES_CORE_CONTROL_UNIT_n_421;
  wire AES_CORE_CONTROL_UNIT_n_422;
  wire AES_CORE_CONTROL_UNIT_n_423;
  wire AES_CORE_CONTROL_UNIT_n_424;
  wire AES_CORE_CONTROL_UNIT_n_425;
  wire AES_CORE_CONTROL_UNIT_n_426;
  wire AES_CORE_CONTROL_UNIT_n_427;
  wire AES_CORE_CONTROL_UNIT_n_428;
  wire AES_CORE_CONTROL_UNIT_n_429;
  wire AES_CORE_CONTROL_UNIT_n_430;
  wire AES_CORE_CONTROL_UNIT_n_431;
  wire AES_CORE_CONTROL_UNIT_n_432;
  wire AES_CORE_CONTROL_UNIT_n_433;
  wire AES_CORE_CONTROL_UNIT_n_434;
  wire AES_CORE_CONTROL_UNIT_n_436;
  wire AES_CORE_CONTROL_UNIT_n_437;
  wire AES_CORE_CONTROL_UNIT_n_438;
  wire AES_CORE_CONTROL_UNIT_n_90;
  wire AES_CORE_CONTROL_UNIT_n_91;
  wire AES_CORE_CONTROL_UNIT_n_92;
  wire AES_CORE_CONTROL_UNIT_n_93;
  wire AES_CORE_CONTROL_UNIT_n_94;
  wire AES_CORE_CONTROL_UNIT_n_95;
  wire AES_CORE_CONTROL_UNIT_n_96;
  wire AES_CORE_CONTROL_UNIT_n_97;
  wire AES_CORE_CONTROL_UNIT_n_98;
  wire AES_CORE_CONTROL_UNIT_n_99;
  wire AES_CORE_DATAPATH_n_126;
  wire AES_CORE_DATAPATH_n_127;
  wire AES_CORE_DATAPATH_n_128;
  wire AES_CORE_DATAPATH_n_129;
  wire AES_CORE_DATAPATH_n_130;
  wire AES_CORE_DATAPATH_n_131;
  wire AES_CORE_DATAPATH_n_132;
  wire AES_CORE_DATAPATH_n_144;
  wire AES_CORE_DATAPATH_n_145;
  wire AES_CORE_DATAPATH_n_146;
  wire AES_CORE_DATAPATH_n_147;
  wire AES_CORE_DATAPATH_n_148;
  wire AES_CORE_DATAPATH_n_149;
  wire AES_CORE_DATAPATH_n_150;
  wire AES_CORE_DATAPATH_n_151;
  wire AES_CORE_DATAPATH_n_152;
  wire AES_CORE_DATAPATH_n_153;
  wire AES_CORE_DATAPATH_n_154;
  wire AES_CORE_DATAPATH_n_155;
  wire AES_CORE_DATAPATH_n_156;
  wire AES_CORE_DATAPATH_n_157;
  wire AES_CORE_DATAPATH_n_158;
  wire AES_CORE_DATAPATH_n_159;
  wire AES_CORE_DATAPATH_n_160;
  wire AES_CORE_DATAPATH_n_161;
  wire AES_CORE_DATAPATH_n_162;
  wire AES_CORE_DATAPATH_n_163;
  wire AES_CORE_DATAPATH_n_164;
  wire AES_CORE_DATAPATH_n_165;
  wire AES_CORE_DATAPATH_n_166;
  wire AES_CORE_DATAPATH_n_167;
  wire AES_CORE_DATAPATH_n_168;
  wire AES_CORE_DATAPATH_n_169;
  wire AES_CORE_DATAPATH_n_170;
  wire AES_CORE_DATAPATH_n_171;
  wire AES_CORE_DATAPATH_n_172;
  wire AES_CORE_DATAPATH_n_173;
  wire AES_CORE_DATAPATH_n_174;
  wire AES_CORE_DATAPATH_n_175;
  wire AES_CORE_DATAPATH_n_176;
  wire AES_CORE_DATAPATH_n_177;
  wire AES_CORE_DATAPATH_n_178;
  wire AES_CORE_DATAPATH_n_2;
  wire AES_CORE_DATAPATH_n_325;
  wire AES_CORE_DATAPATH_n_35;
  wire AES_CORE_DATAPATH_n_36;
  wire AES_CORE_DATAPATH_n_37;
  wire AES_CORE_DATAPATH_n_38;
  wire AES_CORE_DATAPATH_n_39;
  wire AES_CORE_DATAPATH_n_406;
  wire AES_CORE_DATAPATH_n_407;
  wire AES_CORE_DATAPATH_n_408;
  wire AES_CORE_DATAPATH_n_409;
  wire AES_CORE_DATAPATH_n_410;
  wire AES_CORE_DATAPATH_n_411;
  wire AES_CORE_DATAPATH_n_412;
  wire AES_CORE_DATAPATH_n_413;
  wire AES_CORE_DATAPATH_n_414;
  wire AES_CORE_DATAPATH_n_415;
  wire AES_CORE_DATAPATH_n_416;
  wire AES_CORE_DATAPATH_n_417;
  wire AES_CORE_DATAPATH_n_418;
  wire AES_CORE_DATAPATH_n_419;
  wire AES_CORE_DATAPATH_n_420;
  wire AES_CORE_DATAPATH_n_421;
  wire AES_CORE_DATAPATH_n_450;
  wire AES_CORE_DATAPATH_n_451;
  wire AES_CORE_DATAPATH_n_452;
  wire AES_CORE_DATAPATH_n_453;
  wire AES_CORE_DATAPATH_n_454;
  wire AES_CORE_DATAPATH_n_455;
  wire AES_CORE_DATAPATH_n_456;
  wire AES_CORE_DATAPATH_n_457;
  wire AES_CORE_DATAPATH_n_458;
  wire AES_CORE_DATAPATH_n_459;
  wire AES_CORE_DATAPATH_n_460;
  wire AES_CORE_DATAPATH_n_461;
  wire AES_CORE_DATAPATH_n_462;
  wire AES_CORE_DATAPATH_n_463;
  wire AES_CORE_DATAPATH_n_464;
  wire AES_CORE_DATAPATH_n_465;
  wire AES_CORE_DATAPATH_n_466;
  wire AES_CORE_DATAPATH_n_467;
  wire AES_CORE_DATAPATH_n_468;
  wire AES_CORE_DATAPATH_n_469;
  wire AES_CORE_DATAPATH_n_470;
  wire AES_CORE_DATAPATH_n_535;
  wire AES_CORE_DATAPATH_n_536;
  wire AES_CORE_DATAPATH_n_537;
  wire AES_CORE_DATAPATH_n_538;
  wire AES_CORE_DATAPATH_n_539;
  wire AES_CORE_DATAPATH_n_540;
  wire AES_CORE_DATAPATH_n_541;
  wire AES_CORE_DATAPATH_n_542;
  wire AES_CORE_DATAPATH_n_543;
  wire AES_CORE_DATAPATH_n_544;
  wire AES_CORE_DATAPATH_n_545;
  wire AES_CORE_DATAPATH_n_546;
  wire AES_CORE_DATAPATH_n_547;
  wire AES_CORE_DATAPATH_n_548;
  wire AES_CORE_DATAPATH_n_549;
  wire AES_CORE_DATAPATH_n_550;
  wire AES_CORE_DATAPATH_n_551;
  wire AES_CORE_DATAPATH_n_552;
  wire AES_CORE_DATAPATH_n_553;
  wire AES_CORE_DATAPATH_n_554;
  wire AES_CORE_DATAPATH_n_555;
  wire AES_CORE_DATAPATH_n_556;
  wire AES_CORE_DATAPATH_n_557;
  wire AES_CORE_DATAPATH_n_558;
  wire AES_CORE_DATAPATH_n_559;
  wire AES_CORE_DATAPATH_n_560;
  wire AES_CORE_DATAPATH_n_561;
  wire AES_CORE_DATAPATH_n_562;
  wire AES_CORE_DATAPATH_n_563;
  wire AES_CORE_DATAPATH_n_564;
  wire AES_CORE_DATAPATH_n_62;
  wire AES_CORE_DATAPATH_n_631;
  wire AES_CORE_DATAPATH_n_664;
  wire AES_CORE_DATAPATH_n_665;
  wire AES_CORE_DATAPATH_n_666;
  wire AES_CORE_DATAPATH_n_667;
  wire AES_CORE_DATAPATH_n_668;
  wire AES_CORE_DATAPATH_n_669;
  wire AES_CORE_DATAPATH_n_670;
  wire AES_CORE_DATAPATH_n_671;
  wire AES_CORE_DATAPATH_n_672;
  wire AES_CORE_DATAPATH_n_673;
  wire AES_CORE_DATAPATH_n_674;
  wire AES_CORE_DATAPATH_n_675;
  wire AES_CORE_DATAPATH_n_676;
  wire AES_CORE_DATAPATH_n_677;
  wire AES_CORE_DATAPATH_n_678;
  wire AES_CORE_DATAPATH_n_679;
  wire AES_CORE_DATAPATH_n_680;
  wire AES_CORE_DATAPATH_n_681;
  wire AES_CORE_DATAPATH_n_682;
  wire AES_CORE_DATAPATH_n_683;
  wire AES_CORE_DATAPATH_n_684;
  wire AES_CORE_DATAPATH_n_685;
  wire AES_CORE_DATAPATH_n_686;
  wire AES_CORE_DATAPATH_n_687;
  wire AES_CORE_DATAPATH_n_688;
  wire AES_CORE_DATAPATH_n_689;
  wire AES_CORE_DATAPATH_n_690;
  wire AES_CORE_DATAPATH_n_691;
  wire AES_CORE_DATAPATH_n_692;
  wire AES_CORE_DATAPATH_n_693;
  wire AES_CORE_DATAPATH_n_694;
  wire AES_CORE_DATAPATH_n_695;
  wire AES_CORE_DATAPATH_n_696;
  wire AES_CORE_DATAPATH_n_697;
  wire AES_CORE_DATAPATH_n_698;
  wire AES_CORE_DATAPATH_n_699;
  wire AES_CORE_DATAPATH_n_700;
  wire AES_CORE_DATAPATH_n_701;
  wire AES_CORE_DATAPATH_n_702;
  wire AES_CORE_DATAPATH_n_703;
  wire AES_CORE_DATAPATH_n_704;
  wire AES_CORE_DATAPATH_n_705;
  wire AES_CORE_DATAPATH_n_706;
  wire AES_CORE_DATAPATH_n_707;
  wire AES_CORE_DATAPATH_n_708;
  wire AES_CORE_DATAPATH_n_709;
  wire AES_CORE_DATAPATH_n_710;
  wire AES_CORE_DATAPATH_n_711;
  wire AES_CORE_DATAPATH_n_712;
  wire AES_CORE_DATAPATH_n_713;
  wire AES_CORE_DATAPATH_n_714;
  wire AES_CORE_DATAPATH_n_715;
  wire AES_CORE_DATAPATH_n_716;
  wire AES_CORE_DATAPATH_n_717;
  wire AES_CORE_DATAPATH_n_718;
  wire AES_CORE_DATAPATH_n_719;
  wire AES_CORE_DATAPATH_n_720;
  wire AES_CORE_DATAPATH_n_93;
  wire \CD[0].col[3][0]_i_2 ;
  wire \CD[0].col[3][0]_i_2_0 ;
  wire \CD[0].col[3][0]_i_4 ;
  wire \CD[0].col[3][10]_i_12 ;
  wire \CD[0].col[3][10]_i_6 ;
  wire \CD[0].col[3][31]_i_22 ;
  wire \CD[0].col[3][5]_i_2 ;
  wire [31:0]\CD[0].col_reg[3]_8 ;
  wire [31:0]\CD[2].col_reg[1][31] ;
  wire [1:0]\CD[3].col_reg[0][31] ;
  wire \CD[3].col_reg[0][31]_0 ;
  wire [31:0]\CD[3].col_reg[0]_9 ;
  wire [7:0]D;
  wire [0:0]E;
  wire \FSM_sequential_state_reg[0] ;
  wire \FSM_sequential_state_reg[0]_0 ;
  wire \FSM_sequential_state_reg[0]_1 ;
  wire \FSM_sequential_state_reg[0]_2 ;
  wire \FSM_sequential_state_reg[0]_3 ;
  wire [0:0]\FSM_sequential_state_reg[1] ;
  wire \FSM_sequential_state_reg[2] ;
  wire \FSM_sequential_state_reg[2]_0 ;
  wire [0:0]\FSM_sequential_state_reg[2]_1 ;
  wire \FSM_sequential_state_reg[2]_2 ;
  wire \FSM_sequential_state_reg[2]_3 ;
  wire \FSM_sequential_state_reg[3] ;
  wire \FSM_sequential_state_reg[3]_0 ;
  wire \FSM_sequential_state_reg[3]_1 ;
  wire \FSM_sequential_state_reg[3]_2 ;
  wire \FSM_sequential_state_reg[3]_3 ;
  wire \FSM_sequential_state_reg[3]_4 ;
  wire [31:0]\IV_BKP_REGISTERS[0].bkp_1_reg[0][31] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][0] ;
  wire [0:0]\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ;
  wire [7:0]\IV_BKP_REGISTERS[0].bkp_reg[0][15] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][16] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][17] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][18] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][19] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][1] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][20] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][21] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][22] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][23] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][24] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][25] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][26] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][27] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][28] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][29] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][2] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][30] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][31] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][3] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][4] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][5] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][6] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][7] ;
  wire [31:0]\IV_BKP_REGISTERS[0].bkp_reg[0]_17 ;
  wire [31:0]\IV_BKP_REGISTERS[0].iv_reg[0]_7 ;
  wire [31:0]\IV_BKP_REGISTERS[1].bkp_1_reg[1][31] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][0] ;
  wire [0:0]\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][10] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][11] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][12] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][13] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][14] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][15] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][16] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][17] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][18] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][19] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][1] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][20] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][21] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][22] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][23] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][2] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][31] ;
  wire [7:0]\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][3] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][4] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][5] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][6] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][7] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][8] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][9] ;
  wire [31:0]\IV_BKP_REGISTERS[1].bkp_reg[1]_15 ;
  wire [31:0]\IV_BKP_REGISTERS[1].iv_reg[1]_6 ;
  wire [31:0]\IV_BKP_REGISTERS[2].bkp_1_reg[2][31] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][0] ;
  wire [0:0]\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][10] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][11] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][12] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][13] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][14] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][15] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][16] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][17] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][18] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][19] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][1] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][20] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][21] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][22] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][23] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][2] ;
  wire [7:0]\IV_BKP_REGISTERS[2].bkp_reg[2][31] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][3] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][4] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][5] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][6] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][7] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][8] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][9] ;
  wire [31:0]\IV_BKP_REGISTERS[2].iv_reg[2]_5 ;
  wire [31:0]\IV_BKP_REGISTERS[3].bkp_1_reg[3][31] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][0] ;
  wire [0:0]\IV_BKP_REGISTERS[3].bkp_reg[3][0]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][16] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][17] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][18] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][19] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][1] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][20] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][21] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][22] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][23] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][24] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][25] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][26] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][27] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][28] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][29] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][2] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][30] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][31] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][3] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][4] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][5] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][6] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][7] ;
  wire [0:0]\IV_BKP_REGISTERS[3].iv_reg[3][0] ;
  wire [31:0]\IV_BKP_REGISTERS[3].iv_reg[3]_4 ;
  wire [27:26]\KEY_EXPANDER/g_func ;
  wire [0:0]\KR[1].key_host_reg[2][0] ;
  wire [5:0]\KR[1].key_reg[2][12] ;
  wire [0:0]\KR[2].key_host_reg[1][0] ;
  wire [31:0]\KR[2].key_host_reg[1]_2 ;
  wire [0:0]\KR[3].key_host_reg[0][0] ;
  wire \KR[3].key_reg[0][31] ;
  wire [3:0]Q;
  wire \SBOX/SBOX[0]/isomorphism_inv_return033_out ;
  wire \SBOX/SBOX[0]/isomorphism_inv_return03_out ;
  wire \SBOX/SBOX[0]/isomorphism_inv_return05_out ;
  wire \SBOX/SBOX[0]/isomorphism_return114_out ;
  wire \SBOX/SBOX[0]/isomorphism_return179_out ;
  wire \SBOX/SBOX[0]/p_16_in ;
  wire \SBOX/SBOX[0]/p_86_in ;
  wire \SBOX/SBOX[0]/p_93_in ;
  wire \SBOX/SBOX[1]/isomorphism_inv_return033_out ;
  wire \SBOX/SBOX[1]/isomorphism_inv_return03_out ;
  wire \SBOX/SBOX[1]/isomorphism_inv_return05_out ;
  wire \SBOX/SBOX[1]/isomorphism_return114_out ;
  wire \SBOX/SBOX[1]/isomorphism_return179_out ;
  wire \SBOX/SBOX[1]/p_16_in ;
  wire \SBOX/SBOX[1]/p_86_in ;
  wire \SBOX/SBOX[1]/p_93_in ;
  wire \SBOX/SBOX[2]/isomorphism_inv_return033_out ;
  wire \SBOX/SBOX[2]/isomorphism_inv_return03_out ;
  wire \SBOX/SBOX[2]/isomorphism_inv_return05_out ;
  wire \SBOX/SBOX[2]/isomorphism_return114_out ;
  wire \SBOX/SBOX[2]/isomorphism_return179_out ;
  wire \SBOX/SBOX[2]/p_16_in ;
  wire \SBOX/SBOX[2]/p_86_in ;
  wire \SBOX/SBOX[2]/p_93_in ;
  wire \SBOX/SBOX[3]/isomorphism_return114_out ;
  wire \SBOX/SBOX[3]/isomorphism_return179_out ;
  wire [23:0]add_rk_out;
  wire add_rk_sel;
  wire [2:0]\aes_cr_reg[2] ;
  wire \aes_cr_reg[4] ;
  wire \aes_cr_reg[5] ;
  wire \aes_cr_reg[5]_0 ;
  wire [31:0]bus_swap;
  wire bypass_key_en;
  wire bypass_rk;
  wire ccf;
  wire ccf_reg;
  wire ccf_reg_0;
  wire clk_i;
  wire [2:0]col_en_cnt_unit;
  wire \col_en_cnt_unit_pp1_reg[3] ;
  wire [3:0]\col_en_cnt_unit_pp2_reg[3] ;
  wire [3:0]col_en_host;
  wire [31:4]col_out;
  wire [1:0]col_sel;
  wire \col_sel_pp1_reg[1] ;
  wire [1:0]col_sel_pp2;
  wire [15:0]data_in;
  wire [31:0]enable_i;
  wire \enable_i[6]_0 ;
  wire enable_i_0_sn_1;
  wire enable_i_2_sn_1;
  wire enable_i_3_sn_1;
  wire enable_i_6_sn_1;
  wire enc_dec;
  wire enc_dec_sbox;
  wire first_block;
  wire [27:0]info_o;
  wire \info_o[0]_0 ;
  wire [6:0]\info_o[0]_1 ;
  wire \info_o[28]_INST_0_i_15 ;
  wire \info_o[28]_INST_0_i_15_0 ;
  wire \info_o[31] ;
  wire \info_o[31]_0 ;
  wire \info_o[31]_INST_0_i_12 ;
  wire info_o_0_sn_1;
  wire info_o_10_sn_1;
  wire info_o_11_sn_1;
  wire info_o_12_sn_1;
  wire info_o_4_sn_1;
  wire info_o_6_sn_1;
  wire info_o_9_sn_1;
  wire [2:0]iv_en;
  wire iv_mux_out13_out;
  wire iv_mux_out16_out;
  wire key_derivation_en;
  wire [3:0]key_en;
  wire [3:0]key_en_cnt_unit;
  wire [3:0]key_en_pp1;
  wire \key_en_pp1_reg[3] ;
  wire [127:0]key_in;
  wire [31:0]key_out;
  wire [1:1]key_out_sel_pp1;
  wire [1:1]key_out_sel_pp2;
  wire key_sel;
  wire key_sel_mux;
  wire key_sel_pp1;
  wire [0:0]key_sel_rd;
  wire last_round;
  wire [15:0]last_round_pp2_reg;
  wire [31:0]p_0_in1_in;
  wire p_12_out;
  wire p_16_out;
  wire p_1_in;
  wire p_1_in2_in;
  wire p_1_in5_in;
  wire p_20_out;
  wire [31:0]p_2_in;
  wire p_8_out;
  wire [0:0]\rd_count_reg[2] ;
  wire \rd_count_reg[3] ;
  wire rk_out_sel;
  wire rk_out_sel_pp2;
  wire [1:0]rk_sel;
  wire [3:0]round;
  wire rst_i;
  wire [19:2]sbox_out_enc;
  wire \sbox_pp2_reg[31] ;
  wire [1:0]sbox_sel;
  wire [87:32]sr_input;

  assign enable_i_0_sp_1 = enable_i_0_sn_1;
  assign enable_i_2_sp_1 = enable_i_2_sn_1;
  assign enable_i_3_sp_1 = enable_i_3_sn_1;
  assign enable_i_6_sp_1 = enable_i_6_sn_1;
  assign info_o_0_sn_1 = info_o_0_sp_1;
  assign info_o_10_sn_1 = info_o_10_sp_1;
  assign info_o_11_sn_1 = info_o_11_sp_1;
  assign info_o_12_sn_1 = info_o_12_sp_1;
  assign info_o_4_sn_1 = info_o_4_sp_1;
  assign info_o_6_sn_1 = info_o_6_sp_1;
  assign info_o_9_sn_1 = info_o_9_sp_1;
  switch_elements_control_unit AES_CORE_CONTROL_UNIT
       (.\CD[0].col[3][0]_i_2_0 (AES_CORE_DATAPATH_n_664),
        .\CD[0].col[3][0]_i_4_0 (\CD[0].col[3][0]_i_4 ),
        .\CD[0].col[3][10]_i_12_0 (\CD[0].col[3][10]_i_12 ),
        .\CD[0].col[3][10]_i_3_0 (AES_CORE_DATAPATH_n_543),
        .\CD[0].col[3][10]_i_6_0 (\CD[0].col[3][10]_i_6 ),
        .\CD[0].col[3][11]_i_3_0 (AES_CORE_DATAPATH_n_544),
        .\CD[0].col[3][12]_i_3_0 (AES_CORE_DATAPATH_n_545),
        .\CD[0].col[3][13]_i_3_0 (AES_CORE_DATAPATH_n_546),
        .\CD[0].col[3][14]_i_3_0 (AES_CORE_DATAPATH_n_673),
        .\CD[0].col[3][15]_i_5_0 (AES_CORE_DATAPATH_n_674),
        .\CD[0].col[3][16]_i_2_0 (AES_CORE_DATAPATH_n_549),
        .\CD[0].col[3][16]_i_2_1 (AES_CORE_DATAPATH_n_675),
        .\CD[0].col[3][17]_i_2_0 (AES_CORE_DATAPATH_n_550),
        .\CD[0].col[3][17]_i_2_1 (AES_CORE_DATAPATH_n_676),
        .\CD[0].col[3][18]_i_2_0 (AES_CORE_DATAPATH_n_551),
        .\CD[0].col[3][18]_i_2_1 (AES_CORE_DATAPATH_n_677),
        .\CD[0].col[3][19]_i_2_0 (AES_CORE_DATAPATH_n_552),
        .\CD[0].col[3][19]_i_2_1 (AES_CORE_DATAPATH_n_678),
        .\CD[0].col[3][1]_i_2_0 (AES_CORE_DATAPATH_n_535),
        .\CD[0].col[3][1]_i_2_1 (AES_CORE_DATAPATH_n_665),
        .\CD[0].col[3][20]_i_2_0 (AES_CORE_DATAPATH_n_553),
        .\CD[0].col[3][20]_i_2_1 (AES_CORE_DATAPATH_n_679),
        .\CD[0].col[3][21]_i_2_0 (AES_CORE_DATAPATH_n_554),
        .\CD[0].col[3][21]_i_2_1 (AES_CORE_DATAPATH_n_680),
        .\CD[0].col[3][22]_i_2_0 (AES_CORE_DATAPATH_n_555),
        .\CD[0].col[3][22]_i_2_1 (AES_CORE_DATAPATH_n_681),
        .\CD[0].col[3][23]_i_2_0 (AES_CORE_DATAPATH_n_556),
        .\CD[0].col[3][23]_i_2_1 (AES_CORE_DATAPATH_n_682),
        .\CD[0].col[3][24]_i_2_0 (AES_CORE_DATAPATH_n_683),
        .\CD[0].col[3][25]_i_2_0 (AES_CORE_DATAPATH_n_684),
        .\CD[0].col[3][26]_i_2_0 (AES_CORE_DATAPATH_n_685),
        .\CD[0].col[3][27]_i_2_0 (AES_CORE_DATAPATH_n_686),
        .\CD[0].col[3][28]_i_2_0 (AES_CORE_DATAPATH_n_561),
        .\CD[0].col[3][29]_i_2_0 (AES_CORE_DATAPATH_n_687),
        .\CD[0].col[3][2]_i_2_0 (AES_CORE_DATAPATH_n_536),
        .\CD[0].col[3][2]_i_2_1 (AES_CORE_DATAPATH_n_666),
        .\CD[0].col[3][30]_i_2_0 (AES_CORE_DATAPATH_n_688),
        .\CD[0].col[3][31]_i_10_0 (\IV_BKP_REGISTERS[0].bkp_reg[0]_17 ),
        .\CD[0].col[3][31]_i_13_0 (\IV_BKP_REGISTERS[1].iv_reg[1]_6 ),
        .\CD[0].col[3][31]_i_13_1 (\IV_BKP_REGISTERS[0].iv_reg[0]_7 ),
        .\CD[0].col[3][31]_i_22 (\CD[0].col[3][31]_i_22 ),
        .\CD[0].col[3][31]_i_5_0 (\IV_BKP_REGISTERS[1].bkp_reg[1]_15 ),
        .\CD[0].col[3][31]_i_5_1 (AES_CORE_DATAPATH_n_689),
        .\CD[0].col[3][31]_i_7_0 (col_sel_pp2),
        .\CD[0].col[3][3]_i_2_0 (AES_CORE_DATAPATH_n_537),
        .\CD[0].col[3][3]_i_2_1 (AES_CORE_DATAPATH_n_667),
        .\CD[0].col[3][4]_i_2_0 (AES_CORE_DATAPATH_n_538),
        .\CD[0].col[3][4]_i_2_1 (AES_CORE_DATAPATH_n_668),
        .\CD[0].col[3][5]_i_2_0 (AES_CORE_DATAPATH_n_421),
        .\CD[0].col[3][5]_i_2_1 (AES_CORE_DATAPATH_n_631),
        .\CD[0].col[3][5]_i_2_2 (\CD[0].col[3][5]_i_2 ),
        .\CD[0].col[3][6]_i_2_0 (AES_CORE_DATAPATH_n_539),
        .\CD[0].col[3][6]_i_2_1 (AES_CORE_DATAPATH_n_669),
        .\CD[0].col[3][7]_i_2_0 (AES_CORE_DATAPATH_n_540),
        .\CD[0].col[3][7]_i_2_1 (AES_CORE_DATAPATH_n_670),
        .\CD[0].col[3][8]_i_3_0 (AES_CORE_DATAPATH_n_671),
        .\CD[0].col[3][9]_i_3_0 (AES_CORE_DATAPATH_n_672),
        .\CD[0].col_reg[3][31] ({AES_CORE_CONTROL_UNIT_n_138,AES_CORE_CONTROL_UNIT_n_139,AES_CORE_CONTROL_UNIT_n_140,AES_CORE_CONTROL_UNIT_n_141,AES_CORE_CONTROL_UNIT_n_142,AES_CORE_CONTROL_UNIT_n_143,AES_CORE_CONTROL_UNIT_n_144,AES_CORE_CONTROL_UNIT_n_145,AES_CORE_CONTROL_UNIT_n_146,AES_CORE_CONTROL_UNIT_n_147,AES_CORE_CONTROL_UNIT_n_148,AES_CORE_CONTROL_UNIT_n_149,AES_CORE_CONTROL_UNIT_n_150,AES_CORE_CONTROL_UNIT_n_151,AES_CORE_CONTROL_UNIT_n_152,AES_CORE_CONTROL_UNIT_n_153,AES_CORE_CONTROL_UNIT_n_154,AES_CORE_CONTROL_UNIT_n_155,AES_CORE_CONTROL_UNIT_n_156,AES_CORE_CONTROL_UNIT_n_157,AES_CORE_CONTROL_UNIT_n_158,AES_CORE_CONTROL_UNIT_n_159,AES_CORE_CONTROL_UNIT_n_160,AES_CORE_CONTROL_UNIT_n_161}),
        .\CD[0].col_reg[3][31]_0 ({AES_CORE_CONTROL_UNIT_n_194,AES_CORE_CONTROL_UNIT_n_195,AES_CORE_CONTROL_UNIT_n_196,AES_CORE_CONTROL_UNIT_n_197,AES_CORE_CONTROL_UNIT_n_198,AES_CORE_CONTROL_UNIT_n_199,AES_CORE_CONTROL_UNIT_n_200,AES_CORE_CONTROL_UNIT_n_201,AES_CORE_CONTROL_UNIT_n_202,AES_CORE_CONTROL_UNIT_n_203,AES_CORE_CONTROL_UNIT_n_204,AES_CORE_CONTROL_UNIT_n_205,AES_CORE_CONTROL_UNIT_n_206,AES_CORE_CONTROL_UNIT_n_207,AES_CORE_CONTROL_UNIT_n_208,AES_CORE_CONTROL_UNIT_n_209,AES_CORE_CONTROL_UNIT_n_210,AES_CORE_CONTROL_UNIT_n_211,AES_CORE_CONTROL_UNIT_n_212,AES_CORE_CONTROL_UNIT_n_213,AES_CORE_CONTROL_UNIT_n_214,AES_CORE_CONTROL_UNIT_n_215,AES_CORE_CONTROL_UNIT_n_216,AES_CORE_CONTROL_UNIT_n_217,AES_CORE_CONTROL_UNIT_n_218,AES_CORE_CONTROL_UNIT_n_219,AES_CORE_CONTROL_UNIT_n_220,AES_CORE_CONTROL_UNIT_n_221,AES_CORE_CONTROL_UNIT_n_222,AES_CORE_CONTROL_UNIT_n_223,AES_CORE_CONTROL_UNIT_n_224,AES_CORE_CONTROL_UNIT_n_225}),
        .\CD[0].col_reg[3][31]_1 (\col_en_cnt_unit_pp2_reg[3] ),
        .\CD[1].col_reg[2][10] (last_round_pp2_reg[2]),
        .\CD[1].col_reg[2][10]_0 (AES_CORE_DATAPATH_n_458),
        .\CD[1].col_reg[2][10]_1 (AES_CORE_DATAPATH_n_148),
        .\CD[1].col_reg[2][11] (last_round_pp2_reg[3]),
        .\CD[1].col_reg[2][11]_0 (AES_CORE_DATAPATH_n_459),
        .\CD[1].col_reg[2][11]_1 (AES_CORE_DATAPATH_n_149),
        .\CD[1].col_reg[2][12] (last_round_pp2_reg[4]),
        .\CD[1].col_reg[2][12]_0 (AES_CORE_DATAPATH_n_460),
        .\CD[1].col_reg[2][12]_1 (AES_CORE_DATAPATH_n_150),
        .\CD[1].col_reg[2][13] (last_round_pp2_reg[5]),
        .\CD[1].col_reg[2][13]_0 (AES_CORE_DATAPATH_n_461),
        .\CD[1].col_reg[2][13]_1 (AES_CORE_DATAPATH_n_151),
        .\CD[1].col_reg[2][14] (last_round_pp2_reg[6]),
        .\CD[1].col_reg[2][14]_0 (AES_CORE_DATAPATH_n_153),
        .\CD[1].col_reg[2][14]_1 (AES_CORE_DATAPATH_n_152),
        .\CD[1].col_reg[2][15] (last_round_pp2_reg[7]),
        .\CD[1].col_reg[2][15]_0 (AES_CORE_DATAPATH_n_155),
        .\CD[1].col_reg[2][15]_1 (AES_CORE_DATAPATH_n_154),
        .\CD[1].col_reg[2][16] (AES_CORE_DATAPATH_n_462),
        .\CD[1].col_reg[2][16]_0 (AES_CORE_DATAPATH_n_156),
        .\CD[1].col_reg[2][17] (AES_CORE_DATAPATH_n_463),
        .\CD[1].col_reg[2][17]_0 (AES_CORE_DATAPATH_n_157),
        .\CD[1].col_reg[2][18] (AES_CORE_DATAPATH_n_464),
        .\CD[1].col_reg[2][18]_0 (AES_CORE_DATAPATH_n_158),
        .\CD[1].col_reg[2][19] (AES_CORE_DATAPATH_n_465),
        .\CD[1].col_reg[2][19]_0 (AES_CORE_DATAPATH_n_159),
        .\CD[1].col_reg[2][20] (AES_CORE_DATAPATH_n_466),
        .\CD[1].col_reg[2][20]_0 (AES_CORE_DATAPATH_n_160),
        .\CD[1].col_reg[2][21] (AES_CORE_DATAPATH_n_467),
        .\CD[1].col_reg[2][21]_0 (AES_CORE_DATAPATH_n_161),
        .\CD[1].col_reg[2][22] (AES_CORE_DATAPATH_n_468),
        .\CD[1].col_reg[2][22]_0 (AES_CORE_DATAPATH_n_162),
        .\CD[1].col_reg[2][23] ({AES_CORE_CONTROL_UNIT_n_90,AES_CORE_CONTROL_UNIT_n_91,AES_CORE_CONTROL_UNIT_n_92,AES_CORE_CONTROL_UNIT_n_93,AES_CORE_CONTROL_UNIT_n_94,AES_CORE_CONTROL_UNIT_n_95,AES_CORE_CONTROL_UNIT_n_96,AES_CORE_CONTROL_UNIT_n_97,AES_CORE_CONTROL_UNIT_n_98,AES_CORE_CONTROL_UNIT_n_99,AES_CORE_CONTROL_UNIT_n_100,AES_CORE_CONTROL_UNIT_n_101,AES_CORE_CONTROL_UNIT_n_102,AES_CORE_CONTROL_UNIT_n_103,AES_CORE_CONTROL_UNIT_n_104,AES_CORE_CONTROL_UNIT_n_105,AES_CORE_CONTROL_UNIT_n_106,AES_CORE_CONTROL_UNIT_n_107,AES_CORE_CONTROL_UNIT_n_108,AES_CORE_CONTROL_UNIT_n_109,AES_CORE_CONTROL_UNIT_n_110,AES_CORE_CONTROL_UNIT_n_111,AES_CORE_CONTROL_UNIT_n_112,AES_CORE_CONTROL_UNIT_n_113}),
        .\CD[1].col_reg[2][23]_0 (AES_CORE_DATAPATH_n_469),
        .\CD[1].col_reg[2][23]_1 (AES_CORE_DATAPATH_n_163),
        .\CD[1].col_reg[2][31] ({AES_CORE_CONTROL_UNIT_n_226,AES_CORE_CONTROL_UNIT_n_227,AES_CORE_CONTROL_UNIT_n_228,AES_CORE_CONTROL_UNIT_n_229,AES_CORE_CONTROL_UNIT_n_230,AES_CORE_CONTROL_UNIT_n_231,AES_CORE_CONTROL_UNIT_n_232,AES_CORE_CONTROL_UNIT_n_233,AES_CORE_CONTROL_UNIT_n_234,AES_CORE_CONTROL_UNIT_n_235,AES_CORE_CONTROL_UNIT_n_236,AES_CORE_CONTROL_UNIT_n_237,AES_CORE_CONTROL_UNIT_n_238,AES_CORE_CONTROL_UNIT_n_239,AES_CORE_CONTROL_UNIT_n_240,AES_CORE_CONTROL_UNIT_n_241,AES_CORE_CONTROL_UNIT_n_242,AES_CORE_CONTROL_UNIT_n_243,AES_CORE_CONTROL_UNIT_n_244,AES_CORE_CONTROL_UNIT_n_245,AES_CORE_CONTROL_UNIT_n_246,AES_CORE_CONTROL_UNIT_n_247,AES_CORE_CONTROL_UNIT_n_248,AES_CORE_CONTROL_UNIT_n_249,AES_CORE_CONTROL_UNIT_n_250,AES_CORE_CONTROL_UNIT_n_251,AES_CORE_CONTROL_UNIT_n_252,AES_CORE_CONTROL_UNIT_n_253,AES_CORE_CONTROL_UNIT_n_254,AES_CORE_CONTROL_UNIT_n_255,AES_CORE_CONTROL_UNIT_n_256,AES_CORE_CONTROL_UNIT_n_257}),
        .\CD[1].col_reg[2][31]_0 ({\CD[2].col_reg[1][31] [15:8],sr_input[55:48],\CD[2].col_reg[1][31] [7:0],sr_input[39:32]}),
        .\CD[1].col_reg[2][8] (last_round_pp2_reg[0]),
        .\CD[1].col_reg[2][8]_0 (AES_CORE_DATAPATH_n_145),
        .\CD[1].col_reg[2][8]_1 (AES_CORE_DATAPATH_n_144),
        .\CD[1].col_reg[2][9] (last_round_pp2_reg[1]),
        .\CD[1].col_reg[2][9]_0 (AES_CORE_DATAPATH_n_147),
        .\CD[1].col_reg[2][9]_1 (AES_CORE_DATAPATH_n_146),
        .\CD[2].col_reg[1][0] (AES_CORE_DATAPATH_n_450),
        .\CD[2].col_reg[1][0]_0 (AES_CORE_DATAPATH_n_93),
        .\CD[2].col_reg[1][1] (AES_CORE_DATAPATH_n_451),
        .\CD[2].col_reg[1][1]_0 (AES_CORE_DATAPATH_n_126),
        .\CD[2].col_reg[1][23] ({AES_CORE_CONTROL_UNIT_n_114,AES_CORE_CONTROL_UNIT_n_115,AES_CORE_CONTROL_UNIT_n_116,AES_CORE_CONTROL_UNIT_n_117,AES_CORE_CONTROL_UNIT_n_118,AES_CORE_CONTROL_UNIT_n_119,AES_CORE_CONTROL_UNIT_n_120,AES_CORE_CONTROL_UNIT_n_121,AES_CORE_CONTROL_UNIT_n_122,AES_CORE_CONTROL_UNIT_n_123,AES_CORE_CONTROL_UNIT_n_124,AES_CORE_CONTROL_UNIT_n_125,AES_CORE_CONTROL_UNIT_n_126,AES_CORE_CONTROL_UNIT_n_127,AES_CORE_CONTROL_UNIT_n_128,AES_CORE_CONTROL_UNIT_n_129,AES_CORE_CONTROL_UNIT_n_130,AES_CORE_CONTROL_UNIT_n_131,AES_CORE_CONTROL_UNIT_n_132,AES_CORE_CONTROL_UNIT_n_133,AES_CORE_CONTROL_UNIT_n_134,AES_CORE_CONTROL_UNIT_n_135,AES_CORE_CONTROL_UNIT_n_136,AES_CORE_CONTROL_UNIT_n_137}),
        .\CD[2].col_reg[1][24] (last_round_pp2_reg[8]),
        .\CD[2].col_reg[1][24]_0 (AES_CORE_DATAPATH_n_165),
        .\CD[2].col_reg[1][24]_1 (AES_CORE_DATAPATH_n_164),
        .\CD[2].col_reg[1][25] (last_round_pp2_reg[9]),
        .\CD[2].col_reg[1][25]_0 (AES_CORE_DATAPATH_n_167),
        .\CD[2].col_reg[1][25]_1 (AES_CORE_DATAPATH_n_166),
        .\CD[2].col_reg[1][26] (last_round_pp2_reg[10]),
        .\CD[2].col_reg[1][26]_0 (AES_CORE_DATAPATH_n_169),
        .\CD[2].col_reg[1][26]_1 (AES_CORE_DATAPATH_n_168),
        .\CD[2].col_reg[1][27] (last_round_pp2_reg[11]),
        .\CD[2].col_reg[1][27]_0 (AES_CORE_DATAPATH_n_171),
        .\CD[2].col_reg[1][27]_1 (AES_CORE_DATAPATH_n_170),
        .\CD[2].col_reg[1][28] (last_round_pp2_reg[12]),
        .\CD[2].col_reg[1][28]_0 (AES_CORE_DATAPATH_n_470),
        .\CD[2].col_reg[1][28]_1 (AES_CORE_DATAPATH_n_172),
        .\CD[2].col_reg[1][29] (last_round_pp2_reg[13]),
        .\CD[2].col_reg[1][29]_0 (AES_CORE_DATAPATH_n_174),
        .\CD[2].col_reg[1][29]_1 (AES_CORE_DATAPATH_n_173),
        .\CD[2].col_reg[1][2] (AES_CORE_DATAPATH_n_452),
        .\CD[2].col_reg[1][2]_0 (AES_CORE_DATAPATH_n_127),
        .\CD[2].col_reg[1][30] (last_round_pp2_reg[14]),
        .\CD[2].col_reg[1][30]_0 (AES_CORE_DATAPATH_n_176),
        .\CD[2].col_reg[1][30]_1 (AES_CORE_DATAPATH_n_175),
        .\CD[2].col_reg[1][31] ({AES_CORE_CONTROL_UNIT_n_258,AES_CORE_CONTROL_UNIT_n_259,AES_CORE_CONTROL_UNIT_n_260,AES_CORE_CONTROL_UNIT_n_261,AES_CORE_CONTROL_UNIT_n_262,AES_CORE_CONTROL_UNIT_n_263,AES_CORE_CONTROL_UNIT_n_264,AES_CORE_CONTROL_UNIT_n_265,AES_CORE_CONTROL_UNIT_n_266,AES_CORE_CONTROL_UNIT_n_267,AES_CORE_CONTROL_UNIT_n_268,AES_CORE_CONTROL_UNIT_n_269,AES_CORE_CONTROL_UNIT_n_270,AES_CORE_CONTROL_UNIT_n_271,AES_CORE_CONTROL_UNIT_n_272,AES_CORE_CONTROL_UNIT_n_273,AES_CORE_CONTROL_UNIT_n_274,AES_CORE_CONTROL_UNIT_n_275,AES_CORE_CONTROL_UNIT_n_276,AES_CORE_CONTROL_UNIT_n_277,AES_CORE_CONTROL_UNIT_n_278,AES_CORE_CONTROL_UNIT_n_279,AES_CORE_CONTROL_UNIT_n_280,AES_CORE_CONTROL_UNIT_n_281,AES_CORE_CONTROL_UNIT_n_282,AES_CORE_CONTROL_UNIT_n_283,AES_CORE_CONTROL_UNIT_n_284,AES_CORE_CONTROL_UNIT_n_285,AES_CORE_CONTROL_UNIT_n_286,AES_CORE_CONTROL_UNIT_n_287,AES_CORE_CONTROL_UNIT_n_288,AES_CORE_CONTROL_UNIT_n_289}),
        .\CD[2].col_reg[1][31]_0 ({\CD[2].col_reg[1][31] [31:24],sr_input[87:80],\CD[2].col_reg[1][31] [23:16],sr_input[71:64]}),
        .\CD[2].col_reg[1][31]_1 (\IV_BKP_REGISTERS[1].bkp_reg[1][31] ),
        .\CD[2].col_reg[1][31]_2 (last_round_pp2_reg[15]),
        .\CD[2].col_reg[1][31]_3 (AES_CORE_DATAPATH_n_178),
        .\CD[2].col_reg[1][31]_4 (AES_CORE_DATAPATH_n_177),
        .\CD[2].col_reg[1][3] (AES_CORE_DATAPATH_n_453),
        .\CD[2].col_reg[1][3]_0 (AES_CORE_DATAPATH_n_128),
        .\CD[2].col_reg[1][4] (AES_CORE_DATAPATH_n_454),
        .\CD[2].col_reg[1][4]_0 (AES_CORE_DATAPATH_n_129),
        .\CD[2].col_reg[1][5] (AES_CORE_DATAPATH_n_455),
        .\CD[2].col_reg[1][5]_0 (AES_CORE_DATAPATH_n_130),
        .\CD[2].col_reg[1][6] (AES_CORE_DATAPATH_n_456),
        .\CD[2].col_reg[1][6]_0 (AES_CORE_DATAPATH_n_131),
        .\CD[2].col_reg[1][7] (AES_CORE_DATAPATH_n_457),
        .\CD[2].col_reg[1][7]_0 (AES_CORE_DATAPATH_n_132),
        .\CD[3].col_reg[0][0] (AES_CORE_CONTROL_UNIT_n_339),
        .\CD[3].col_reg[0][10] (AES_CORE_CONTROL_UNIT_n_360),
        .\CD[3].col_reg[0][11] (AES_CORE_CONTROL_UNIT_n_358),
        .\CD[3].col_reg[0][12] (AES_CORE_CONTROL_UNIT_n_356),
        .\CD[3].col_reg[0][13] (AES_CORE_CONTROL_UNIT_n_352),
        .\CD[3].col_reg[0][14] (AES_CORE_CONTROL_UNIT_n_348),
        .\CD[3].col_reg[0][15] (AES_CORE_CONTROL_UNIT_n_344),
        .\CD[3].col_reg[0][16] (AES_CORE_CONTROL_UNIT_n_373),
        .\CD[3].col_reg[0][17] (AES_CORE_CONTROL_UNIT_n_372),
        .\CD[3].col_reg[0][18] (AES_CORE_CONTROL_UNIT_n_371),
        .\CD[3].col_reg[0][19] (AES_CORE_CONTROL_UNIT_n_370),
        .\CD[3].col_reg[0][1] (AES_CORE_CONTROL_UNIT_n_346),
        .\CD[3].col_reg[0][20] (AES_CORE_CONTROL_UNIT_n_369),
        .\CD[3].col_reg[0][21] (AES_CORE_CONTROL_UNIT_n_368),
        .\CD[3].col_reg[0][22] (AES_CORE_CONTROL_UNIT_n_367),
        .\CD[3].col_reg[0][23] (AES_CORE_CONTROL_UNIT_n_366),
        .\CD[3].col_reg[0][24] (AES_CORE_CONTROL_UNIT_n_365),
        .\CD[3].col_reg[0][25] (AES_CORE_CONTROL_UNIT_n_363),
        .\CD[3].col_reg[0][26] (AES_CORE_CONTROL_UNIT_n_361),
        .\CD[3].col_reg[0][27] (AES_CORE_CONTROL_UNIT_n_359),
        .\CD[3].col_reg[0][28] (AES_CORE_CONTROL_UNIT_n_357),
        .\CD[3].col_reg[0][29] (AES_CORE_CONTROL_UNIT_n_353),
        .\CD[3].col_reg[0][2] (AES_CORE_CONTROL_UNIT_n_350),
        .\CD[3].col_reg[0][30] (AES_CORE_CONTROL_UNIT_n_349),
        .\CD[3].col_reg[0][31] ({p_0_in1_in[31:16],p_0_in1_in[7:0]}),
        .\CD[3].col_reg[0][31]_0 (p_2_in),
        .\CD[3].col_reg[0][31]_1 (AES_CORE_CONTROL_UNIT_n_345),
        .\CD[3].col_reg[0][31]_2 (\CD[3].col_reg[0][31] ),
        .\CD[3].col_reg[0][31]_3 (\CD[3].col_reg[0][31]_0 ),
        .\CD[3].col_reg[0][3] (AES_CORE_CONTROL_UNIT_n_354),
        .\CD[3].col_reg[0][4] (AES_CORE_CONTROL_UNIT_n_355),
        .\CD[3].col_reg[0][5] (AES_CORE_CONTROL_UNIT_n_351),
        .\CD[3].col_reg[0][6] (AES_CORE_CONTROL_UNIT_n_347),
        .\CD[3].col_reg[0][7] (AES_CORE_CONTROL_UNIT_n_343),
        .\CD[3].col_reg[0][8] (AES_CORE_CONTROL_UNIT_n_364),
        .\CD[3].col_reg[0][9] (AES_CORE_CONTROL_UNIT_n_362),
        .D(col_sel),
        .E(p_1_in5_in),
        .\FSM_sequential_state_reg[0]_0 (\FSM_sequential_state_reg[0] ),
        .\FSM_sequential_state_reg[0]_1 (key_en_cnt_unit),
        .\FSM_sequential_state_reg[0]_2 (\FSM_sequential_state_reg[0]_0 ),
        .\FSM_sequential_state_reg[0]_3 (\FSM_sequential_state_reg[0]_1 ),
        .\FSM_sequential_state_reg[0]_4 (\FSM_sequential_state_reg[0]_2 ),
        .\FSM_sequential_state_reg[0]_5 (\FSM_sequential_state_reg[0]_3 ),
        .\FSM_sequential_state_reg[1]_0 (rk_sel),
        .\FSM_sequential_state_reg[1]_1 (\FSM_sequential_state_reg[1] ),
        .\FSM_sequential_state_reg[2]_0 (\FSM_sequential_state_reg[2] ),
        .\FSM_sequential_state_reg[2]_1 (\FSM_sequential_state_reg[2]_0 ),
        .\FSM_sequential_state_reg[2]_2 ({\FSM_sequential_state_reg[2]_1 ,col_en_cnt_unit}),
        .\FSM_sequential_state_reg[2]_3 (sbox_sel),
        .\FSM_sequential_state_reg[2]_4 (\FSM_sequential_state_reg[2]_2 ),
        .\FSM_sequential_state_reg[2]_5 (bypass_rk),
        .\FSM_sequential_state_reg[2]_6 (AES_CORE_CONTROL_UNIT_n_340),
        .\FSM_sequential_state_reg[2]_7 (\FSM_sequential_state_reg[2]_3 ),
        .\FSM_sequential_state_reg[3]_0 (\FSM_sequential_state_reg[3] ),
        .\FSM_sequential_state_reg[3]_1 (\FSM_sequential_state_reg[3]_0 ),
        .\FSM_sequential_state_reg[3]_10 (\FSM_sequential_state_reg[3]_3 ),
        .\FSM_sequential_state_reg[3]_11 (\FSM_sequential_state_reg[3]_4 ),
        .\FSM_sequential_state_reg[3]_2 (\FSM_sequential_state_reg[3]_1 ),
        .\FSM_sequential_state_reg[3]_3 (AES_CORE_CONTROL_UNIT_n_341),
        .\FSM_sequential_state_reg[3]_4 (AES_CORE_CONTROL_UNIT_n_342),
        .\FSM_sequential_state_reg[3]_5 (AES_CORE_CONTROL_UNIT_n_394),
        .\FSM_sequential_state_reg[3]_6 (AES_CORE_CONTROL_UNIT_n_395),
        .\FSM_sequential_state_reg[3]_7 (AES_CORE_CONTROL_UNIT_n_436),
        .\FSM_sequential_state_reg[3]_8 (AES_CORE_CONTROL_UNIT_n_437),
        .\FSM_sequential_state_reg[3]_9 (\FSM_sequential_state_reg[3]_2 ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][0] (\IV_BKP_REGISTERS[0].bkp_reg[0][0] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][16] (\IV_BKP_REGISTERS[0].bkp_reg[0][16] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][17] (\IV_BKP_REGISTERS[0].bkp_reg[0][17] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][18] (\IV_BKP_REGISTERS[0].bkp_reg[0][18] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][19] (\IV_BKP_REGISTERS[0].bkp_reg[0][19] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][1] (\IV_BKP_REGISTERS[0].bkp_reg[0][1] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][20] (\IV_BKP_REGISTERS[0].bkp_reg[0][20] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][21] (\IV_BKP_REGISTERS[0].bkp_reg[0][21] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][22] (\IV_BKP_REGISTERS[0].bkp_reg[0][22] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][23] (\IV_BKP_REGISTERS[0].bkp_reg[0][23] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][24] (\IV_BKP_REGISTERS[0].bkp_reg[0][24] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][25] (\IV_BKP_REGISTERS[0].bkp_reg[0][25] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][26] (\IV_BKP_REGISTERS[0].bkp_reg[0][26] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][27] (\IV_BKP_REGISTERS[0].bkp_reg[0][27] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][28] (\IV_BKP_REGISTERS[0].bkp_reg[0][28] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][29] (\IV_BKP_REGISTERS[0].bkp_reg[0][29] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][2] (\IV_BKP_REGISTERS[0].bkp_reg[0][2] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][30] (\IV_BKP_REGISTERS[0].bkp_reg[0][30] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][31] (\CD[0].col_reg[3]_8 ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 (\IV_BKP_REGISTERS[0].bkp_reg[0][31] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][3] (\IV_BKP_REGISTERS[0].bkp_reg[0][3] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][4] (\IV_BKP_REGISTERS[0].bkp_reg[0][4] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][5] (\IV_BKP_REGISTERS[0].bkp_reg[0][5] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][6] (\IV_BKP_REGISTERS[0].bkp_reg[0][6] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][7] (\IV_BKP_REGISTERS[0].bkp_reg[0][7] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][0] (\IV_BKP_REGISTERS[1].bkp_reg[1][0] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][10] (\IV_BKP_REGISTERS[1].bkp_reg[1][10] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][11] (\IV_BKP_REGISTERS[1].bkp_reg[1][11] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][12] (\IV_BKP_REGISTERS[1].bkp_reg[1][12] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][13] (\IV_BKP_REGISTERS[1].bkp_reg[1][13] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][14] (\IV_BKP_REGISTERS[1].bkp_reg[1][14] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][15] (\IV_BKP_REGISTERS[1].bkp_reg[1][15] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][16] (\IV_BKP_REGISTERS[1].bkp_reg[1][16] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][17] (\IV_BKP_REGISTERS[1].bkp_reg[1][17] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][18] (\IV_BKP_REGISTERS[1].bkp_reg[1][18] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][19] (\IV_BKP_REGISTERS[1].bkp_reg[1][19] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][1] (\IV_BKP_REGISTERS[1].bkp_reg[1][1] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][20] (\IV_BKP_REGISTERS[1].bkp_reg[1][20] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][21] (\IV_BKP_REGISTERS[1].bkp_reg[1][21] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][22] (\IV_BKP_REGISTERS[1].bkp_reg[1][22] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][23] (\IV_BKP_REGISTERS[1].bkp_reg[1][23] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][2] (\IV_BKP_REGISTERS[1].bkp_reg[1][2] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][3] (\IV_BKP_REGISTERS[1].bkp_reg[1][3] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][4] (\IV_BKP_REGISTERS[1].bkp_reg[1][4] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][5] (\IV_BKP_REGISTERS[1].bkp_reg[1][5] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][6] (\IV_BKP_REGISTERS[1].bkp_reg[1][6] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][7] (\IV_BKP_REGISTERS[1].bkp_reg[1][7] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][8] (\IV_BKP_REGISTERS[1].bkp_reg[1][8] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][9] (\IV_BKP_REGISTERS[1].bkp_reg[1][9] ),
        .\IV_BKP_REGISTERS[2].bkp[2][24]_i_2 (AES_CORE_DATAPATH_n_557),
        .\IV_BKP_REGISTERS[2].bkp[2][25]_i_2 (AES_CORE_DATAPATH_n_558),
        .\IV_BKP_REGISTERS[2].bkp[2][26]_i_2 (AES_CORE_DATAPATH_n_559),
        .\IV_BKP_REGISTERS[2].bkp[2][27]_i_2 (AES_CORE_DATAPATH_n_560),
        .\IV_BKP_REGISTERS[2].bkp[2][29]_i_2 (AES_CORE_DATAPATH_n_562),
        .\IV_BKP_REGISTERS[2].bkp[2][30]_i_2 (AES_CORE_DATAPATH_n_563),
        .\IV_BKP_REGISTERS[2].bkp[2][31]_i_2 (AES_CORE_DATAPATH_n_564),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][0] (\IV_BKP_REGISTERS[2].bkp_reg[2][0] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][10] (\IV_BKP_REGISTERS[2].bkp_reg[2][10] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][11] (\IV_BKP_REGISTERS[2].bkp_reg[2][11] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][12] (\IV_BKP_REGISTERS[2].bkp_reg[2][12] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][13] (\IV_BKP_REGISTERS[2].bkp_reg[2][13] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][14] (\IV_BKP_REGISTERS[2].bkp_reg[2][14] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][15] (\IV_BKP_REGISTERS[2].bkp_reg[2][15] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][16] (\IV_BKP_REGISTERS[2].bkp_reg[2][16] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][17] (\IV_BKP_REGISTERS[2].bkp_reg[2][17] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][18] (\IV_BKP_REGISTERS[2].bkp_reg[2][18] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][19] (\IV_BKP_REGISTERS[2].bkp_reg[2][19] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][1] (\IV_BKP_REGISTERS[2].bkp_reg[2][1] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][20] (\IV_BKP_REGISTERS[2].bkp_reg[2][20] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][21] (\IV_BKP_REGISTERS[2].bkp_reg[2][21] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][22] (\IV_BKP_REGISTERS[2].bkp_reg[2][22] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][23] (\IV_BKP_REGISTERS[2].bkp_reg[2][23] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][2] (\IV_BKP_REGISTERS[2].bkp_reg[2][2] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][3] (\IV_BKP_REGISTERS[2].bkp_reg[2][3] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][4] (\IV_BKP_REGISTERS[2].bkp_reg[2][4] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][5] (\IV_BKP_REGISTERS[2].bkp_reg[2][5] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][6] (\IV_BKP_REGISTERS[2].bkp_reg[2][6] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][7] (\IV_BKP_REGISTERS[2].bkp_reg[2][7] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][8] (\IV_BKP_REGISTERS[2].bkp_reg[2][8] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][9] (\IV_BKP_REGISTERS[2].bkp_reg[2][9] ),
        .\IV_BKP_REGISTERS[2].iv_reg[2][14] (AES_CORE_CONTROL_UNIT_n_298),
        .\IV_BKP_REGISTERS[2].iv_reg[2][15] (AES_CORE_CONTROL_UNIT_n_299),
        .\IV_BKP_REGISTERS[2].iv_reg[2][24] (AES_CORE_CONTROL_UNIT_n_300),
        .\IV_BKP_REGISTERS[2].iv_reg[2][25] (AES_CORE_CONTROL_UNIT_n_301),
        .\IV_BKP_REGISTERS[2].iv_reg[2][26] (AES_CORE_CONTROL_UNIT_n_302),
        .\IV_BKP_REGISTERS[2].iv_reg[2][27] (AES_CORE_CONTROL_UNIT_n_303),
        .\IV_BKP_REGISTERS[2].iv_reg[2][29] (AES_CORE_CONTROL_UNIT_n_304),
        .\IV_BKP_REGISTERS[2].iv_reg[2][30] (AES_CORE_CONTROL_UNIT_n_305),
        .\IV_BKP_REGISTERS[2].iv_reg[2][31] (AES_CORE_CONTROL_UNIT_n_306),
        .\IV_BKP_REGISTERS[2].iv_reg[2][8] (AES_CORE_CONTROL_UNIT_n_291),
        .\IV_BKP_REGISTERS[2].iv_reg[2][9] (AES_CORE_CONTROL_UNIT_n_292),
        .\IV_BKP_REGISTERS[3].bkp[3][14]_i_2 (AES_CORE_DATAPATH_n_547),
        .\IV_BKP_REGISTERS[3].bkp[3][15]_i_4 (AES_CORE_DATAPATH_n_548),
        .\IV_BKP_REGISTERS[3].bkp[3][8]_i_2 (AES_CORE_DATAPATH_n_541),
        .\IV_BKP_REGISTERS[3].bkp[3][9]_i_2 (AES_CORE_DATAPATH_n_542),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][0] (\IV_BKP_REGISTERS[3].bkp_reg[3][0] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][16] (\IV_BKP_REGISTERS[3].bkp_reg[3][16] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][17] (\IV_BKP_REGISTERS[3].bkp_reg[3][17] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][18] (\IV_BKP_REGISTERS[3].bkp_reg[3][18] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][19] (\IV_BKP_REGISTERS[3].bkp_reg[3][19] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][1] (\IV_BKP_REGISTERS[3].bkp_reg[3][1] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][20] (\IV_BKP_REGISTERS[3].bkp_reg[3][20] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][21] (\IV_BKP_REGISTERS[3].bkp_reg[3][21] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][22] (\IV_BKP_REGISTERS[3].bkp_reg[3][22] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][23] (\IV_BKP_REGISTERS[3].bkp_reg[3][23] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][24] (\IV_BKP_REGISTERS[3].bkp_reg[3][24] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][25] (\IV_BKP_REGISTERS[3].bkp_reg[3][25] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][26] (\IV_BKP_REGISTERS[3].bkp_reg[3][26] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][27] (\IV_BKP_REGISTERS[3].bkp_reg[3][27] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][28] (\IV_BKP_REGISTERS[3].bkp_reg[3][28] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][29] (\IV_BKP_REGISTERS[3].bkp_reg[3][29] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][2] (\IV_BKP_REGISTERS[3].bkp_reg[3][2] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][30] (\IV_BKP_REGISTERS[3].bkp_reg[3][30] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][31] (\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 (\CD[3].col_reg[0]_9 ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 (\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][3] (\IV_BKP_REGISTERS[3].bkp_reg[3][3] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][4] (\IV_BKP_REGISTERS[3].bkp_reg[3][4] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][5] (\IV_BKP_REGISTERS[3].bkp_reg[3][5] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][6] (\IV_BKP_REGISTERS[3].bkp_reg[3][6] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][7] (\IV_BKP_REGISTERS[3].bkp_reg[3][7] ),
        .\IV_BKP_REGISTERS[3].iv_reg[3][14] (AES_CORE_CONTROL_UNIT_n_380),
        .\IV_BKP_REGISTERS[3].iv_reg[3][15] (AES_CORE_CONTROL_UNIT_n_381),
        .\IV_BKP_REGISTERS[3].iv_reg[3][16] ({AES_CORE_DATAPATH_n_698,AES_CORE_DATAPATH_n_699,AES_CORE_DATAPATH_n_700,AES_CORE_DATAPATH_n_701,AES_CORE_DATAPATH_n_702,AES_CORE_DATAPATH_n_703,AES_CORE_DATAPATH_n_704,AES_CORE_DATAPATH_n_705}),
        .\IV_BKP_REGISTERS[3].iv_reg[3][24] (AES_CORE_CONTROL_UNIT_n_382),
        .\IV_BKP_REGISTERS[3].iv_reg[3][24]_0 ({AES_CORE_DATAPATH_n_706,AES_CORE_DATAPATH_n_707,AES_CORE_DATAPATH_n_708,AES_CORE_DATAPATH_n_709,AES_CORE_DATAPATH_n_710,AES_CORE_DATAPATH_n_711,AES_CORE_DATAPATH_n_712,AES_CORE_DATAPATH_n_713}),
        .\IV_BKP_REGISTERS[3].iv_reg[3][25] (AES_CORE_CONTROL_UNIT_n_383),
        .\IV_BKP_REGISTERS[3].iv_reg[3][26] (AES_CORE_CONTROL_UNIT_n_384),
        .\IV_BKP_REGISTERS[3].iv_reg[3][27] (AES_CORE_CONTROL_UNIT_n_385),
        .\IV_BKP_REGISTERS[3].iv_reg[3][29] (AES_CORE_CONTROL_UNIT_n_386),
        .\IV_BKP_REGISTERS[3].iv_reg[3][30] (AES_CORE_CONTROL_UNIT_n_387),
        .\IV_BKP_REGISTERS[3].iv_reg[3][31] (AES_CORE_CONTROL_UNIT_n_388),
        .\IV_BKP_REGISTERS[3].iv_reg[3][8] (AES_CORE_CONTROL_UNIT_n_378),
        .\IV_BKP_REGISTERS[3].iv_reg[3][8]_0 ({AES_CORE_DATAPATH_n_690,AES_CORE_DATAPATH_n_691,AES_CORE_DATAPATH_n_692,AES_CORE_DATAPATH_n_693,AES_CORE_DATAPATH_n_694,AES_CORE_DATAPATH_n_695,AES_CORE_DATAPATH_n_696,AES_CORE_DATAPATH_n_697}),
        .\IV_BKP_REGISTERS[3].iv_reg[3][9] (AES_CORE_CONTROL_UNIT_n_379),
        .\KR[0].key_reg[3][31] (key_en_pp1),
        .\KR[2].key_reg[1][24] (AES_CORE_DATAPATH_n_62),
        .\KR[2].key_reg[1][25] (AES_CORE_DATAPATH_n_39),
        .\KR[2].key_reg[1][28] (AES_CORE_DATAPATH_n_36),
        .\KR[2].key_reg[1][29] (AES_CORE_DATAPATH_n_38),
        .\KR[2].key_reg[1][30] (AES_CORE_DATAPATH_n_35),
        .\KR[2].key_reg[1][31] (\KR[2].key_host_reg[1]_2 ),
        .\KR[2].key_reg[1][31]_0 (AES_CORE_DATAPATH_n_37),
        .\KR[3].key_reg[0][31] ({AES_CORE_CONTROL_UNIT_n_307,AES_CORE_CONTROL_UNIT_n_308,AES_CORE_CONTROL_UNIT_n_309,AES_CORE_CONTROL_UNIT_n_310,AES_CORE_CONTROL_UNIT_n_311,AES_CORE_CONTROL_UNIT_n_312,AES_CORE_CONTROL_UNIT_n_313,AES_CORE_CONTROL_UNIT_n_314,AES_CORE_CONTROL_UNIT_n_315,AES_CORE_CONTROL_UNIT_n_316,AES_CORE_CONTROL_UNIT_n_317,AES_CORE_CONTROL_UNIT_n_318,AES_CORE_CONTROL_UNIT_n_319,AES_CORE_CONTROL_UNIT_n_320,AES_CORE_CONTROL_UNIT_n_321,AES_CORE_CONTROL_UNIT_n_322,AES_CORE_CONTROL_UNIT_n_323,AES_CORE_CONTROL_UNIT_n_324,AES_CORE_CONTROL_UNIT_n_325,AES_CORE_CONTROL_UNIT_n_326,AES_CORE_CONTROL_UNIT_n_327,AES_CORE_CONTROL_UNIT_n_328,AES_CORE_CONTROL_UNIT_n_329,AES_CORE_CONTROL_UNIT_n_330,AES_CORE_CONTROL_UNIT_n_331,AES_CORE_CONTROL_UNIT_n_332,AES_CORE_CONTROL_UNIT_n_333,AES_CORE_CONTROL_UNIT_n_334,AES_CORE_CONTROL_UNIT_n_335,AES_CORE_CONTROL_UNIT_n_336,AES_CORE_CONTROL_UNIT_n_337,AES_CORE_CONTROL_UNIT_n_338}),
        .\KR[3].key_reg[0][31]_0 (\KR[3].key_reg[0][31] ),
        .O({AES_CORE_DATAPATH_n_714,AES_CORE_DATAPATH_n_715,AES_CORE_DATAPATH_n_716,AES_CORE_DATAPATH_n_717,AES_CORE_DATAPATH_n_718,AES_CORE_DATAPATH_n_719,AES_CORE_DATAPATH_n_720}),
        .Q(Q),
        .add_rk_out({add_rk_out[23:16],add_rk_out[7:0]}),
        .add_rk_sel(add_rk_sel),
        .\aes_cr_reg[4] (\aes_cr_reg[4] ),
        .\aes_cr_reg[5] (\aes_cr_reg[5] ),
        .\aes_cr_reg[5]_0 (\aes_cr_reg[5]_0 ),
        .\aes_cr_reg[7] (AES_CORE_CONTROL_UNIT_n_28),
        .\base_new_pp_reg[7] (AES_CORE_DATAPATH_n_409),
        .\base_new_pp_reg[7]_0 (AES_CORE_DATAPATH_n_416),
        .\base_new_pp_reg[7]_1 (AES_CORE_DATAPATH_n_414),
        .\base_new_pp_reg[7]_10 (AES_CORE_DATAPATH_n_406),
        .\base_new_pp_reg[7]_2 (AES_CORE_DATAPATH_n_417),
        .\base_new_pp_reg[7]_3 (AES_CORE_DATAPATH_n_420),
        .\base_new_pp_reg[7]_4 (AES_CORE_DATAPATH_n_419),
        .\base_new_pp_reg[7]_5 (AES_CORE_DATAPATH_n_408),
        .\base_new_pp_reg[7]_6 (AES_CORE_DATAPATH_n_415),
        .\base_new_pp_reg[7]_7 (AES_CORE_DATAPATH_n_413),
        .\base_new_pp_reg[7]_8 (AES_CORE_DATAPATH_n_407),
        .\base_new_pp_reg[7]_9 (AES_CORE_DATAPATH_n_325),
        .bus_swap(bus_swap),
        .bypass_key_en(bypass_key_en),
        .ccf(ccf),
        .ccf_reg(ccf_reg),
        .ccf_reg_0(ccf_reg_0),
        .clk_i(clk_i),
        .\col_en_cnt_unit_pp1_reg[3] (\col_en_cnt_unit_pp1_reg[3] ),
        .\col_en_cnt_unit_pp2_reg[0] (AES_CORE_CONTROL_UNIT_n_392),
        .\col_en_cnt_unit_pp2_reg[1] (p_1_in),
        .\col_en_cnt_unit_pp2_reg[2] (p_1_in2_in),
        .\col_en_cnt_unit_pp2_reg[3] (iv_mux_out16_out),
        .col_en_host(col_en_host),
        .col_out({col_out[31:6],col_out[4]}),
        .\col_sel_pp1_reg[1] (\col_sel_pp1_reg[1] ),
        .data_in({data_in[12],data_in[5:2]}),
        .enable_i(enable_i),
        .\enable_i[31] ({AES_CORE_CONTROL_UNIT_n_403,AES_CORE_CONTROL_UNIT_n_404,AES_CORE_CONTROL_UNIT_n_405,AES_CORE_CONTROL_UNIT_n_406,AES_CORE_CONTROL_UNIT_n_407,AES_CORE_CONTROL_UNIT_n_408,AES_CORE_CONTROL_UNIT_n_409,AES_CORE_CONTROL_UNIT_n_410,AES_CORE_CONTROL_UNIT_n_411,AES_CORE_CONTROL_UNIT_n_412,AES_CORE_CONTROL_UNIT_n_413,AES_CORE_CONTROL_UNIT_n_414,AES_CORE_CONTROL_UNIT_n_415,AES_CORE_CONTROL_UNIT_n_416,AES_CORE_CONTROL_UNIT_n_417,AES_CORE_CONTROL_UNIT_n_418,AES_CORE_CONTROL_UNIT_n_419,AES_CORE_CONTROL_UNIT_n_420,AES_CORE_CONTROL_UNIT_n_421,AES_CORE_CONTROL_UNIT_n_422,AES_CORE_CONTROL_UNIT_n_423,AES_CORE_CONTROL_UNIT_n_424,AES_CORE_CONTROL_UNIT_n_425,AES_CORE_CONTROL_UNIT_n_426,AES_CORE_CONTROL_UNIT_n_427,AES_CORE_CONTROL_UNIT_n_428,AES_CORE_CONTROL_UNIT_n_429,AES_CORE_CONTROL_UNIT_n_430,AES_CORE_CONTROL_UNIT_n_431,AES_CORE_CONTROL_UNIT_n_432,AES_CORE_CONTROL_UNIT_n_433,AES_CORE_CONTROL_UNIT_n_434}),
        .enc_dec(enc_dec),
        .enc_dec_sbox(enc_dec_sbox),
        .first_block(first_block),
        .first_block_reg(AES_CORE_CONTROL_UNIT_n_374),
        .first_block_reg_0(AES_CORE_CONTROL_UNIT_n_377),
        .first_block_reg_1(AES_CORE_CONTROL_UNIT_n_438),
        .g_func(\KEY_EXPANDER/g_func ),
        .info_o(info_o),
        .\info_o[0]_0 (\info_o[0]_1 [6:2]),
        .\info_o[28]_INST_0_i_15 (\info_o[28]_INST_0_i_15 ),
        .\info_o[28]_INST_0_i_15_0 (\info_o[28]_INST_0_i_15_0 ),
        .\info_o[31] (\info_o[31] ),
        .\info_o[31]_0 (\info_o[31]_0 ),
        .\info_o[31]_1 (enable_i_0_sn_1),
        .\info_o[31]_2 (\IV_BKP_REGISTERS[2].iv_reg[2]_5 ),
        .\info_o[31]_3 ({\IV_BKP_REGISTERS[3].iv_reg[3]_4 [31:6],\IV_BKP_REGISTERS[3].iv_reg[3]_4 [4],\IV_BKP_REGISTERS[3].iv_reg[3]_4 [0]}),
        .\info_o[31]_INST_0_i_12_0 (\info_o[31]_INST_0_i_12 ),
        .\info_o[31]_INST_0_i_4 (key_out_sel_pp1),
        .\info_o[31]_INST_0_i_4_0 (\sbox_pp2_reg[31] ),
        .\info_o[31]_INST_0_i_4_1 (key_out_sel_pp2),
        .info_o_0_sp_1(AES_CORE_DATAPATH_n_2),
        .info_o_10_sp_1(info_o_10_sn_1),
        .info_o_11_sp_1(info_o_11_sn_1),
        .info_o_12_sp_1(info_o_12_sn_1),
        .info_o_4_sp_1(info_o_4_sn_1),
        .info_o_6_sp_1(info_o_6_sn_1),
        .info_o_9_sp_1(info_o_9_sn_1),
        .isomorphism_inv_return033_out(\SBOX/SBOX[2]/isomorphism_inv_return033_out ),
        .isomorphism_inv_return033_out_12(\SBOX/SBOX[0]/isomorphism_inv_return033_out ),
        .isomorphism_inv_return033_out_6(\SBOX/SBOX[1]/isomorphism_inv_return033_out ),
        .isomorphism_inv_return03_out(\SBOX/SBOX[2]/isomorphism_inv_return03_out ),
        .isomorphism_inv_return03_out_13(\SBOX/SBOX[0]/isomorphism_inv_return03_out ),
        .isomorphism_inv_return03_out_7(\SBOX/SBOX[1]/isomorphism_inv_return03_out ),
        .isomorphism_inv_return05_out(\SBOX/SBOX[2]/isomorphism_inv_return05_out ),
        .isomorphism_inv_return05_out_14(\SBOX/SBOX[0]/isomorphism_inv_return05_out ),
        .isomorphism_inv_return05_out_8(\SBOX/SBOX[1]/isomorphism_inv_return05_out ),
        .isomorphism_return114_out(\SBOX/SBOX[3]/isomorphism_return114_out ),
        .isomorphism_return114_out_1(\SBOX/SBOX[2]/isomorphism_return114_out ),
        .isomorphism_return114_out_3(\SBOX/SBOX[1]/isomorphism_return114_out ),
        .isomorphism_return114_out_5(\SBOX/SBOX[0]/isomorphism_return114_out ),
        .isomorphism_return179_out(\SBOX/SBOX[3]/isomorphism_return179_out ),
        .isomorphism_return179_out_0(\SBOX/SBOX[2]/isomorphism_return179_out ),
        .isomorphism_return179_out_2(\SBOX/SBOX[1]/isomorphism_return179_out ),
        .isomorphism_return179_out_4(\SBOX/SBOX[0]/isomorphism_return179_out ),
        .iv_mux_out13_out(iv_mux_out13_out),
        .key_en(key_en),
        .\key_en_pp1_reg[0] (p_8_out),
        .\key_en_pp1_reg[1] (p_12_out),
        .\key_en_pp1_reg[2] (p_16_out),
        .\key_en_pp1_reg[3] (p_20_out),
        .\key_en_pp1_reg[3]_0 (\key_en_pp1_reg[3] ),
        .key_in(key_in),
        .key_out({key_out[31:13],key_out[8:7],key_out[0]}),
        .\key_out_sel_pp1_reg[1] (AES_CORE_CONTROL_UNIT_n_402),
        .key_sel(key_sel),
        .key_sel_mux(key_sel_mux),
        .key_sel_pp1(key_sel_pp1),
        .last_round(last_round),
        .\out_gf_pp[1]_i_2 (AES_CORE_DATAPATH_n_412),
        .\out_gf_pp[1]_i_2__0 (AES_CORE_DATAPATH_n_418),
        .\out_gf_pp[1]_i_2__1 (AES_CORE_DATAPATH_n_411),
        .\out_gf_pp[1]_i_2__2 (AES_CORE_DATAPATH_n_410),
        .p_16_in(\SBOX/SBOX[2]/p_16_in ),
        .p_16_in_11(\SBOX/SBOX[1]/p_16_in ),
        .p_16_in_17(\SBOX/SBOX[0]/p_16_in ),
        .p_86_in(\SBOX/SBOX[2]/p_86_in ),
        .p_86_in_15(\SBOX/SBOX[0]/p_86_in ),
        .p_86_in_9(\SBOX/SBOX[1]/p_86_in ),
        .p_93_in(\SBOX/SBOX[2]/p_93_in ),
        .p_93_in_10(\SBOX/SBOX[1]/p_93_in ),
        .p_93_in_16(\SBOX/SBOX[0]/p_93_in ),
        .\rd_count_reg[3]_0 (\rd_count_reg[3] ),
        .\rd_count_reg[3]_1 ({round[3],\rd_count_reg[2] ,round[1:0]}),
        .rk_out_sel_pp2(rk_out_sel_pp2),
        .rst_i(rst_i),
        .sbox_out_enc({sbox_out_enc[19:18],sbox_out_enc[11:10],sbox_out_enc[3:2]}));
  switch_elements_datapath AES_CORE_DATAPATH
       (.\CD[0].col[3][0]_i_2 (\CD[0].col[3][0]_i_2 ),
        .\CD[0].col[3][0]_i_2_0 (\CD[0].col[3][0]_i_2_0 ),
        .\CD[0].col[3][0]_i_6_0 (AES_CORE_CONTROL_UNIT_n_339),
        .\CD[0].col[3][10]_i_8_0 (AES_CORE_CONTROL_UNIT_n_360),
        .\CD[0].col[3][12]_i_8_0 (AES_CORE_CONTROL_UNIT_n_356),
        .\CD[0].col[3][13]_i_8_0 (AES_CORE_CONTROL_UNIT_n_352),
        .\CD[0].col[3][15]_i_11_0 (AES_CORE_CONTROL_UNIT_n_344),
        .\CD[0].col[3][16]_i_6_0 (AES_CORE_CONTROL_UNIT_n_373),
        .\CD[0].col[3][17]_i_6_0 (AES_CORE_CONTROL_UNIT_n_372),
        .\CD[0].col[3][18]_i_6_0 (AES_CORE_CONTROL_UNIT_n_371),
        .\CD[0].col[3][1]_i_6_0 (AES_CORE_CONTROL_UNIT_n_346),
        .\CD[0].col[3][20]_i_6_0 (AES_CORE_CONTROL_UNIT_n_369),
        .\CD[0].col[3][21]_i_6_0 (AES_CORE_CONTROL_UNIT_n_368),
        .\CD[0].col[3][23]_i_7_0 (AES_CORE_CONTROL_UNIT_n_366),
        .\CD[0].col[3][24]_i_6_0 (AES_CORE_CONTROL_UNIT_n_365),
        .\CD[0].col[3][25]_i_6_0 (AES_CORE_CONTROL_UNIT_n_363),
        .\CD[0].col[3][26]_i_6_0 (AES_CORE_CONTROL_UNIT_n_361),
        .\CD[0].col[3][28]_i_6_0 (AES_CORE_CONTROL_UNIT_n_357),
        .\CD[0].col[3][29]_i_6_0 (AES_CORE_CONTROL_UNIT_n_353),
        .\CD[0].col[3][2]_i_6_0 (AES_CORE_CONTROL_UNIT_n_350),
        .\CD[0].col[3][31]_i_12_0 (AES_CORE_CONTROL_UNIT_n_345),
        .\CD[0].col[3][31]_i_5 (AES_CORE_CONTROL_UNIT_n_438),
        .\CD[0].col[3][4]_i_6_0 (AES_CORE_CONTROL_UNIT_n_355),
        .\CD[0].col[3][5]_i_6_0 (AES_CORE_CONTROL_UNIT_n_351),
        .\CD[0].col[3][5]_i_7 (iv_mux_out16_out),
        .\CD[0].col[3][7]_i_7_0 (AES_CORE_CONTROL_UNIT_n_343),
        .\CD[0].col[3][7]_i_9_0 (AES_CORE_CONTROL_UNIT_n_436),
        .\CD[0].col[3][7]_i_9_1 (AES_CORE_CONTROL_UNIT_n_437),
        .\CD[0].col[3][8]_i_8_0 (AES_CORE_CONTROL_UNIT_n_364),
        .\CD[0].col[3][9]_i_8_0 (AES_CORE_CONTROL_UNIT_n_362),
        .\CD[0].col[3][9]_i_8_1 (Q[3:2]),
        .\CD[0].col_reg[3][31]_0 (p_1_in5_in),
        .\CD[0].col_reg[3][31]_1 ({AES_CORE_CONTROL_UNIT_n_194,AES_CORE_CONTROL_UNIT_n_195,AES_CORE_CONTROL_UNIT_n_196,AES_CORE_CONTROL_UNIT_n_197,AES_CORE_CONTROL_UNIT_n_198,AES_CORE_CONTROL_UNIT_n_199,AES_CORE_CONTROL_UNIT_n_200,AES_CORE_CONTROL_UNIT_n_201,AES_CORE_CONTROL_UNIT_n_202,AES_CORE_CONTROL_UNIT_n_203,AES_CORE_CONTROL_UNIT_n_204,AES_CORE_CONTROL_UNIT_n_205,AES_CORE_CONTROL_UNIT_n_206,AES_CORE_CONTROL_UNIT_n_207,AES_CORE_CONTROL_UNIT_n_208,AES_CORE_CONTROL_UNIT_n_209,AES_CORE_CONTROL_UNIT_n_210,AES_CORE_CONTROL_UNIT_n_211,AES_CORE_CONTROL_UNIT_n_212,AES_CORE_CONTROL_UNIT_n_213,AES_CORE_CONTROL_UNIT_n_214,AES_CORE_CONTROL_UNIT_n_215,AES_CORE_CONTROL_UNIT_n_216,AES_CORE_CONTROL_UNIT_n_217,AES_CORE_CONTROL_UNIT_n_218,AES_CORE_CONTROL_UNIT_n_219,AES_CORE_CONTROL_UNIT_n_220,AES_CORE_CONTROL_UNIT_n_221,AES_CORE_CONTROL_UNIT_n_222,AES_CORE_CONTROL_UNIT_n_223,AES_CORE_CONTROL_UNIT_n_224,AES_CORE_CONTROL_UNIT_n_225}),
        .\CD[1].col_reg[2][31]_0 ({\CD[2].col_reg[1][31] [15:8],sr_input[55:48],\CD[2].col_reg[1][31] [7:0],sr_input[39:32]}),
        .\CD[1].col_reg[2][31]_1 (p_1_in2_in),
        .\CD[1].col_reg[2][31]_2 ({AES_CORE_CONTROL_UNIT_n_226,AES_CORE_CONTROL_UNIT_n_227,AES_CORE_CONTROL_UNIT_n_228,AES_CORE_CONTROL_UNIT_n_229,AES_CORE_CONTROL_UNIT_n_230,AES_CORE_CONTROL_UNIT_n_231,AES_CORE_CONTROL_UNIT_n_232,AES_CORE_CONTROL_UNIT_n_233,AES_CORE_CONTROL_UNIT_n_234,AES_CORE_CONTROL_UNIT_n_235,AES_CORE_CONTROL_UNIT_n_236,AES_CORE_CONTROL_UNIT_n_237,AES_CORE_CONTROL_UNIT_n_238,AES_CORE_CONTROL_UNIT_n_239,AES_CORE_CONTROL_UNIT_n_240,AES_CORE_CONTROL_UNIT_n_241,AES_CORE_CONTROL_UNIT_n_242,AES_CORE_CONTROL_UNIT_n_243,AES_CORE_CONTROL_UNIT_n_244,AES_CORE_CONTROL_UNIT_n_245,AES_CORE_CONTROL_UNIT_n_246,AES_CORE_CONTROL_UNIT_n_247,AES_CORE_CONTROL_UNIT_n_248,AES_CORE_CONTROL_UNIT_n_249,AES_CORE_CONTROL_UNIT_n_250,AES_CORE_CONTROL_UNIT_n_251,AES_CORE_CONTROL_UNIT_n_252,AES_CORE_CONTROL_UNIT_n_253,AES_CORE_CONTROL_UNIT_n_254,AES_CORE_CONTROL_UNIT_n_255,AES_CORE_CONTROL_UNIT_n_256,AES_CORE_CONTROL_UNIT_n_257}),
        .\CD[2].col_reg[1][0]_0 (AES_CORE_DATAPATH_n_325),
        .\CD[2].col_reg[1][13]_0 (AES_CORE_DATAPATH_n_411),
        .\CD[2].col_reg[1][14]_0 (AES_CORE_DATAPATH_n_408),
        .\CD[2].col_reg[1][16]_0 (AES_CORE_DATAPATH_n_420),
        .\CD[2].col_reg[1][17]_0 (AES_CORE_DATAPATH_n_419),
        .\CD[2].col_reg[1][1]_0 (AES_CORE_DATAPATH_n_406),
        .\CD[2].col_reg[1][21]_0 (AES_CORE_DATAPATH_n_418),
        .\CD[2].col_reg[1][22]_0 (AES_CORE_DATAPATH_n_417),
        .\CD[2].col_reg[1][24]_0 (AES_CORE_DATAPATH_n_416),
        .\CD[2].col_reg[1][25]_0 (AES_CORE_DATAPATH_n_414),
        .\CD[2].col_reg[1][29]_0 (AES_CORE_DATAPATH_n_412),
        .\CD[2].col_reg[1][30]_0 (AES_CORE_DATAPATH_n_409),
        .\CD[2].col_reg[1][31]_0 ({\CD[2].col_reg[1][31] [31:24],sr_input[87:80],\CD[2].col_reg[1][31] [23:16],sr_input[71:64]}),
        .\CD[2].col_reg[1][31]_1 (p_1_in),
        .\CD[2].col_reg[1][31]_2 ({AES_CORE_CONTROL_UNIT_n_258,AES_CORE_CONTROL_UNIT_n_259,AES_CORE_CONTROL_UNIT_n_260,AES_CORE_CONTROL_UNIT_n_261,AES_CORE_CONTROL_UNIT_n_262,AES_CORE_CONTROL_UNIT_n_263,AES_CORE_CONTROL_UNIT_n_264,AES_CORE_CONTROL_UNIT_n_265,AES_CORE_CONTROL_UNIT_n_266,AES_CORE_CONTROL_UNIT_n_267,AES_CORE_CONTROL_UNIT_n_268,AES_CORE_CONTROL_UNIT_n_269,AES_CORE_CONTROL_UNIT_n_270,AES_CORE_CONTROL_UNIT_n_271,AES_CORE_CONTROL_UNIT_n_272,AES_CORE_CONTROL_UNIT_n_273,AES_CORE_CONTROL_UNIT_n_274,AES_CORE_CONTROL_UNIT_n_275,AES_CORE_CONTROL_UNIT_n_276,AES_CORE_CONTROL_UNIT_n_277,AES_CORE_CONTROL_UNIT_n_278,AES_CORE_CONTROL_UNIT_n_279,AES_CORE_CONTROL_UNIT_n_280,AES_CORE_CONTROL_UNIT_n_281,AES_CORE_CONTROL_UNIT_n_282,AES_CORE_CONTROL_UNIT_n_283,AES_CORE_CONTROL_UNIT_n_284,AES_CORE_CONTROL_UNIT_n_285,AES_CORE_CONTROL_UNIT_n_286,AES_CORE_CONTROL_UNIT_n_287,AES_CORE_CONTROL_UNIT_n_288,AES_CORE_CONTROL_UNIT_n_289}),
        .\CD[2].col_reg[1][5]_0 (AES_CORE_DATAPATH_n_410),
        .\CD[2].col_reg[1][6]_0 (AES_CORE_DATAPATH_n_407),
        .\CD[2].col_reg[1][8]_0 (AES_CORE_DATAPATH_n_415),
        .\CD[2].col_reg[1][9]_0 (AES_CORE_DATAPATH_n_413),
        .\CD[3].col_reg[0][31]_0 (\CD[3].col_reg[0]_9 ),
        .\CD[3].col_reg[0][31]_1 (AES_CORE_CONTROL_UNIT_n_392),
        .\CD[3].col_reg[0][31]_2 (p_2_in),
        .D(sbox_sel),
        .E(AES_CORE_CONTROL_UNIT_n_394),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 (\IV_BKP_REGISTERS[0].bkp_1_reg[0][31] ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 (\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][14]_0 (AES_CORE_CONTROL_UNIT_n_298),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][14]_1 (AES_CORE_CONTROL_UNIT_n_380),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][15]_0 (AES_CORE_CONTROL_UNIT_n_299),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][15]_1 (AES_CORE_CONTROL_UNIT_n_381),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 (\IV_BKP_REGISTERS[0].bkp_reg[0]_17 ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 ({AES_CORE_CONTROL_UNIT_n_138,AES_CORE_CONTROL_UNIT_n_139,AES_CORE_CONTROL_UNIT_n_140,AES_CORE_CONTROL_UNIT_n_141,AES_CORE_CONTROL_UNIT_n_142,AES_CORE_CONTROL_UNIT_n_143,AES_CORE_CONTROL_UNIT_n_144,AES_CORE_CONTROL_UNIT_n_145,AES_CORE_CONTROL_UNIT_n_146,AES_CORE_CONTROL_UNIT_n_147,AES_CORE_CONTROL_UNIT_n_148,AES_CORE_CONTROL_UNIT_n_149,AES_CORE_CONTROL_UNIT_n_150,AES_CORE_CONTROL_UNIT_n_151,AES_CORE_CONTROL_UNIT_n_152,AES_CORE_CONTROL_UNIT_n_153,\IV_BKP_REGISTERS[0].bkp_reg[0][15] ,AES_CORE_CONTROL_UNIT_n_154,AES_CORE_CONTROL_UNIT_n_155,AES_CORE_CONTROL_UNIT_n_156,AES_CORE_CONTROL_UNIT_n_157,AES_CORE_CONTROL_UNIT_n_158,AES_CORE_CONTROL_UNIT_n_159,AES_CORE_CONTROL_UNIT_n_160,AES_CORE_CONTROL_UNIT_n_161}),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][8]_0 (AES_CORE_CONTROL_UNIT_n_291),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][8]_1 (AES_CORE_CONTROL_UNIT_n_378),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][9]_0 (AES_CORE_CONTROL_UNIT_n_292),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][9]_1 (AES_CORE_CONTROL_UNIT_n_379),
        .\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 (\IV_BKP_REGISTERS[0].iv_reg[0]_7 ),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 (\IV_BKP_REGISTERS[1].bkp_1_reg[1][31] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 (\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][24]_0 (AES_CORE_CONTROL_UNIT_n_300),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][24]_1 (AES_CORE_CONTROL_UNIT_n_382),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][25]_0 (AES_CORE_CONTROL_UNIT_n_301),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][25]_1 (AES_CORE_CONTROL_UNIT_n_383),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][26]_0 (AES_CORE_CONTROL_UNIT_n_302),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][26]_1 (AES_CORE_CONTROL_UNIT_n_384),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][27]_0 (AES_CORE_CONTROL_UNIT_n_303),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][27]_1 (AES_CORE_CONTROL_UNIT_n_385),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][29]_0 (AES_CORE_CONTROL_UNIT_n_304),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][29]_1 (AES_CORE_CONTROL_UNIT_n_386),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][30]_0 (AES_CORE_CONTROL_UNIT_n_305),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][30]_1 (AES_CORE_CONTROL_UNIT_n_387),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 (\IV_BKP_REGISTERS[1].bkp_reg[1]_15 ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 (\IV_BKP_REGISTERS[1].bkp_reg[1][31] ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][31]_2 (AES_CORE_CONTROL_UNIT_n_306),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][31]_3 (AES_CORE_CONTROL_UNIT_n_388),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 ({\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 ,AES_CORE_CONTROL_UNIT_n_114,AES_CORE_CONTROL_UNIT_n_115,AES_CORE_CONTROL_UNIT_n_116,AES_CORE_CONTROL_UNIT_n_117,AES_CORE_CONTROL_UNIT_n_118,AES_CORE_CONTROL_UNIT_n_119,AES_CORE_CONTROL_UNIT_n_120,AES_CORE_CONTROL_UNIT_n_121,AES_CORE_CONTROL_UNIT_n_122,AES_CORE_CONTROL_UNIT_n_123,AES_CORE_CONTROL_UNIT_n_124,AES_CORE_CONTROL_UNIT_n_125,AES_CORE_CONTROL_UNIT_n_126,AES_CORE_CONTROL_UNIT_n_127,AES_CORE_CONTROL_UNIT_n_128,AES_CORE_CONTROL_UNIT_n_129,AES_CORE_CONTROL_UNIT_n_130,AES_CORE_CONTROL_UNIT_n_131,AES_CORE_CONTROL_UNIT_n_132,AES_CORE_CONTROL_UNIT_n_133,AES_CORE_CONTROL_UNIT_n_134,AES_CORE_CONTROL_UNIT_n_135,AES_CORE_CONTROL_UNIT_n_136,AES_CORE_CONTROL_UNIT_n_137}),
        .\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 (\IV_BKP_REGISTERS[1].iv_reg[1]_6 ),
        .\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 (AES_CORE_CONTROL_UNIT_n_374),
        .\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 (AES_CORE_CONTROL_UNIT_n_377),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 (\IV_BKP_REGISTERS[2].bkp_1_reg[2][31] ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 (\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 ({\IV_BKP_REGISTERS[2].bkp_reg[2][31] ,AES_CORE_CONTROL_UNIT_n_90,AES_CORE_CONTROL_UNIT_n_91,AES_CORE_CONTROL_UNIT_n_92,AES_CORE_CONTROL_UNIT_n_93,AES_CORE_CONTROL_UNIT_n_94,AES_CORE_CONTROL_UNIT_n_95,AES_CORE_CONTROL_UNIT_n_96,AES_CORE_CONTROL_UNIT_n_97,AES_CORE_CONTROL_UNIT_n_98,AES_CORE_CONTROL_UNIT_n_99,AES_CORE_CONTROL_UNIT_n_100,AES_CORE_CONTROL_UNIT_n_101,AES_CORE_CONTROL_UNIT_n_102,AES_CORE_CONTROL_UNIT_n_103,AES_CORE_CONTROL_UNIT_n_104,AES_CORE_CONTROL_UNIT_n_105,AES_CORE_CONTROL_UNIT_n_106,AES_CORE_CONTROL_UNIT_n_107,AES_CORE_CONTROL_UNIT_n_108,AES_CORE_CONTROL_UNIT_n_109,AES_CORE_CONTROL_UNIT_n_110,AES_CORE_CONTROL_UNIT_n_111,AES_CORE_CONTROL_UNIT_n_112,AES_CORE_CONTROL_UNIT_n_113}),
        .\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 (\IV_BKP_REGISTERS[2].iv_reg[2]_5 ),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 (\IV_BKP_REGISTERS[3].bkp_1_reg[3][31] ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][0]_0 (AES_CORE_DATAPATH_n_450),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 (\IV_BKP_REGISTERS[3].bkp_reg[3][0]_0 ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][10]_0 (AES_CORE_DATAPATH_n_458),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][11]_0 (AES_CORE_DATAPATH_n_459),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][12]_0 (AES_CORE_DATAPATH_n_460),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][13]_0 (AES_CORE_DATAPATH_n_461),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][14]_0 (AES_CORE_DATAPATH_n_153),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][15]_0 (AES_CORE_DATAPATH_n_155),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][16]_0 (AES_CORE_DATAPATH_n_462),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][17]_0 (AES_CORE_DATAPATH_n_463),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][18]_0 (AES_CORE_DATAPATH_n_464),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][19]_0 (AES_CORE_DATAPATH_n_465),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][1]_0 (AES_CORE_DATAPATH_n_451),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][20]_0 (AES_CORE_DATAPATH_n_466),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][21]_0 (AES_CORE_DATAPATH_n_467),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][22]_0 (AES_CORE_DATAPATH_n_468),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][23]_0 (AES_CORE_DATAPATH_n_469),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][24]_0 (AES_CORE_DATAPATH_n_165),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][25]_0 (AES_CORE_DATAPATH_n_167),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][26]_0 (AES_CORE_DATAPATH_n_169),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][27]_0 (AES_CORE_DATAPATH_n_171),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][28]_0 (AES_CORE_DATAPATH_n_470),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][29]_0 (AES_CORE_DATAPATH_n_174),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][2]_0 (AES_CORE_DATAPATH_n_452),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][30]_0 (AES_CORE_DATAPATH_n_176),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 (AES_CORE_DATAPATH_n_178),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 ({p_0_in1_in[31:16],D,p_0_in1_in[7:0]}),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][3]_0 (AES_CORE_DATAPATH_n_453),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][4]_0 (AES_CORE_DATAPATH_n_454),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][5]_0 (AES_CORE_DATAPATH_n_455),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][6]_0 (AES_CORE_DATAPATH_n_456),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][7]_0 (AES_CORE_DATAPATH_n_457),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][8]_0 (AES_CORE_DATAPATH_n_145),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][9]_0 (AES_CORE_DATAPATH_n_147),
        .\IV_BKP_REGISTERS[3].iv_reg[3][0]_0 (AES_CORE_DATAPATH_n_664),
        .\IV_BKP_REGISTERS[3].iv_reg[3][0]_1 ({AES_CORE_DATAPATH_n_690,AES_CORE_DATAPATH_n_691,AES_CORE_DATAPATH_n_692,AES_CORE_DATAPATH_n_693,AES_CORE_DATAPATH_n_694,AES_CORE_DATAPATH_n_695,AES_CORE_DATAPATH_n_696,AES_CORE_DATAPATH_n_697}),
        .\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 (\IV_BKP_REGISTERS[3].iv_reg[3][0] ),
        .\IV_BKP_REGISTERS[3].iv_reg[3][10]_0 (AES_CORE_DATAPATH_n_543),
        .\IV_BKP_REGISTERS[3].iv_reg[3][11]_0 (AES_CORE_DATAPATH_n_544),
        .\IV_BKP_REGISTERS[3].iv_reg[3][12]_0 (AES_CORE_DATAPATH_n_545),
        .\IV_BKP_REGISTERS[3].iv_reg[3][13]_0 (AES_CORE_DATAPATH_n_546),
        .\IV_BKP_REGISTERS[3].iv_reg[3][14]_0 (AES_CORE_DATAPATH_n_547),
        .\IV_BKP_REGISTERS[3].iv_reg[3][14]_1 (AES_CORE_DATAPATH_n_673),
        .\IV_BKP_REGISTERS[3].iv_reg[3][15]_0 (AES_CORE_DATAPATH_n_548),
        .\IV_BKP_REGISTERS[3].iv_reg[3][15]_1 (AES_CORE_DATAPATH_n_674),
        .\IV_BKP_REGISTERS[3].iv_reg[3][16]_0 (AES_CORE_DATAPATH_n_549),
        .\IV_BKP_REGISTERS[3].iv_reg[3][16]_1 (AES_CORE_DATAPATH_n_675),
        .\IV_BKP_REGISTERS[3].iv_reg[3][16]_2 ({AES_CORE_DATAPATH_n_698,AES_CORE_DATAPATH_n_699,AES_CORE_DATAPATH_n_700,AES_CORE_DATAPATH_n_701,AES_CORE_DATAPATH_n_702,AES_CORE_DATAPATH_n_703,AES_CORE_DATAPATH_n_704,AES_CORE_DATAPATH_n_705}),
        .\IV_BKP_REGISTERS[3].iv_reg[3][17]_0 (AES_CORE_DATAPATH_n_550),
        .\IV_BKP_REGISTERS[3].iv_reg[3][17]_1 (AES_CORE_DATAPATH_n_676),
        .\IV_BKP_REGISTERS[3].iv_reg[3][18]_0 (AES_CORE_DATAPATH_n_551),
        .\IV_BKP_REGISTERS[3].iv_reg[3][18]_1 (AES_CORE_DATAPATH_n_677),
        .\IV_BKP_REGISTERS[3].iv_reg[3][19]_0 (AES_CORE_DATAPATH_n_552),
        .\IV_BKP_REGISTERS[3].iv_reg[3][19]_1 (AES_CORE_DATAPATH_n_678),
        .\IV_BKP_REGISTERS[3].iv_reg[3][1]_0 (AES_CORE_DATAPATH_n_535),
        .\IV_BKP_REGISTERS[3].iv_reg[3][1]_1 (AES_CORE_DATAPATH_n_665),
        .\IV_BKP_REGISTERS[3].iv_reg[3][20]_0 (AES_CORE_DATAPATH_n_553),
        .\IV_BKP_REGISTERS[3].iv_reg[3][20]_1 (AES_CORE_DATAPATH_n_679),
        .\IV_BKP_REGISTERS[3].iv_reg[3][21]_0 (AES_CORE_DATAPATH_n_554),
        .\IV_BKP_REGISTERS[3].iv_reg[3][21]_1 (AES_CORE_DATAPATH_n_680),
        .\IV_BKP_REGISTERS[3].iv_reg[3][22]_0 (AES_CORE_DATAPATH_n_555),
        .\IV_BKP_REGISTERS[3].iv_reg[3][22]_1 (AES_CORE_DATAPATH_n_681),
        .\IV_BKP_REGISTERS[3].iv_reg[3][23]_0 (AES_CORE_DATAPATH_n_556),
        .\IV_BKP_REGISTERS[3].iv_reg[3][23]_1 (AES_CORE_DATAPATH_n_682),
        .\IV_BKP_REGISTERS[3].iv_reg[3][24]_0 (AES_CORE_DATAPATH_n_557),
        .\IV_BKP_REGISTERS[3].iv_reg[3][24]_1 (AES_CORE_DATAPATH_n_683),
        .\IV_BKP_REGISTERS[3].iv_reg[3][24]_2 ({AES_CORE_DATAPATH_n_706,AES_CORE_DATAPATH_n_707,AES_CORE_DATAPATH_n_708,AES_CORE_DATAPATH_n_709,AES_CORE_DATAPATH_n_710,AES_CORE_DATAPATH_n_711,AES_CORE_DATAPATH_n_712,AES_CORE_DATAPATH_n_713}),
        .\IV_BKP_REGISTERS[3].iv_reg[3][25]_0 (AES_CORE_DATAPATH_n_558),
        .\IV_BKP_REGISTERS[3].iv_reg[3][25]_1 (AES_CORE_DATAPATH_n_684),
        .\IV_BKP_REGISTERS[3].iv_reg[3][26]_0 (AES_CORE_DATAPATH_n_559),
        .\IV_BKP_REGISTERS[3].iv_reg[3][26]_1 (AES_CORE_DATAPATH_n_685),
        .\IV_BKP_REGISTERS[3].iv_reg[3][27]_0 (AES_CORE_DATAPATH_n_560),
        .\IV_BKP_REGISTERS[3].iv_reg[3][27]_1 (AES_CORE_DATAPATH_n_686),
        .\IV_BKP_REGISTERS[3].iv_reg[3][28]_0 (AES_CORE_DATAPATH_n_561),
        .\IV_BKP_REGISTERS[3].iv_reg[3][29]_0 (AES_CORE_DATAPATH_n_562),
        .\IV_BKP_REGISTERS[3].iv_reg[3][29]_1 (AES_CORE_DATAPATH_n_687),
        .\IV_BKP_REGISTERS[3].iv_reg[3][2]_0 (AES_CORE_DATAPATH_n_536),
        .\IV_BKP_REGISTERS[3].iv_reg[3][2]_1 (AES_CORE_DATAPATH_n_666),
        .\IV_BKP_REGISTERS[3].iv_reg[3][30]_0 (AES_CORE_DATAPATH_n_563),
        .\IV_BKP_REGISTERS[3].iv_reg[3][30]_1 (AES_CORE_DATAPATH_n_688),
        .\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 ({\IV_BKP_REGISTERS[3].iv_reg[3]_4 [31:6],\IV_BKP_REGISTERS[3].iv_reg[3]_4 [4],\IV_BKP_REGISTERS[3].iv_reg[3]_4 [0]}),
        .\IV_BKP_REGISTERS[3].iv_reg[3][31]_1 (AES_CORE_DATAPATH_n_564),
        .\IV_BKP_REGISTERS[3].iv_reg[3][31]_2 (AES_CORE_DATAPATH_n_689),
        .\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 ({AES_CORE_CONTROL_UNIT_n_403,AES_CORE_CONTROL_UNIT_n_404,AES_CORE_CONTROL_UNIT_n_405,AES_CORE_CONTROL_UNIT_n_406,AES_CORE_CONTROL_UNIT_n_407,AES_CORE_CONTROL_UNIT_n_408,AES_CORE_CONTROL_UNIT_n_409,AES_CORE_CONTROL_UNIT_n_410,AES_CORE_CONTROL_UNIT_n_411,AES_CORE_CONTROL_UNIT_n_412,AES_CORE_CONTROL_UNIT_n_413,AES_CORE_CONTROL_UNIT_n_414,AES_CORE_CONTROL_UNIT_n_415,AES_CORE_CONTROL_UNIT_n_416,AES_CORE_CONTROL_UNIT_n_417,AES_CORE_CONTROL_UNIT_n_418,AES_CORE_CONTROL_UNIT_n_419,AES_CORE_CONTROL_UNIT_n_420,AES_CORE_CONTROL_UNIT_n_421,AES_CORE_CONTROL_UNIT_n_422,AES_CORE_CONTROL_UNIT_n_423,AES_CORE_CONTROL_UNIT_n_424,AES_CORE_CONTROL_UNIT_n_425,AES_CORE_CONTROL_UNIT_n_426,AES_CORE_CONTROL_UNIT_n_427,AES_CORE_CONTROL_UNIT_n_428,AES_CORE_CONTROL_UNIT_n_429,AES_CORE_CONTROL_UNIT_n_430,AES_CORE_CONTROL_UNIT_n_431,AES_CORE_CONTROL_UNIT_n_432,AES_CORE_CONTROL_UNIT_n_433,AES_CORE_CONTROL_UNIT_n_434}),
        .\IV_BKP_REGISTERS[3].iv_reg[3][3]_0 (AES_CORE_DATAPATH_n_537),
        .\IV_BKP_REGISTERS[3].iv_reg[3][3]_1 (AES_CORE_DATAPATH_n_667),
        .\IV_BKP_REGISTERS[3].iv_reg[3][4]_0 (AES_CORE_DATAPATH_n_538),
        .\IV_BKP_REGISTERS[3].iv_reg[3][4]_1 (AES_CORE_DATAPATH_n_668),
        .\IV_BKP_REGISTERS[3].iv_reg[3][5]_0 (AES_CORE_DATAPATH_n_421),
        .\IV_BKP_REGISTERS[3].iv_reg[3][5]_1 (AES_CORE_DATAPATH_n_631),
        .\IV_BKP_REGISTERS[3].iv_reg[3][6]_0 (AES_CORE_DATAPATH_n_539),
        .\IV_BKP_REGISTERS[3].iv_reg[3][6]_1 (AES_CORE_DATAPATH_n_669),
        .\IV_BKP_REGISTERS[3].iv_reg[3][7]_0 (AES_CORE_DATAPATH_n_540),
        .\IV_BKP_REGISTERS[3].iv_reg[3][7]_1 (AES_CORE_DATAPATH_n_670),
        .\IV_BKP_REGISTERS[3].iv_reg[3][8]_0 (AES_CORE_DATAPATH_n_541),
        .\IV_BKP_REGISTERS[3].iv_reg[3][8]_1 (AES_CORE_DATAPATH_n_671),
        .\IV_BKP_REGISTERS[3].iv_reg[3][9]_0 (AES_CORE_DATAPATH_n_542),
        .\IV_BKP_REGISTERS[3].iv_reg[3][9]_1 (AES_CORE_DATAPATH_n_672),
        .\KR[0].key_host_reg[3][0]_0 (E),
        .\KR[0].key_reg[3][31]_0 (p_20_out),
        .\KR[1].key_host_reg[2][0]_0 (\KR[1].key_host_reg[2][0] ),
        .\KR[1].key_reg[2][10]_0 (\KR[1].key_reg[2][12] [3]),
        .\KR[1].key_reg[2][11]_0 (\KR[1].key_reg[2][12] [4]),
        .\KR[1].key_reg[2][12]_0 (\KR[1].key_reg[2][12] [5]),
        .\KR[1].key_reg[2][31]_0 (p_16_out),
        .\KR[1].key_reg[2][4]_0 (\KR[1].key_reg[2][12] [0]),
        .\KR[1].key_reg[2][6]_0 (\KR[1].key_reg[2][12] [1]),
        .\KR[1].key_reg[2][9]_0 (\KR[1].key_reg[2][12] [2]),
        .\KR[2].key_host_reg[1][0]_0 (\KR[2].key_host_reg[1][0] ),
        .\KR[2].key_host_reg[1][31]_0 (\KR[2].key_host_reg[1]_2 ),
        .\KR[2].key_reg[1][31]_0 (p_12_out),
        .\KR[2].key_reg[1][31]_1 ({AES_CORE_CONTROL_UNIT_n_307,AES_CORE_CONTROL_UNIT_n_308,AES_CORE_CONTROL_UNIT_n_309,AES_CORE_CONTROL_UNIT_n_310,AES_CORE_CONTROL_UNIT_n_311,AES_CORE_CONTROL_UNIT_n_312,AES_CORE_CONTROL_UNIT_n_313,AES_CORE_CONTROL_UNIT_n_314,AES_CORE_CONTROL_UNIT_n_315,AES_CORE_CONTROL_UNIT_n_316,AES_CORE_CONTROL_UNIT_n_317,AES_CORE_CONTROL_UNIT_n_318,AES_CORE_CONTROL_UNIT_n_319,AES_CORE_CONTROL_UNIT_n_320,AES_CORE_CONTROL_UNIT_n_321,AES_CORE_CONTROL_UNIT_n_322,AES_CORE_CONTROL_UNIT_n_323,AES_CORE_CONTROL_UNIT_n_324,AES_CORE_CONTROL_UNIT_n_325,AES_CORE_CONTROL_UNIT_n_326,AES_CORE_CONTROL_UNIT_n_327,AES_CORE_CONTROL_UNIT_n_328,AES_CORE_CONTROL_UNIT_n_329,AES_CORE_CONTROL_UNIT_n_330,AES_CORE_CONTROL_UNIT_n_331,AES_CORE_CONTROL_UNIT_n_332,AES_CORE_CONTROL_UNIT_n_333,AES_CORE_CONTROL_UNIT_n_334,AES_CORE_CONTROL_UNIT_n_335,AES_CORE_CONTROL_UNIT_n_336,AES_CORE_CONTROL_UNIT_n_337,AES_CORE_CONTROL_UNIT_n_338}),
        .\KR[3].key_host_reg[0][0]_0 (\KR[3].key_host_reg[0][0] ),
        .\KR[3].key_reg[0][31]_0 (p_8_out),
        .O({AES_CORE_DATAPATH_n_714,AES_CORE_DATAPATH_n_715,AES_CORE_DATAPATH_n_716,AES_CORE_DATAPATH_n_717,AES_CORE_DATAPATH_n_718,AES_CORE_DATAPATH_n_719,AES_CORE_DATAPATH_n_720}),
        .Q(\CD[0].col_reg[3]_8 ),
        .add_rk_out({add_rk_out[23:16],add_rk_out[7:0]}),
        .add_rk_sel(add_rk_sel),
        .\aes_cr_reg[0] (AES_CORE_DATAPATH_n_2),
        .\aes_cr_reg[2] ({col_out[31:6],col_out[4]}),
        .\aes_cr_reg[2]_0 (\aes_cr_reg[2] ),
        .\base_new_pp_reg[3] (AES_CORE_CONTROL_UNIT_n_354),
        .\base_new_pp_reg[3]_0 (AES_CORE_CONTROL_UNIT_n_358),
        .\base_new_pp_reg[3]_1 (AES_CORE_CONTROL_UNIT_n_359),
        .\base_new_pp_reg[3]_2 (AES_CORE_CONTROL_UNIT_n_370),
        .\base_new_pp_reg[4] (AES_CORE_CONTROL_UNIT_n_342),
        .\base_new_pp_reg[4]_0 (AES_CORE_CONTROL_UNIT_n_347),
        .\base_new_pp_reg[4]_1 (AES_CORE_CONTROL_UNIT_n_348),
        .\base_new_pp_reg[4]_2 (AES_CORE_CONTROL_UNIT_n_349),
        .\base_new_pp_reg[4]_3 (AES_CORE_CONTROL_UNIT_n_367),
        .bus_swap(bus_swap),
        .bypass_key_en(bypass_key_en),
        .clk_i(clk_i),
        .\col_en_cnt_unit_pp1_reg[0]_0 (AES_CORE_CONTROL_UNIT_n_395),
        .\col_en_cnt_unit_pp1_reg[3]_0 ({\FSM_sequential_state_reg[2]_1 ,col_en_cnt_unit}),
        .\col_en_cnt_unit_pp2_reg[3]_0 (\col_en_cnt_unit_pp2_reg[3] ),
        .\col_sel_pp1_reg[1]_0 (col_sel),
        .\col_sel_pp2_reg[1]_0 (col_sel_pp2),
        .data_in({data_in[15:13],data_in[11:6],data_in[1:0]}),
        .enable_i(enable_i),
        .\enable_i[0]_0 (AES_CORE_DATAPATH_n_156),
        .\enable_i[2]_0 (AES_CORE_DATAPATH_n_158),
        .\enable_i[3]_0 (AES_CORE_DATAPATH_n_159),
        .\enable_i[6]_0 (\enable_i[6]_0 ),
        .\enable_i[6]_1 (AES_CORE_DATAPATH_n_162),
        .enable_i_0_sp_1(enable_i_0_sn_1),
        .enable_i_10_sp_1(AES_CORE_DATAPATH_n_168),
        .enable_i_11_sp_1(AES_CORE_DATAPATH_n_170),
        .enable_i_12_sp_1(AES_CORE_DATAPATH_n_172),
        .enable_i_13_sp_1(AES_CORE_DATAPATH_n_173),
        .enable_i_14_sp_1(AES_CORE_DATAPATH_n_175),
        .enable_i_15_sp_1(AES_CORE_DATAPATH_n_177),
        .enable_i_16_sp_1(AES_CORE_DATAPATH_n_93),
        .enable_i_17_sp_1(AES_CORE_DATAPATH_n_126),
        .enable_i_18_sp_1(AES_CORE_DATAPATH_n_127),
        .enable_i_19_sp_1(AES_CORE_DATAPATH_n_128),
        .enable_i_1_sp_1(AES_CORE_DATAPATH_n_157),
        .enable_i_20_sp_1(AES_CORE_DATAPATH_n_129),
        .enable_i_21_sp_1(AES_CORE_DATAPATH_n_130),
        .enable_i_22_sp_1(AES_CORE_DATAPATH_n_131),
        .enable_i_23_sp_1(AES_CORE_DATAPATH_n_132),
        .enable_i_24_sp_1(AES_CORE_DATAPATH_n_144),
        .enable_i_25_sp_1(AES_CORE_DATAPATH_n_146),
        .enable_i_26_sp_1(AES_CORE_DATAPATH_n_148),
        .enable_i_27_sp_1(AES_CORE_DATAPATH_n_149),
        .enable_i_28_sp_1(AES_CORE_DATAPATH_n_150),
        .enable_i_29_sp_1(AES_CORE_DATAPATH_n_151),
        .enable_i_2_sp_1(enable_i_2_sn_1),
        .enable_i_30_sp_1(AES_CORE_DATAPATH_n_152),
        .enable_i_31_sp_1(AES_CORE_DATAPATH_n_154),
        .enable_i_3_sp_1(enable_i_3_sn_1),
        .enable_i_4_sp_1(AES_CORE_DATAPATH_n_160),
        .enable_i_5_sp_1(AES_CORE_DATAPATH_n_161),
        .enable_i_6_sp_1(enable_i_6_sn_1),
        .enable_i_7_sp_1(AES_CORE_DATAPATH_n_163),
        .enable_i_8_sp_1(AES_CORE_DATAPATH_n_164),
        .enable_i_9_sp_1(AES_CORE_DATAPATH_n_166),
        .enc_dec_sbox(enc_dec_sbox),
        .g_func(\KEY_EXPANDER/g_func ),
        .\info_o[0] (info_o_0_sn_1),
        .\info_o[0]_0 (AES_CORE_CONTROL_UNIT_n_28),
        .\info_o[0]_1 (\FSM_sequential_state_reg[3]_2 ),
        .\info_o[0]_2 (\info_o[0]_0 ),
        .\info_o[1] (\info_o[0]_1 [1:0]),
        .\info_o[28]_INST_0_i_7 (AES_CORE_CONTROL_UNIT_n_341),
        .\info_o[28]_INST_0_i_7_0 (AES_CORE_CONTROL_UNIT_n_340),
        .isomorphism_inv_return033_out(\SBOX/SBOX[2]/isomorphism_inv_return033_out ),
        .isomorphism_inv_return033_out_3(\SBOX/SBOX[1]/isomorphism_inv_return033_out ),
        .isomorphism_inv_return033_out_9(\SBOX/SBOX[0]/isomorphism_inv_return033_out ),
        .isomorphism_inv_return03_out(\SBOX/SBOX[2]/isomorphism_inv_return03_out ),
        .isomorphism_inv_return03_out_1(\SBOX/SBOX[1]/isomorphism_inv_return03_out ),
        .isomorphism_inv_return03_out_7(\SBOX/SBOX[0]/isomorphism_inv_return03_out ),
        .isomorphism_inv_return05_out(\SBOX/SBOX[2]/isomorphism_inv_return05_out ),
        .isomorphism_inv_return05_out_10(\SBOX/SBOX[0]/isomorphism_inv_return05_out ),
        .isomorphism_inv_return05_out_4(\SBOX/SBOX[1]/isomorphism_inv_return05_out ),
        .isomorphism_return114_out(\SBOX/SBOX[3]/isomorphism_return114_out ),
        .isomorphism_return114_out_13(\SBOX/SBOX[2]/isomorphism_return114_out ),
        .isomorphism_return114_out_15(\SBOX/SBOX[1]/isomorphism_return114_out ),
        .isomorphism_return114_out_17(\SBOX/SBOX[0]/isomorphism_return114_out ),
        .isomorphism_return179_out(\SBOX/SBOX[3]/isomorphism_return179_out ),
        .isomorphism_return179_out_12(\SBOX/SBOX[2]/isomorphism_return179_out ),
        .isomorphism_return179_out_14(\SBOX/SBOX[1]/isomorphism_return179_out ),
        .isomorphism_return179_out_16(\SBOX/SBOX[0]/isomorphism_return179_out ),
        .iv_en(iv_en),
        .iv_mux_out13_out(iv_mux_out13_out),
        .key_derivation_en(key_derivation_en),
        .key_en({key_en[3:2],key_en[0]}),
        .\key_en_pp1_reg[3]_0 (key_en_pp1),
        .\key_en_pp1_reg[3]_1 (key_en_cnt_unit),
        .key_in(key_in),
        .key_out({key_out[31:13],key_out[8:7],key_out[0]}),
        .\key_out_sel_pp1_reg[1]_0 (key_out_sel_pp1),
        .\key_out_sel_pp2_reg[1]_0 (key_out_sel_pp2),
        .key_sel(key_sel),
        .key_sel_mux(key_sel_mux),
        .key_sel_pp1(key_sel_pp1),
        .key_sel_rd(key_sel_rd),
        .last_round(last_round),
        .last_round_pp2_reg_0(last_round_pp2_reg),
        .p_16_in(\SBOX/SBOX[2]/p_16_in ),
        .p_16_in_0(\SBOX/SBOX[1]/p_16_in ),
        .p_16_in_6(\SBOX/SBOX[0]/p_16_in ),
        .p_86_in(\SBOX/SBOX[2]/p_86_in ),
        .p_86_in_11(\SBOX/SBOX[0]/p_86_in ),
        .p_86_in_5(\SBOX/SBOX[1]/p_86_in ),
        .p_93_in(\SBOX/SBOX[2]/p_93_in ),
        .p_93_in_2(\SBOX/SBOX[1]/p_93_in ),
        .p_93_in_8(\SBOX/SBOX[0]/p_93_in ),
        .rk_out_sel(rk_out_sel),
        .rk_out_sel_pp2(rk_out_sel_pp2),
        .\rk_sel_pp1_reg[1]_0 (rk_sel),
        .\round_pp1_reg[0]_0 (AES_CORE_DATAPATH_n_35),
        .\round_pp1_reg[0]_1 (AES_CORE_DATAPATH_n_38),
        .\round_pp1_reg[0]_2 (AES_CORE_DATAPATH_n_62),
        .\round_pp1_reg[3]_0 (AES_CORE_DATAPATH_n_36),
        .\round_pp1_reg[3]_1 (AES_CORE_DATAPATH_n_37),
        .\round_pp1_reg[3]_2 (AES_CORE_DATAPATH_n_39),
        .\round_pp1_reg[3]_3 ({round[3],\rd_count_reg[2] ,round[1:0]}),
        .rst_i(rst_i),
        .sbox_out_enc({sbox_out_enc[19:18],sbox_out_enc[11:10],sbox_out_enc[3:2]}),
        .\sbox_pp2_reg[31]_0 (\sbox_pp2_reg[31] ),
        .\sbox_pp2_reg[5]_0 (AES_CORE_CONTROL_UNIT_n_402));
endmodule

(* ORIG_REF_NAME = "aes_ip" *) 
module switch_elements_aes_ip
   (info_o,
    clk_i,
    rst_i,
    info_o_3_sp_1,
    enable_i,
    \info_o[0]_INST_0_i_4 ,
    info_o_2_sp_1);
  output [30:0]info_o;
  input clk_i;
  input rst_i;
  input info_o_3_sp_1;
  input [31:0]enable_i;
  input \info_o[0]_INST_0_i_4 ;
  input info_o_2_sp_1;

  wire [3:0]\AES_CORE_CONTROL_UNIT/state ;
  wire [31:0]\AES_CORE_DATAPATH/IV_BKP_REGISTERS[0].bkp_1_reg[0]_16 ;
  wire [31:0]\AES_CORE_DATAPATH/IV_BKP_REGISTERS[1].bkp_1_reg[1]_14 ;
  wire [31:0]\AES_CORE_DATAPATH/IV_BKP_REGISTERS[2].bkp_1_reg[2]_12 ;
  wire [31:0]\AES_CORE_DATAPATH/IV_BKP_REGISTERS[3].bkp_1_reg[3]_10 ;
  wire [31:8]\AES_CORE_DATAPATH/add_rk_out ;
  wire [31:0]\AES_CORE_DATAPATH/bus_swap ;
  wire [3:0]\AES_CORE_DATAPATH/col_en_cnt_unit_pp2 ;
  wire [31:8]\AES_CORE_DATAPATH/data_in ;
  wire \AES_CORE_DATAPATH/iv ;
  wire \AES_CORE_DATAPATH/iv_mux_out16_out ;
  wire \AES_CORE_DATAPATH/p_0_in ;
  wire [15:8]\AES_CORE_DATAPATH/p_0_in1_in ;
  wire \AES_CORE_DATAPATH/p_13_out ;
  wire \AES_CORE_DATAPATH/p_17_out ;
  wire \AES_CORE_DATAPATH/p_21_out ;
  wire \AES_CORE_DATAPATH/p_9_out ;
  wire \AES_CORE_DATAPATH/rk_out_sel ;
  wire [95:40]\AES_CORE_DATAPATH/sr_input ;
  wire AES_CORE_n_139;
  wire AES_CORE_n_161;
  wire AES_CORE_n_162;
  wire AES_CORE_n_34;
  wire AES_CORE_n_38;
  wire AES_CORE_n_43;
  wire AES_CORE_n_44;
  wire AES_CORE_n_45;
  wire AES_CORE_n_46;
  wire AES_CORE_n_47;
  wire AES_CORE_n_48;
  wire AES_CORE_n_49;
  wire AES_CORE_n_50;
  wire AES_CORE_n_53;
  wire AES_CORE_n_54;
  wire AES_CORE_n_55;
  wire AES_CORE_n_56;
  wire AES_CORE_n_57;
  wire HOST_INTERFACE_n_100;
  wire HOST_INTERFACE_n_101;
  wire HOST_INTERFACE_n_110;
  wire HOST_INTERFACE_n_111;
  wire HOST_INTERFACE_n_112;
  wire HOST_INTERFACE_n_113;
  wire HOST_INTERFACE_n_114;
  wire HOST_INTERFACE_n_115;
  wire HOST_INTERFACE_n_116;
  wire HOST_INTERFACE_n_117;
  wire HOST_INTERFACE_n_118;
  wire HOST_INTERFACE_n_119;
  wire HOST_INTERFACE_n_120;
  wire HOST_INTERFACE_n_121;
  wire HOST_INTERFACE_n_122;
  wire HOST_INTERFACE_n_123;
  wire HOST_INTERFACE_n_124;
  wire HOST_INTERFACE_n_125;
  wire HOST_INTERFACE_n_126;
  wire HOST_INTERFACE_n_127;
  wire HOST_INTERFACE_n_128;
  wire HOST_INTERFACE_n_129;
  wire HOST_INTERFACE_n_130;
  wire HOST_INTERFACE_n_131;
  wire HOST_INTERFACE_n_132;
  wire HOST_INTERFACE_n_133;
  wire HOST_INTERFACE_n_134;
  wire HOST_INTERFACE_n_135;
  wire HOST_INTERFACE_n_136;
  wire HOST_INTERFACE_n_137;
  wire HOST_INTERFACE_n_138;
  wire HOST_INTERFACE_n_139;
  wire HOST_INTERFACE_n_14;
  wire HOST_INTERFACE_n_140;
  wire HOST_INTERFACE_n_141;
  wire HOST_INTERFACE_n_142;
  wire HOST_INTERFACE_n_143;
  wire HOST_INTERFACE_n_144;
  wire HOST_INTERFACE_n_145;
  wire HOST_INTERFACE_n_146;
  wire HOST_INTERFACE_n_147;
  wire HOST_INTERFACE_n_148;
  wire HOST_INTERFACE_n_149;
  wire HOST_INTERFACE_n_15;
  wire HOST_INTERFACE_n_150;
  wire HOST_INTERFACE_n_151;
  wire HOST_INTERFACE_n_152;
  wire HOST_INTERFACE_n_153;
  wire HOST_INTERFACE_n_154;
  wire HOST_INTERFACE_n_155;
  wire HOST_INTERFACE_n_156;
  wire HOST_INTERFACE_n_157;
  wire HOST_INTERFACE_n_158;
  wire HOST_INTERFACE_n_159;
  wire HOST_INTERFACE_n_16;
  wire HOST_INTERFACE_n_160;
  wire HOST_INTERFACE_n_161;
  wire HOST_INTERFACE_n_162;
  wire HOST_INTERFACE_n_163;
  wire HOST_INTERFACE_n_164;
  wire HOST_INTERFACE_n_165;
  wire HOST_INTERFACE_n_166;
  wire HOST_INTERFACE_n_167;
  wire HOST_INTERFACE_n_168;
  wire HOST_INTERFACE_n_169;
  wire HOST_INTERFACE_n_17;
  wire HOST_INTERFACE_n_170;
  wire HOST_INTERFACE_n_171;
  wire HOST_INTERFACE_n_172;
  wire HOST_INTERFACE_n_173;
  wire HOST_INTERFACE_n_174;
  wire HOST_INTERFACE_n_175;
  wire HOST_INTERFACE_n_176;
  wire HOST_INTERFACE_n_177;
  wire HOST_INTERFACE_n_178;
  wire HOST_INTERFACE_n_179;
  wire HOST_INTERFACE_n_18;
  wire HOST_INTERFACE_n_180;
  wire HOST_INTERFACE_n_181;
  wire HOST_INTERFACE_n_182;
  wire HOST_INTERFACE_n_183;
  wire HOST_INTERFACE_n_184;
  wire HOST_INTERFACE_n_185;
  wire HOST_INTERFACE_n_186;
  wire HOST_INTERFACE_n_187;
  wire HOST_INTERFACE_n_19;
  wire HOST_INTERFACE_n_192;
  wire HOST_INTERFACE_n_193;
  wire HOST_INTERFACE_n_196;
  wire HOST_INTERFACE_n_197;
  wire HOST_INTERFACE_n_198;
  wire HOST_INTERFACE_n_20;
  wire HOST_INTERFACE_n_200;
  wire HOST_INTERFACE_n_201;
  wire HOST_INTERFACE_n_21;
  wire HOST_INTERFACE_n_22;
  wire HOST_INTERFACE_n_23;
  wire HOST_INTERFACE_n_24;
  wire HOST_INTERFACE_n_25;
  wire HOST_INTERFACE_n_26;
  wire HOST_INTERFACE_n_27;
  wire HOST_INTERFACE_n_31;
  wire HOST_INTERFACE_n_36;
  wire HOST_INTERFACE_n_38;
  wire HOST_INTERFACE_n_39;
  wire HOST_INTERFACE_n_40;
  wire HOST_INTERFACE_n_46;
  wire HOST_INTERFACE_n_47;
  wire HOST_INTERFACE_n_48;
  wire HOST_INTERFACE_n_49;
  wire HOST_INTERFACE_n_50;
  wire HOST_INTERFACE_n_51;
  wire HOST_INTERFACE_n_52;
  wire HOST_INTERFACE_n_53;
  wire HOST_INTERFACE_n_55;
  wire HOST_INTERFACE_n_56;
  wire HOST_INTERFACE_n_57;
  wire HOST_INTERFACE_n_58;
  wire HOST_INTERFACE_n_59;
  wire HOST_INTERFACE_n_60;
  wire HOST_INTERFACE_n_61;
  wire HOST_INTERFACE_n_62;
  wire HOST_INTERFACE_n_63;
  wire HOST_INTERFACE_n_64;
  wire HOST_INTERFACE_n_65;
  wire HOST_INTERFACE_n_66;
  wire HOST_INTERFACE_n_67;
  wire HOST_INTERFACE_n_68;
  wire HOST_INTERFACE_n_69;
  wire HOST_INTERFACE_n_70;
  wire HOST_INTERFACE_n_71;
  wire HOST_INTERFACE_n_72;
  wire HOST_INTERFACE_n_73;
  wire HOST_INTERFACE_n_74;
  wire HOST_INTERFACE_n_75;
  wire HOST_INTERFACE_n_76;
  wire HOST_INTERFACE_n_77;
  wire HOST_INTERFACE_n_78;
  wire HOST_INTERFACE_n_79;
  wire HOST_INTERFACE_n_80;
  wire HOST_INTERFACE_n_81;
  wire HOST_INTERFACE_n_82;
  wire HOST_INTERFACE_n_83;
  wire HOST_INTERFACE_n_84;
  wire HOST_INTERFACE_n_85;
  wire HOST_INTERFACE_n_86;
  wire HOST_INTERFACE_n_87;
  wire HOST_INTERFACE_n_88;
  wire HOST_INTERFACE_n_89;
  wire HOST_INTERFACE_n_90;
  wire HOST_INTERFACE_n_91;
  wire HOST_INTERFACE_n_92;
  wire HOST_INTERFACE_n_93;
  wire HOST_INTERFACE_n_94;
  wire HOST_INTERFACE_n_95;
  wire HOST_INTERFACE_n_96;
  wire HOST_INTERFACE_n_97;
  wire HOST_INTERFACE_n_98;
  wire HOST_INTERFACE_n_99;
  wire [1:0]addr;
  wire [1:0]aes_mode;
  wire bypass_rk;
  wire ccf;
  wire ccf_ie;
  wire clk_i;
  wire [3:3]col_en_cnt_unit;
  wire [3:0]col_en_host;
  wire [3:1]col_out;
  wire [1:0]data_type;
  wire [31:0]enable_i;
  wire enc_dec;
  wire first_block;
  wire [30:0]info_o;
  wire \info_o[0]_INST_0_i_4 ;
  wire info_o_2_sn_1;
  wire info_o_3_sn_1;
  wire [2:0]iv_en;
  wire key_derivation_en;
  wire [3:0]key_en;
  wire [12:4]key_out;
  wire [0:0]key_sel_rd;
  wire [1:0]op_mode;
  wire [2:2]round;
  wire rst_i;

  assign info_o_2_sn_1 = info_o_2_sp_1;
  assign info_o_3_sn_1 = info_o_3_sp_1;
  switch_elements_aes_core AES_CORE
       (.\CD[0].col[3][0]_i_2 (HOST_INTERFACE_n_57),
        .\CD[0].col[3][0]_i_2_0 (HOST_INTERFACE_n_192),
        .\CD[0].col[3][0]_i_4 (HOST_INTERFACE_n_58),
        .\CD[0].col[3][10]_i_12 (HOST_INTERFACE_n_38),
        .\CD[0].col[3][10]_i_6 (HOST_INTERFACE_n_193),
        .\CD[0].col[3][31]_i_22 (HOST_INTERFACE_n_31),
        .\CD[0].col[3][5]_i_2 (HOST_INTERFACE_n_201),
        .\CD[2].col_reg[1][31] ({\AES_CORE_DATAPATH/sr_input [95:88],\AES_CORE_DATAPATH/sr_input [79:72],\AES_CORE_DATAPATH/sr_input [63:56],\AES_CORE_DATAPATH/sr_input [47:40]}),
        .\CD[3].col_reg[0][31] (addr),
        .\CD[3].col_reg[0][31]_0 (HOST_INTERFACE_n_23),
        .D(\AES_CORE_DATAPATH/p_0_in1_in ),
        .E(\AES_CORE_DATAPATH/p_21_out ),
        .\FSM_sequential_state_reg[0] (AES_CORE_n_46),
        .\FSM_sequential_state_reg[0]_0 (AES_CORE_n_139),
        .\FSM_sequential_state_reg[0]_1 (HOST_INTERFACE_n_27),
        .\FSM_sequential_state_reg[0]_2 (HOST_INTERFACE_n_46),
        .\FSM_sequential_state_reg[0]_3 (HOST_INTERFACE_n_21),
        .\FSM_sequential_state_reg[1] (HOST_INTERFACE_n_24),
        .\FSM_sequential_state_reg[2] (AES_CORE_n_43),
        .\FSM_sequential_state_reg[2]_0 (AES_CORE_n_45),
        .\FSM_sequential_state_reg[2]_1 (col_en_cnt_unit),
        .\FSM_sequential_state_reg[2]_2 (AES_CORE_n_57),
        .\FSM_sequential_state_reg[2]_3 (HOST_INTERFACE_n_51),
        .\FSM_sequential_state_reg[3] (AES_CORE_n_44),
        .\FSM_sequential_state_reg[3]_0 (AES_CORE_n_54),
        .\FSM_sequential_state_reg[3]_1 (AES_CORE_n_55),
        .\FSM_sequential_state_reg[3]_2 (HOST_INTERFACE_n_22),
        .\FSM_sequential_state_reg[3]_3 (HOST_INTERFACE_n_47),
        .\FSM_sequential_state_reg[3]_4 (HOST_INTERFACE_n_52),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][31] (\AES_CORE_DATAPATH/IV_BKP_REGISTERS[0].bkp_1_reg[0]_16 ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][0] (HOST_INTERFACE_n_63),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 (\AES_CORE_DATAPATH/p_0_in ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][15] ({HOST_INTERFACE_n_94,HOST_INTERFACE_n_95,HOST_INTERFACE_n_96,HOST_INTERFACE_n_97,HOST_INTERFACE_n_98,HOST_INTERFACE_n_99,HOST_INTERFACE_n_100,HOST_INTERFACE_n_101}),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][16] (HOST_INTERFACE_n_127),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][17] (HOST_INTERFACE_n_131),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][18] (HOST_INTERFACE_n_135),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][19] (HOST_INTERFACE_n_139),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][1] (HOST_INTERFACE_n_67),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][20] (HOST_INTERFACE_n_143),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][21] (HOST_INTERFACE_n_147),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][22] (HOST_INTERFACE_n_151),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][23] (HOST_INTERFACE_n_155),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][24] (HOST_INTERFACE_n_172),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][25] (HOST_INTERFACE_n_174),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][26] (HOST_INTERFACE_n_176),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][27] (HOST_INTERFACE_n_178),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][28] (HOST_INTERFACE_n_180),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][29] (HOST_INTERFACE_n_182),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][2] (HOST_INTERFACE_n_71),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][30] (HOST_INTERFACE_n_184),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][31] (HOST_INTERFACE_n_186),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][3] (HOST_INTERFACE_n_75),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][4] (HOST_INTERFACE_n_79),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][5] (HOST_INTERFACE_n_83),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][6] (HOST_INTERFACE_n_87),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][7] (HOST_INTERFACE_n_91),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][31] (\AES_CORE_DATAPATH/IV_BKP_REGISTERS[1].bkp_1_reg[1]_14 ),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][0] (HOST_INTERFACE_n_62),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 (HOST_INTERFACE_n_198),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][10] (HOST_INTERFACE_n_113),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][11] (HOST_INTERFACE_n_115),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][12] (HOST_INTERFACE_n_117),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][13] (HOST_INTERFACE_n_119),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][14] (HOST_INTERFACE_n_121),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][15] (HOST_INTERFACE_n_123),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][16] (HOST_INTERFACE_n_126),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][17] (HOST_INTERFACE_n_130),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][18] (HOST_INTERFACE_n_134),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][19] (HOST_INTERFACE_n_138),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][1] (HOST_INTERFACE_n_66),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][20] (HOST_INTERFACE_n_142),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][21] (HOST_INTERFACE_n_146),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][22] (HOST_INTERFACE_n_150),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][23] (HOST_INTERFACE_n_154),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][2] (HOST_INTERFACE_n_70),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][31] (HOST_INTERFACE_n_200),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 ({HOST_INTERFACE_n_156,HOST_INTERFACE_n_157,HOST_INTERFACE_n_158,HOST_INTERFACE_n_159,HOST_INTERFACE_n_160,HOST_INTERFACE_n_161,HOST_INTERFACE_n_162,HOST_INTERFACE_n_163}),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][3] (HOST_INTERFACE_n_74),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][4] (HOST_INTERFACE_n_78),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][5] (HOST_INTERFACE_n_82),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][6] (HOST_INTERFACE_n_86),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][7] (HOST_INTERFACE_n_90),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][8] (HOST_INTERFACE_n_93),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][9] (HOST_INTERFACE_n_111),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][31] (\AES_CORE_DATAPATH/IV_BKP_REGISTERS[2].bkp_1_reg[2]_12 ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][0] (HOST_INTERFACE_n_61),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 (HOST_INTERFACE_n_197),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][10] (HOST_INTERFACE_n_112),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][11] (HOST_INTERFACE_n_114),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][12] (HOST_INTERFACE_n_116),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][13] (HOST_INTERFACE_n_118),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][14] (HOST_INTERFACE_n_120),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][15] (HOST_INTERFACE_n_122),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][16] (HOST_INTERFACE_n_125),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][17] (HOST_INTERFACE_n_129),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][18] (HOST_INTERFACE_n_133),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][19] (HOST_INTERFACE_n_137),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][1] (HOST_INTERFACE_n_65),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][20] (HOST_INTERFACE_n_141),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][21] (HOST_INTERFACE_n_145),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][22] (HOST_INTERFACE_n_149),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][23] (HOST_INTERFACE_n_153),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][2] (HOST_INTERFACE_n_69),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][31] ({HOST_INTERFACE_n_164,HOST_INTERFACE_n_165,HOST_INTERFACE_n_166,HOST_INTERFACE_n_167,HOST_INTERFACE_n_168,HOST_INTERFACE_n_169,HOST_INTERFACE_n_170,HOST_INTERFACE_n_171}),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][3] (HOST_INTERFACE_n_73),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][4] (HOST_INTERFACE_n_77),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][5] (HOST_INTERFACE_n_81),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][6] (HOST_INTERFACE_n_85),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][7] (HOST_INTERFACE_n_89),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][8] (HOST_INTERFACE_n_92),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][9] (HOST_INTERFACE_n_110),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][31] (\AES_CORE_DATAPATH/IV_BKP_REGISTERS[3].bkp_1_reg[3]_10 ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][0] (HOST_INTERFACE_n_60),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][0]_0 (HOST_INTERFACE_n_196),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][16] (HOST_INTERFACE_n_124),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][17] (HOST_INTERFACE_n_128),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][18] (HOST_INTERFACE_n_132),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][19] (HOST_INTERFACE_n_136),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][1] (HOST_INTERFACE_n_64),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][20] (HOST_INTERFACE_n_140),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][21] (HOST_INTERFACE_n_144),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][22] (HOST_INTERFACE_n_148),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][23] (HOST_INTERFACE_n_152),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][24] (HOST_INTERFACE_n_173),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][25] (HOST_INTERFACE_n_175),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][26] (HOST_INTERFACE_n_177),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][27] (HOST_INTERFACE_n_179),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][28] (HOST_INTERFACE_n_181),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][29] (HOST_INTERFACE_n_183),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][2] (HOST_INTERFACE_n_68),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][30] (HOST_INTERFACE_n_185),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][31] (HOST_INTERFACE_n_56),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 (HOST_INTERFACE_n_187),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][3] (HOST_INTERFACE_n_72),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][4] (HOST_INTERFACE_n_76),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][5] (HOST_INTERFACE_n_80),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][6] (HOST_INTERFACE_n_84),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][7] (HOST_INTERFACE_n_88),
        .\IV_BKP_REGISTERS[3].iv_reg[3][0] (\AES_CORE_DATAPATH/iv ),
        .\KR[1].key_host_reg[2][0] (\AES_CORE_DATAPATH/p_17_out ),
        .\KR[1].key_reg[2][12] ({key_out[12:9],key_out[6],key_out[4]}),
        .\KR[2].key_host_reg[1][0] (\AES_CORE_DATAPATH/p_13_out ),
        .\KR[3].key_host_reg[0][0] (\AES_CORE_DATAPATH/p_9_out ),
        .\KR[3].key_reg[0][31] (HOST_INTERFACE_n_26),
        .Q(\AES_CORE_CONTROL_UNIT/state ),
        .\aes_cr_reg[2] (col_out),
        .\aes_cr_reg[4] (AES_CORE_n_53),
        .\aes_cr_reg[5] (AES_CORE_n_161),
        .\aes_cr_reg[5]_0 (AES_CORE_n_162),
        .bus_swap(\AES_CORE_DATAPATH/bus_swap ),
        .bypass_rk(bypass_rk),
        .ccf(ccf),
        .ccf_reg(AES_CORE_n_38),
        .ccf_reg_0(HOST_INTERFACE_n_40),
        .clk_i(clk_i),
        .\col_en_cnt_unit_pp1_reg[3] (HOST_INTERFACE_n_55),
        .\col_en_cnt_unit_pp2_reg[3] (\AES_CORE_DATAPATH/col_en_cnt_unit_pp2 ),
        .col_en_host(col_en_host),
        .\col_sel_pp1_reg[1] (HOST_INTERFACE_n_53),
        .data_in({\AES_CORE_DATAPATH/data_in [31:24],\AES_CORE_DATAPATH/data_in [15:8]}),
        .enable_i(enable_i),
        .\enable_i[6]_0 (AES_CORE_n_49),
        .enable_i_0_sp_1(AES_CORE_n_34),
        .enable_i_2_sp_1(AES_CORE_n_56),
        .enable_i_3_sp_1(AES_CORE_n_48),
        .enable_i_6_sp_1(AES_CORE_n_47),
        .enc_dec(enc_dec),
        .first_block(first_block),
        .info_o({info_o[30:4],info_o[0]}),
        .\info_o[0]_0 (info_o_3_sn_1),
        .\info_o[0]_1 ({ccf_ie,aes_mode,op_mode,data_type}),
        .\info_o[28]_INST_0_i_15 (HOST_INTERFACE_n_49),
        .\info_o[28]_INST_0_i_15_0 (HOST_INTERFACE_n_50),
        .\info_o[31] (HOST_INTERFACE_n_48),
        .\info_o[31]_0 (HOST_INTERFACE_n_15),
        .\info_o[31]_INST_0_i_12 (HOST_INTERFACE_n_36),
        .info_o_0_sp_1(HOST_INTERFACE_n_39),
        .info_o_10_sp_1(HOST_INTERFACE_n_18),
        .info_o_11_sp_1(HOST_INTERFACE_n_19),
        .info_o_12_sp_1(HOST_INTERFACE_n_20),
        .info_o_4_sp_1(HOST_INTERFACE_n_14),
        .info_o_6_sp_1(HOST_INTERFACE_n_16),
        .info_o_9_sp_1(HOST_INTERFACE_n_17),
        .iv_en(iv_en),
        .iv_mux_out16_out(\AES_CORE_DATAPATH/iv_mux_out16_out ),
        .key_derivation_en(key_derivation_en),
        .key_en(key_en),
        .\key_en_pp1_reg[3] (HOST_INTERFACE_n_25),
        .key_sel_rd(key_sel_rd),
        .last_round_pp2_reg({\AES_CORE_DATAPATH/add_rk_out [31:24],\AES_CORE_DATAPATH/add_rk_out [15:8]}),
        .\rd_count_reg[2] (round),
        .\rd_count_reg[3] (AES_CORE_n_50),
        .rk_out_sel(\AES_CORE_DATAPATH/rk_out_sel ),
        .rst_i(rst_i),
        .\sbox_pp2_reg[31] (HOST_INTERFACE_n_59));
  switch_elements_host_interface HOST_INTERFACE
       (.\CD[0].col[3][10]_i_12 (col_en_cnt_unit),
        .\CD[1].col_reg[2][31] ({HOST_INTERFACE_n_156,HOST_INTERFACE_n_157,HOST_INTERFACE_n_158,HOST_INTERFACE_n_159,HOST_INTERFACE_n_160,HOST_INTERFACE_n_161,HOST_INTERFACE_n_162,HOST_INTERFACE_n_163}),
        .\CD[2].col_reg[1][15] ({HOST_INTERFACE_n_94,HOST_INTERFACE_n_95,HOST_INTERFACE_n_96,HOST_INTERFACE_n_97,HOST_INTERFACE_n_98,HOST_INTERFACE_n_99,HOST_INTERFACE_n_100,HOST_INTERFACE_n_101}),
        .\CD[2].col_reg[1][31] ({HOST_INTERFACE_n_164,HOST_INTERFACE_n_165,HOST_INTERFACE_n_166,HOST_INTERFACE_n_167,HOST_INTERFACE_n_168,HOST_INTERFACE_n_169,HOST_INTERFACE_n_170,HOST_INTERFACE_n_171}),
        .D(\AES_CORE_DATAPATH/p_0_in1_in ),
        .E(\AES_CORE_DATAPATH/p_21_out ),
        .\FSM_sequential_state_reg[0]_0 (HOST_INTERFACE_n_23),
        .\FSM_sequential_state_reg[0]_1 (HOST_INTERFACE_n_36),
        .\FSM_sequential_state_reg[0]_2 (AES_CORE_n_43),
        .\FSM_sequential_state_reg[0]_3 (round),
        .\FSM_sequential_state_reg[0]_4 (AES_CORE_n_55),
        .\FSM_sequential_state_reg[1]_0 (AES_CORE_n_57),
        .\FSM_sequential_state_reg[1]_1 (AES_CORE_n_44),
        .\FSM_sequential_state_reg[1]_2 (AES_CORE_n_53),
        .\FSM_sequential_state_reg[2]_0 (HOST_INTERFACE_n_26),
        .\FSM_sequential_state_reg[2]_1 (HOST_INTERFACE_n_27),
        .\FSM_sequential_state_reg[2]_2 (HOST_INTERFACE_n_49),
        .\FSM_sequential_state_reg[2]_3 (HOST_INTERFACE_n_50),
        .\FSM_sequential_state_reg[2]_4 (HOST_INTERFACE_n_56),
        .\FSM_sequential_state_reg[2]_5 (\AES_CORE_DATAPATH/p_13_out ),
        .\FSM_sequential_state_reg[3] (HOST_INTERFACE_n_46),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][0] (HOST_INTERFACE_n_63),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][16] (HOST_INTERFACE_n_127),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][17] (HOST_INTERFACE_n_131),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][18] (HOST_INTERFACE_n_135),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][19] (HOST_INTERFACE_n_139),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][1] (HOST_INTERFACE_n_67),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][20] (HOST_INTERFACE_n_143),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][21] (HOST_INTERFACE_n_147),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][22] (HOST_INTERFACE_n_151),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][23] (HOST_INTERFACE_n_155),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][2] (HOST_INTERFACE_n_71),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][3] (HOST_INTERFACE_n_75),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][4] (HOST_INTERFACE_n_79),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][5] (HOST_INTERFACE_n_83),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][6] (HOST_INTERFACE_n_87),
        .\IV_BKP_REGISTERS[0].bkp_1_reg[0][7] (HOST_INTERFACE_n_91),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][31] (\AES_CORE_DATAPATH/IV_BKP_REGISTERS[0].bkp_1_reg[0]_16 ),
        .\IV_BKP_REGISTERS[0].bkp_reg[0][8] (AES_CORE_n_162),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][0] (HOST_INTERFACE_n_62),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][16] (HOST_INTERFACE_n_126),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][17] (HOST_INTERFACE_n_130),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][18] (HOST_INTERFACE_n_134),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][19] (HOST_INTERFACE_n_138),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][1] (HOST_INTERFACE_n_66),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][20] (HOST_INTERFACE_n_142),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][21] (HOST_INTERFACE_n_146),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][22] (HOST_INTERFACE_n_150),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][23] (HOST_INTERFACE_n_154),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][2] (HOST_INTERFACE_n_70),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][3] (HOST_INTERFACE_n_74),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][4] (HOST_INTERFACE_n_78),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][5] (HOST_INTERFACE_n_82),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][6] (HOST_INTERFACE_n_86),
        .\IV_BKP_REGISTERS[1].bkp_1_reg[1][7] (HOST_INTERFACE_n_90),
        .\IV_BKP_REGISTERS[1].bkp_reg[1][31] (\AES_CORE_DATAPATH/IV_BKP_REGISTERS[1].bkp_1_reg[1]_14 ),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][0] (HOST_INTERFACE_n_61),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][16] (HOST_INTERFACE_n_125),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][17] (HOST_INTERFACE_n_129),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][18] (HOST_INTERFACE_n_133),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][19] (HOST_INTERFACE_n_137),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][1] (HOST_INTERFACE_n_65),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][20] (HOST_INTERFACE_n_141),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][21] (HOST_INTERFACE_n_145),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][22] (HOST_INTERFACE_n_149),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][23] (HOST_INTERFACE_n_153),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][2] (HOST_INTERFACE_n_69),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][3] (HOST_INTERFACE_n_73),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][4] (HOST_INTERFACE_n_77),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][5] (HOST_INTERFACE_n_81),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][6] (HOST_INTERFACE_n_85),
        .\IV_BKP_REGISTERS[2].bkp_1_reg[2][7] (HOST_INTERFACE_n_89),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][31] (\AES_CORE_DATAPATH/IV_BKP_REGISTERS[2].bkp_1_reg[2]_12 ),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 ({\AES_CORE_DATAPATH/sr_input [95:88],\AES_CORE_DATAPATH/sr_input [79:72],\AES_CORE_DATAPATH/sr_input [63:56],\AES_CORE_DATAPATH/sr_input [47:40]}),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 ({\AES_CORE_DATAPATH/add_rk_out [31:24],\AES_CORE_DATAPATH/add_rk_out [15:8]}),
        .\IV_BKP_REGISTERS[2].bkp_reg[2][31]_2 (AES_CORE_n_139),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][0] (HOST_INTERFACE_n_60),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][16] (HOST_INTERFACE_n_124),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][17] (HOST_INTERFACE_n_128),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][18] (HOST_INTERFACE_n_132),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][19] (HOST_INTERFACE_n_136),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][1] (HOST_INTERFACE_n_64),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][20] (HOST_INTERFACE_n_140),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][21] (HOST_INTERFACE_n_144),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][22] (HOST_INTERFACE_n_148),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][23] (HOST_INTERFACE_n_152),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][2] (HOST_INTERFACE_n_68),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][3] (HOST_INTERFACE_n_72),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][4] (HOST_INTERFACE_n_76),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][5] (HOST_INTERFACE_n_80),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][6] (HOST_INTERFACE_n_84),
        .\IV_BKP_REGISTERS[3].bkp_1_reg[3][7] (HOST_INTERFACE_n_88),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][0] (\AES_CORE_DATAPATH/col_en_cnt_unit_pp2 ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][31] (\AES_CORE_DATAPATH/IV_BKP_REGISTERS[3].bkp_1_reg[3]_10 ),
        .\IV_BKP_REGISTERS[3].bkp_reg[3][8] (AES_CORE_n_161),
        .\IV_BKP_REGISTERS[3].iv_reg[3][0] (AES_CORE_n_50),
        .\IV_BKP_REGISTERS[3].iv_reg[3][0]_0 (AES_CORE_n_47),
        .\IV_BKP_REGISTERS[3].iv_reg[3][0]_1 (AES_CORE_n_54),
        .\KR[0].key_host_reg[3][0] (AES_CORE_n_46),
        .\KR[1].key_host_reg[2][0] (AES_CORE_n_49),
        .Q(addr),
        .\aes_cr_reg[0]_0 (HOST_INTERFACE_n_15),
        .\aes_cr_reg[0]_1 (HOST_INTERFACE_n_22),
        .\aes_cr_reg[0]_2 (HOST_INTERFACE_n_48),
        .\aes_cr_reg[0]_3 (AES_CORE_n_48),
        .\aes_cr_reg[10]_0 (HOST_INTERFACE_n_20),
        .\aes_cr_reg[3]_0 (HOST_INTERFACE_n_47),
        .\aes_cr_reg[4]_0 (HOST_INTERFACE_n_14),
        .\aes_cr_reg[4]_1 (HOST_INTERFACE_n_21),
        .\aes_cr_reg[4]_2 (HOST_INTERFACE_n_24),
        .\aes_cr_reg[4]_3 (HOST_INTERFACE_n_51),
        .\aes_cr_reg[4]_4 (HOST_INTERFACE_n_53),
        .\aes_cr_reg[4]_5 (HOST_INTERFACE_n_57),
        .\aes_cr_reg[4]_6 (HOST_INTERFACE_n_59),
        .\aes_cr_reg[5]_0 (HOST_INTERFACE_n_25),
        .\aes_cr_reg[5]_1 (HOST_INTERFACE_n_92),
        .\aes_cr_reg[5]_10 (HOST_INTERFACE_n_117),
        .\aes_cr_reg[5]_11 (HOST_INTERFACE_n_118),
        .\aes_cr_reg[5]_12 (HOST_INTERFACE_n_119),
        .\aes_cr_reg[5]_13 (HOST_INTERFACE_n_120),
        .\aes_cr_reg[5]_14 (HOST_INTERFACE_n_121),
        .\aes_cr_reg[5]_15 (HOST_INTERFACE_n_122),
        .\aes_cr_reg[5]_16 (HOST_INTERFACE_n_123),
        .\aes_cr_reg[5]_17 (HOST_INTERFACE_n_172),
        .\aes_cr_reg[5]_18 (HOST_INTERFACE_n_173),
        .\aes_cr_reg[5]_19 (HOST_INTERFACE_n_174),
        .\aes_cr_reg[5]_2 (HOST_INTERFACE_n_93),
        .\aes_cr_reg[5]_20 (HOST_INTERFACE_n_175),
        .\aes_cr_reg[5]_21 (HOST_INTERFACE_n_176),
        .\aes_cr_reg[5]_22 (HOST_INTERFACE_n_177),
        .\aes_cr_reg[5]_23 (HOST_INTERFACE_n_178),
        .\aes_cr_reg[5]_24 (HOST_INTERFACE_n_179),
        .\aes_cr_reg[5]_25 (HOST_INTERFACE_n_180),
        .\aes_cr_reg[5]_26 (HOST_INTERFACE_n_181),
        .\aes_cr_reg[5]_27 (HOST_INTERFACE_n_182),
        .\aes_cr_reg[5]_28 (HOST_INTERFACE_n_183),
        .\aes_cr_reg[5]_29 (HOST_INTERFACE_n_184),
        .\aes_cr_reg[5]_3 (HOST_INTERFACE_n_110),
        .\aes_cr_reg[5]_30 (HOST_INTERFACE_n_185),
        .\aes_cr_reg[5]_31 (HOST_INTERFACE_n_186),
        .\aes_cr_reg[5]_32 (HOST_INTERFACE_n_187),
        .\aes_cr_reg[5]_33 (\AES_CORE_DATAPATH/iv ),
        .\aes_cr_reg[5]_34 (HOST_INTERFACE_n_200),
        .\aes_cr_reg[5]_35 (HOST_INTERFACE_n_201),
        .\aes_cr_reg[5]_4 (HOST_INTERFACE_n_111),
        .\aes_cr_reg[5]_5 (HOST_INTERFACE_n_112),
        .\aes_cr_reg[5]_6 (HOST_INTERFACE_n_113),
        .\aes_cr_reg[5]_7 (HOST_INTERFACE_n_114),
        .\aes_cr_reg[5]_8 (HOST_INTERFACE_n_115),
        .\aes_cr_reg[5]_9 (HOST_INTERFACE_n_116),
        .\aes_cr_reg[6]_0 (HOST_INTERFACE_n_16),
        .\aes_cr_reg[6]_1 (HOST_INTERFACE_n_52),
        .\aes_cr_reg[6]_2 (HOST_INTERFACE_n_55),
        .\aes_cr_reg[7]_0 ({ccf_ie,aes_mode,op_mode,data_type}),
        .\aes_cr_reg[7]_1 (HOST_INTERFACE_n_17),
        .\aes_cr_reg[8]_0 (HOST_INTERFACE_n_18),
        .\aes_cr_reg[9]_0 (HOST_INTERFACE_n_19),
        .bus_swap(\AES_CORE_DATAPATH/bus_swap ),
        .bypass_rk(bypass_rk),
        .ccf(ccf),
        .ccf_reg_0(AES_CORE_n_45),
        .clk_i(clk_i),
        .\cnt_reg[0]_0 (AES_CORE_n_34),
        .\col_en_cnt_unit_pp2_reg[0] (\AES_CORE_DATAPATH/p_0_in ),
        .\col_en_cnt_unit_pp2_reg[1] (HOST_INTERFACE_n_198),
        .\col_en_cnt_unit_pp2_reg[2] (HOST_INTERFACE_n_197),
        .\col_en_cnt_unit_pp2_reg[3] (HOST_INTERFACE_n_193),
        .\col_en_cnt_unit_pp2_reg[3]_0 (HOST_INTERFACE_n_196),
        .col_en_host(col_en_host),
        .data_in({\AES_CORE_DATAPATH/data_in [31:24],\AES_CORE_DATAPATH/data_in [15:8]}),
        .enable_i({enable_i[12:8],enable_i[6:0]}),
        .\enable_i[1]_0 (HOST_INTERFACE_n_39),
        .\enable_i[2]_0 (HOST_INTERFACE_n_40),
        .\enable_i[2]_1 (\AES_CORE_DATAPATH/p_9_out ),
        .\enable_i[4] (\AES_CORE_DATAPATH/p_17_out ),
        .enable_i_1_sp_1(HOST_INTERFACE_n_31),
        .enable_i_2_sp_1(HOST_INTERFACE_n_38),
        .enc_dec(enc_dec),
        .first_block(first_block),
        .first_block_reg_0(HOST_INTERFACE_n_58),
        .first_block_reg_1(HOST_INTERFACE_n_192),
        .info_o(info_o[3:1]),
        .\info_o[0]_INST_0_i_4 (\info_o[0]_INST_0_i_4 ),
        .\info_o[12] ({key_out[12:9],key_out[6],key_out[4]}),
        .\info_o[31]_INST_0_i_15 (AES_CORE_n_56),
        .\info_o[3] (col_out),
        .\info_o[3]_0 (info_o_3_sn_1),
        .info_o_1_sp_1(AES_CORE_n_38),
        .info_o_2_sp_1(info_o_2_sn_1),
        .iv_en(iv_en),
        .iv_mux_out16_out(\AES_CORE_DATAPATH/iv_mux_out16_out ),
        .key_derivation_en(key_derivation_en),
        .key_en(key_en),
        .key_sel_rd(key_sel_rd),
        .rk_out_sel(\AES_CORE_DATAPATH/rk_out_sel ),
        .rk_out_sel_pp1_reg(\AES_CORE_CONTROL_UNIT/state ),
        .rst_i(rst_i));
endmodule

(* ORIG_REF_NAME = "control_unit" *) 
module switch_elements_control_unit
   (info_o,
    \aes_cr_reg[7] ,
    ccf_reg,
    Q,
    \FSM_sequential_state_reg[2]_0 ,
    \FSM_sequential_state_reg[3]_0 ,
    \FSM_sequential_state_reg[2]_1 ,
    \FSM_sequential_state_reg[0]_0 ,
    D,
    \rd_count_reg[3]_0 ,
    \rd_count_reg[3]_1 ,
    \FSM_sequential_state_reg[1]_0 ,
    \FSM_sequential_state_reg[0]_1 ,
    \FSM_sequential_state_reg[2]_2 ,
    key_sel,
    \aes_cr_reg[4] ,
    \FSM_sequential_state_reg[2]_3 ,
    \FSM_sequential_state_reg[3]_1 ,
    \FSM_sequential_state_reg[3]_2 ,
    \FSM_sequential_state_reg[2]_4 ,
    bypass_key_en,
    last_round,
    \FSM_sequential_state_reg[2]_5 ,
    key_sel_mux,
    \CD[3].col_reg[0][31] ,
    \CD[1].col_reg[2][23] ,
    \CD[2].col_reg[1][23] ,
    \CD[0].col_reg[3][31] ,
    \CD[3].col_reg[0][31]_0 ,
    \CD[0].col_reg[3][31]_0 ,
    \CD[1].col_reg[2][31] ,
    \CD[2].col_reg[1][31] ,
    \FSM_sequential_state_reg[0]_2 ,
    \IV_BKP_REGISTERS[2].iv_reg[2][8] ,
    \IV_BKP_REGISTERS[2].iv_reg[2][9] ,
    data_in,
    \IV_BKP_REGISTERS[2].iv_reg[2][14] ,
    \IV_BKP_REGISTERS[2].iv_reg[2][15] ,
    \IV_BKP_REGISTERS[2].iv_reg[2][24] ,
    \IV_BKP_REGISTERS[2].iv_reg[2][25] ,
    \IV_BKP_REGISTERS[2].iv_reg[2][26] ,
    \IV_BKP_REGISTERS[2].iv_reg[2][27] ,
    \IV_BKP_REGISTERS[2].iv_reg[2][29] ,
    \IV_BKP_REGISTERS[2].iv_reg[2][30] ,
    \IV_BKP_REGISTERS[2].iv_reg[2][31] ,
    \KR[3].key_reg[0][31] ,
    \CD[3].col_reg[0][0] ,
    \FSM_sequential_state_reg[2]_6 ,
    \FSM_sequential_state_reg[3]_3 ,
    \FSM_sequential_state_reg[3]_4 ,
    \CD[3].col_reg[0][7] ,
    \CD[3].col_reg[0][15] ,
    \CD[3].col_reg[0][31]_1 ,
    \CD[3].col_reg[0][1] ,
    \CD[3].col_reg[0][6] ,
    \CD[3].col_reg[0][14] ,
    \CD[3].col_reg[0][30] ,
    \CD[3].col_reg[0][2] ,
    \CD[3].col_reg[0][5] ,
    \CD[3].col_reg[0][13] ,
    \CD[3].col_reg[0][29] ,
    \CD[3].col_reg[0][3] ,
    \CD[3].col_reg[0][4] ,
    \CD[3].col_reg[0][12] ,
    \CD[3].col_reg[0][28] ,
    \CD[3].col_reg[0][11] ,
    \CD[3].col_reg[0][27] ,
    \CD[3].col_reg[0][10] ,
    \CD[3].col_reg[0][26] ,
    \CD[3].col_reg[0][9] ,
    \CD[3].col_reg[0][25] ,
    \CD[3].col_reg[0][8] ,
    \CD[3].col_reg[0][24] ,
    \CD[3].col_reg[0][23] ,
    \CD[3].col_reg[0][22] ,
    \CD[3].col_reg[0][21] ,
    \CD[3].col_reg[0][20] ,
    \CD[3].col_reg[0][19] ,
    \CD[3].col_reg[0][18] ,
    \CD[3].col_reg[0][17] ,
    \CD[3].col_reg[0][16] ,
    first_block_reg,
    iv_mux_out13_out,
    \col_en_cnt_unit_pp2_reg[3] ,
    first_block_reg_0,
    \IV_BKP_REGISTERS[3].iv_reg[3][8] ,
    \IV_BKP_REGISTERS[3].iv_reg[3][9] ,
    \IV_BKP_REGISTERS[3].iv_reg[3][14] ,
    \IV_BKP_REGISTERS[3].iv_reg[3][15] ,
    \IV_BKP_REGISTERS[3].iv_reg[3][24] ,
    \IV_BKP_REGISTERS[3].iv_reg[3][25] ,
    \IV_BKP_REGISTERS[3].iv_reg[3][26] ,
    \IV_BKP_REGISTERS[3].iv_reg[3][27] ,
    \IV_BKP_REGISTERS[3].iv_reg[3][29] ,
    \IV_BKP_REGISTERS[3].iv_reg[3][30] ,
    \IV_BKP_REGISTERS[3].iv_reg[3][31] ,
    E,
    \col_en_cnt_unit_pp2_reg[2] ,
    \col_en_cnt_unit_pp2_reg[1] ,
    \col_en_cnt_unit_pp2_reg[0] ,
    enc_dec_sbox,
    \FSM_sequential_state_reg[3]_5 ,
    \FSM_sequential_state_reg[3]_6 ,
    \key_en_pp1_reg[3] ,
    \key_en_pp1_reg[2] ,
    \key_en_pp1_reg[1] ,
    \key_en_pp1_reg[0] ,
    \aes_cr_reg[5] ,
    \aes_cr_reg[5]_0 ,
    \key_out_sel_pp1_reg[1] ,
    \enable_i[31] ,
    add_rk_sel,
    \FSM_sequential_state_reg[3]_7 ,
    \FSM_sequential_state_reg[3]_8 ,
    first_block_reg_1,
    isomorphism_return179_out,
    isomorphism_return114_out,
    isomorphism_return179_out_0,
    isomorphism_return114_out_1,
    isomorphism_return179_out_2,
    isomorphism_return114_out_3,
    isomorphism_return179_out_4,
    isomorphism_return114_out_5,
    \info_o[31] ,
    key_out,
    \info_o[31]_0 ,
    info_o_0_sp_1,
    col_out,
    info_o_4_sp_1,
    info_o_6_sp_1,
    info_o_9_sp_1,
    info_o_10_sp_1,
    info_o_11_sp_1,
    info_o_12_sp_1,
    \FSM_sequential_state_reg[0]_3 ,
    \col_en_cnt_unit_pp1_reg[3] ,
    \FSM_sequential_state_reg[2]_7 ,
    enable_i,
    ccf,
    ccf_reg_0,
    \col_sel_pp1_reg[1] ,
    \info_o[0]_0 ,
    \info_o[31]_1 ,
    \key_en_pp1_reg[3]_0 ,
    \FSM_sequential_state_reg[3]_9 ,
    \FSM_sequential_state_reg[3]_10 ,
    \FSM_sequential_state_reg[3]_11 ,
    \FSM_sequential_state_reg[0]_4 ,
    \FSM_sequential_state_reg[0]_5 ,
    key_en,
    \KR[2].key_reg[1][31] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][0] ,
    \CD[2].col_reg[1][31]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][31] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][0] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][0] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][0] ,
    \CD[1].col_reg[2][31]_0 ,
    add_rk_out,
    \IV_BKP_REGISTERS[0].bkp_reg[0][31] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 ,
    \CD[2].col_reg[1][31]_1 ,
    \CD[2].col_reg[1][0] ,
    \CD[2].col_reg[1][0]_0 ,
    \info_o[31]_2 ,
    bus_swap,
    \IV_BKP_REGISTERS[3].bkp_reg[3][1] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][1] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][1] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][1] ,
    \CD[2].col_reg[1][1] ,
    \CD[2].col_reg[1][1]_0 ,
    \CD[0].col[3][1]_i_2_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][2] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][2] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][2] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][2] ,
    \CD[2].col_reg[1][2] ,
    \CD[2].col_reg[1][2]_0 ,
    \CD[0].col[3][2]_i_2_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][3] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][3] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][3] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][3] ,
    \CD[2].col_reg[1][3] ,
    \CD[2].col_reg[1][3]_0 ,
    \CD[0].col[3][3]_i_2_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][4] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][4] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][4] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][4] ,
    \CD[2].col_reg[1][4] ,
    \CD[2].col_reg[1][4]_0 ,
    \CD[0].col[3][4]_i_2_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][5] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][5] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][5] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][5] ,
    \CD[2].col_reg[1][5] ,
    \CD[2].col_reg[1][5]_0 ,
    \CD[0].col[3][5]_i_2_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][6] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][6] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][6] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][6] ,
    \CD[2].col_reg[1][6] ,
    \CD[2].col_reg[1][6]_0 ,
    \CD[0].col[3][6]_i_2_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][7] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][7] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][7] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][7] ,
    \CD[2].col_reg[1][7] ,
    \CD[2].col_reg[1][7]_0 ,
    \CD[0].col[3][7]_i_2_0 ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][8] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][8] ,
    \CD[1].col_reg[2][8] ,
    \CD[1].col_reg[2][8]_0 ,
    \CD[1].col_reg[2][8]_1 ,
    \IV_BKP_REGISTERS[3].bkp[3][8]_i_2 ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][9] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][9] ,
    \CD[1].col_reg[2][9] ,
    \CD[1].col_reg[2][9]_0 ,
    \CD[1].col_reg[2][9]_1 ,
    \IV_BKP_REGISTERS[3].bkp[3][9]_i_2 ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][10] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][10] ,
    \CD[1].col_reg[2][10] ,
    \CD[1].col_reg[2][10]_0 ,
    \CD[1].col_reg[2][10]_1 ,
    \CD[0].col[3][10]_i_3_0 ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][11] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][11] ,
    \CD[1].col_reg[2][11] ,
    \CD[1].col_reg[2][11]_0 ,
    \CD[1].col_reg[2][11]_1 ,
    \CD[0].col[3][11]_i_3_0 ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][12] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][12] ,
    \CD[1].col_reg[2][12] ,
    \CD[1].col_reg[2][12]_0 ,
    \CD[1].col_reg[2][12]_1 ,
    \CD[0].col[3][12]_i_3_0 ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][13] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][13] ,
    \CD[1].col_reg[2][13] ,
    \CD[1].col_reg[2][13]_0 ,
    \CD[1].col_reg[2][13]_1 ,
    \CD[0].col[3][13]_i_3_0 ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][14] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][14] ,
    \CD[1].col_reg[2][14] ,
    \CD[1].col_reg[2][14]_0 ,
    \CD[1].col_reg[2][14]_1 ,
    \IV_BKP_REGISTERS[3].bkp[3][14]_i_2 ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][15] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][15] ,
    \CD[1].col_reg[2][15] ,
    \CD[1].col_reg[2][15]_0 ,
    \CD[1].col_reg[2][15]_1 ,
    \IV_BKP_REGISTERS[3].bkp[3][15]_i_4 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][16] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][16] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][16] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][16] ,
    \CD[1].col_reg[2][16] ,
    \CD[1].col_reg[2][16]_0 ,
    \CD[0].col[3][16]_i_2_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][17] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][17] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][17] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][17] ,
    \CD[1].col_reg[2][17] ,
    \CD[1].col_reg[2][17]_0 ,
    \CD[0].col[3][17]_i_2_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][18] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][18] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][18] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][18] ,
    \CD[1].col_reg[2][18] ,
    \CD[1].col_reg[2][18]_0 ,
    \CD[0].col[3][18]_i_2_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][19] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][19] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][19] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][19] ,
    \CD[1].col_reg[2][19] ,
    \CD[1].col_reg[2][19]_0 ,
    \CD[0].col[3][19]_i_2_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][20] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][20] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][20] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][20] ,
    \CD[1].col_reg[2][20] ,
    \CD[1].col_reg[2][20]_0 ,
    \CD[0].col[3][20]_i_2_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][21] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][21] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][21] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][21] ,
    \CD[1].col_reg[2][21] ,
    \CD[1].col_reg[2][21]_0 ,
    \CD[0].col[3][21]_i_2_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][22] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][22] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][22] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][22] ,
    \CD[1].col_reg[2][22] ,
    \CD[1].col_reg[2][22]_0 ,
    \CD[0].col[3][22]_i_2_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][23] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][23] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][23] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][23] ,
    \CD[1].col_reg[2][23]_0 ,
    \CD[1].col_reg[2][23]_1 ,
    \CD[0].col[3][23]_i_2_0 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][24] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][24] ,
    \CD[2].col_reg[1][24] ,
    \CD[2].col_reg[1][24]_0 ,
    \CD[2].col_reg[1][24]_1 ,
    \IV_BKP_REGISTERS[2].bkp[2][24]_i_2 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][25] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][25] ,
    \CD[2].col_reg[1][25] ,
    \CD[2].col_reg[1][25]_0 ,
    \CD[2].col_reg[1][25]_1 ,
    \IV_BKP_REGISTERS[2].bkp[2][25]_i_2 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][26] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][26] ,
    \CD[2].col_reg[1][26] ,
    \CD[2].col_reg[1][26]_0 ,
    \CD[2].col_reg[1][26]_1 ,
    \IV_BKP_REGISTERS[2].bkp[2][26]_i_2 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][27] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][27] ,
    \CD[2].col_reg[1][27] ,
    \CD[2].col_reg[1][27]_0 ,
    \CD[2].col_reg[1][27]_1 ,
    \IV_BKP_REGISTERS[2].bkp[2][27]_i_2 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][28] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][28] ,
    \CD[2].col_reg[1][28] ,
    \CD[2].col_reg[1][28]_0 ,
    \CD[2].col_reg[1][28]_1 ,
    \CD[0].col[3][28]_i_2_0 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][29] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][29] ,
    \CD[2].col_reg[1][29] ,
    \CD[2].col_reg[1][29]_0 ,
    \CD[2].col_reg[1][29]_1 ,
    \IV_BKP_REGISTERS[2].bkp[2][29]_i_2 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][30] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][30] ,
    \CD[2].col_reg[1][30] ,
    \CD[2].col_reg[1][30]_0 ,
    \CD[2].col_reg[1][30]_1 ,
    \IV_BKP_REGISTERS[2].bkp[2][30]_i_2 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 ,
    \CD[2].col_reg[1][31]_2 ,
    \CD[2].col_reg[1][31]_3 ,
    \CD[2].col_reg[1][31]_4 ,
    \IV_BKP_REGISTERS[2].bkp[2][31]_i_2 ,
    \KR[2].key_reg[1][30] ,
    key_in,
    \KR[2].key_reg[1][28] ,
    g_func,
    \KR[2].key_reg[1][31]_0 ,
    \KR[2].key_reg[1][24] ,
    \KR[2].key_reg[1][29] ,
    \KR[2].key_reg[1][25] ,
    isomorphism_inv_return033_out,
    isomorphism_inv_return03_out,
    sbox_out_enc,
    isomorphism_inv_return05_out,
    p_86_in,
    p_93_in,
    p_16_in,
    isomorphism_inv_return033_out_6,
    isomorphism_inv_return03_out_7,
    isomorphism_inv_return05_out_8,
    p_86_in_9,
    p_93_in_10,
    p_16_in_11,
    isomorphism_inv_return033_out_12,
    isomorphism_inv_return03_out_13,
    isomorphism_inv_return05_out_14,
    p_86_in_15,
    p_93_in_16,
    p_16_in_17,
    \CD[0].col[3][31]_i_5_0 ,
    \CD[0].col[3][5]_i_2_1 ,
    \CD[0].col[3][5]_i_2_2 ,
    \CD[0].col[3][0]_i_2_0 ,
    \CD[0].col[3][1]_i_2_1 ,
    \CD[0].col[3][2]_i_2_1 ,
    \CD[0].col[3][3]_i_2_1 ,
    \CD[0].col[3][4]_i_2_1 ,
    \CD[0].col[3][6]_i_2_1 ,
    \CD[0].col[3][7]_i_2_1 ,
    \CD[0].col[3][8]_i_3_0 ,
    \CD[0].col[3][9]_i_3_0 ,
    \CD[0].col[3][31]_i_10_0 ,
    \CD[0].col[3][10]_i_6_0 ,
    \CD[0].col[3][14]_i_3_0 ,
    \CD[0].col[3][15]_i_5_0 ,
    \CD[0].col[3][16]_i_2_1 ,
    \CD[0].col[3][17]_i_2_1 ,
    \CD[0].col[3][18]_i_2_1 ,
    \CD[0].col[3][19]_i_2_1 ,
    \CD[0].col[3][20]_i_2_1 ,
    \CD[0].col[3][21]_i_2_1 ,
    \CD[0].col[3][22]_i_2_1 ,
    \CD[0].col[3][23]_i_2_1 ,
    \CD[0].col[3][24]_i_2_0 ,
    \CD[0].col[3][25]_i_2_0 ,
    \CD[0].col[3][26]_i_2_0 ,
    \CD[0].col[3][27]_i_2_0 ,
    \CD[0].col[3][29]_i_2_0 ,
    \CD[0].col[3][30]_i_2_0 ,
    \CD[0].col[3][31]_i_5_1 ,
    \CD[0].col[3][0]_i_4_0 ,
    first_block,
    \info_o[31]_3 ,
    \CD[0].col[3][31]_i_13_0 ,
    \CD[0].col[3][31]_i_13_1 ,
    \CD[0].col_reg[3][31]_1 ,
    col_en_host,
    \CD[0].col[3][31]_i_22 ,
    \CD[3].col_reg[0][31]_2 ,
    \CD[3].col_reg[0][31]_3 ,
    \CD[0].col[3][10]_i_12_0 ,
    \KR[0].key_reg[3][31] ,
    \KR[3].key_reg[0][31]_0 ,
    \info_o[31]_INST_0_i_4 ,
    \info_o[31]_INST_0_i_4_0 ,
    \info_o[31]_INST_0_i_4_1 ,
    key_sel_pp1,
    O,
    \IV_BKP_REGISTERS[3].iv_reg[3][24]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][16] ,
    \IV_BKP_REGISTERS[3].iv_reg[3][8]_0 ,
    rk_out_sel_pp2,
    \info_o[28]_INST_0_i_15 ,
    \info_o[28]_INST_0_i_15_0 ,
    \CD[0].col[3][31]_i_7_0 ,
    \info_o[31]_INST_0_i_12_0 ,
    enc_dec,
    \base_new_pp_reg[7] ,
    \base_new_pp_reg[7]_0 ,
    \base_new_pp_reg[7]_1 ,
    \out_gf_pp[1]_i_2 ,
    \base_new_pp_reg[7]_2 ,
    \base_new_pp_reg[7]_3 ,
    \base_new_pp_reg[7]_4 ,
    \out_gf_pp[1]_i_2__0 ,
    \base_new_pp_reg[7]_5 ,
    \base_new_pp_reg[7]_6 ,
    \base_new_pp_reg[7]_7 ,
    \out_gf_pp[1]_i_2__1 ,
    \base_new_pp_reg[7]_8 ,
    \base_new_pp_reg[7]_9 ,
    \base_new_pp_reg[7]_10 ,
    \out_gf_pp[1]_i_2__2 ,
    clk_i,
    rst_i,
    \FSM_sequential_state_reg[1]_1 );
  output [27:0]info_o;
  output \aes_cr_reg[7] ;
  output ccf_reg;
  output [3:0]Q;
  output \FSM_sequential_state_reg[2]_0 ;
  output \FSM_sequential_state_reg[3]_0 ;
  output \FSM_sequential_state_reg[2]_1 ;
  output \FSM_sequential_state_reg[0]_0 ;
  output [1:0]D;
  output \rd_count_reg[3]_0 ;
  output [3:0]\rd_count_reg[3]_1 ;
  output [1:0]\FSM_sequential_state_reg[1]_0 ;
  output [3:0]\FSM_sequential_state_reg[0]_1 ;
  output [3:0]\FSM_sequential_state_reg[2]_2 ;
  output key_sel;
  output \aes_cr_reg[4] ;
  output [1:0]\FSM_sequential_state_reg[2]_3 ;
  output \FSM_sequential_state_reg[3]_1 ;
  output \FSM_sequential_state_reg[3]_2 ;
  output \FSM_sequential_state_reg[2]_4 ;
  output bypass_key_en;
  output last_round;
  output \FSM_sequential_state_reg[2]_5 ;
  output key_sel_mux;
  output [23:0]\CD[3].col_reg[0][31] ;
  output [23:0]\CD[1].col_reg[2][23] ;
  output [23:0]\CD[2].col_reg[1][23] ;
  output [23:0]\CD[0].col_reg[3][31] ;
  output [31:0]\CD[3].col_reg[0][31]_0 ;
  output [31:0]\CD[0].col_reg[3][31]_0 ;
  output [31:0]\CD[1].col_reg[2][31] ;
  output [31:0]\CD[2].col_reg[1][31] ;
  output \FSM_sequential_state_reg[0]_2 ;
  output \IV_BKP_REGISTERS[2].iv_reg[2][8] ;
  output \IV_BKP_REGISTERS[2].iv_reg[2][9] ;
  output [4:0]data_in;
  output \IV_BKP_REGISTERS[2].iv_reg[2][14] ;
  output \IV_BKP_REGISTERS[2].iv_reg[2][15] ;
  output \IV_BKP_REGISTERS[2].iv_reg[2][24] ;
  output \IV_BKP_REGISTERS[2].iv_reg[2][25] ;
  output \IV_BKP_REGISTERS[2].iv_reg[2][26] ;
  output \IV_BKP_REGISTERS[2].iv_reg[2][27] ;
  output \IV_BKP_REGISTERS[2].iv_reg[2][29] ;
  output \IV_BKP_REGISTERS[2].iv_reg[2][30] ;
  output \IV_BKP_REGISTERS[2].iv_reg[2][31] ;
  output [31:0]\KR[3].key_reg[0][31] ;
  output \CD[3].col_reg[0][0] ;
  output \FSM_sequential_state_reg[2]_6 ;
  output \FSM_sequential_state_reg[3]_3 ;
  output \FSM_sequential_state_reg[3]_4 ;
  output \CD[3].col_reg[0][7] ;
  output \CD[3].col_reg[0][15] ;
  output \CD[3].col_reg[0][31]_1 ;
  output \CD[3].col_reg[0][1] ;
  output \CD[3].col_reg[0][6] ;
  output \CD[3].col_reg[0][14] ;
  output \CD[3].col_reg[0][30] ;
  output \CD[3].col_reg[0][2] ;
  output \CD[3].col_reg[0][5] ;
  output \CD[3].col_reg[0][13] ;
  output \CD[3].col_reg[0][29] ;
  output \CD[3].col_reg[0][3] ;
  output \CD[3].col_reg[0][4] ;
  output \CD[3].col_reg[0][12] ;
  output \CD[3].col_reg[0][28] ;
  output \CD[3].col_reg[0][11] ;
  output \CD[3].col_reg[0][27] ;
  output \CD[3].col_reg[0][10] ;
  output \CD[3].col_reg[0][26] ;
  output \CD[3].col_reg[0][9] ;
  output \CD[3].col_reg[0][25] ;
  output \CD[3].col_reg[0][8] ;
  output \CD[3].col_reg[0][24] ;
  output \CD[3].col_reg[0][23] ;
  output \CD[3].col_reg[0][22] ;
  output \CD[3].col_reg[0][21] ;
  output \CD[3].col_reg[0][20] ;
  output \CD[3].col_reg[0][19] ;
  output \CD[3].col_reg[0][18] ;
  output \CD[3].col_reg[0][17] ;
  output \CD[3].col_reg[0][16] ;
  output first_block_reg;
  output iv_mux_out13_out;
  output \col_en_cnt_unit_pp2_reg[3] ;
  output first_block_reg_0;
  output \IV_BKP_REGISTERS[3].iv_reg[3][8] ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][9] ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][14] ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][15] ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][24] ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][25] ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][26] ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][27] ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][29] ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][30] ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][31] ;
  output [0:0]E;
  output [0:0]\col_en_cnt_unit_pp2_reg[2] ;
  output [0:0]\col_en_cnt_unit_pp2_reg[1] ;
  output [0:0]\col_en_cnt_unit_pp2_reg[0] ;
  output enc_dec_sbox;
  output [0:0]\FSM_sequential_state_reg[3]_5 ;
  output [0:0]\FSM_sequential_state_reg[3]_6 ;
  output [0:0]\key_en_pp1_reg[3] ;
  output [0:0]\key_en_pp1_reg[2] ;
  output [0:0]\key_en_pp1_reg[1] ;
  output [0:0]\key_en_pp1_reg[0] ;
  output \aes_cr_reg[5] ;
  output \aes_cr_reg[5]_0 ;
  output \key_out_sel_pp1_reg[1] ;
  output [31:0]\enable_i[31] ;
  output add_rk_sel;
  output \FSM_sequential_state_reg[3]_7 ;
  output \FSM_sequential_state_reg[3]_8 ;
  output first_block_reg_1;
  output isomorphism_return179_out;
  output isomorphism_return114_out;
  output isomorphism_return179_out_0;
  output isomorphism_return114_out_1;
  output isomorphism_return179_out_2;
  output isomorphism_return114_out_3;
  output isomorphism_return179_out_4;
  output isomorphism_return114_out_5;
  input \info_o[31] ;
  input [21:0]key_out;
  input \info_o[31]_0 ;
  input info_o_0_sp_1;
  input [26:0]col_out;
  input info_o_4_sp_1;
  input info_o_6_sp_1;
  input info_o_9_sp_1;
  input info_o_10_sp_1;
  input info_o_11_sp_1;
  input info_o_12_sp_1;
  input \FSM_sequential_state_reg[0]_3 ;
  input \col_en_cnt_unit_pp1_reg[3] ;
  input \FSM_sequential_state_reg[2]_7 ;
  input [31:0]enable_i;
  input ccf;
  input ccf_reg_0;
  input \col_sel_pp1_reg[1] ;
  input [4:0]\info_o[0]_0 ;
  input \info_o[31]_1 ;
  input \key_en_pp1_reg[3]_0 ;
  input \FSM_sequential_state_reg[3]_9 ;
  input \FSM_sequential_state_reg[3]_10 ;
  input \FSM_sequential_state_reg[3]_11 ;
  input \FSM_sequential_state_reg[0]_4 ;
  input \FSM_sequential_state_reg[0]_5 ;
  input [3:0]key_en;
  input [31:0]\KR[2].key_reg[1][31] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][0] ;
  input [31:0]\CD[2].col_reg[1][31]_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][31] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][0] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][0] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][0] ;
  input [31:0]\CD[1].col_reg[2][31]_0 ;
  input [15:0]add_rk_out;
  input [31:0]\IV_BKP_REGISTERS[0].bkp_reg[0][31] ;
  input [31:0]\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 ;
  input \CD[2].col_reg[1][31]_1 ;
  input \CD[2].col_reg[1][0] ;
  input \CD[2].col_reg[1][0]_0 ;
  input [31:0]\info_o[31]_2 ;
  input [31:0]bus_swap;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][1] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][1] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][1] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][1] ;
  input \CD[2].col_reg[1][1] ;
  input \CD[2].col_reg[1][1]_0 ;
  input \CD[0].col[3][1]_i_2_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][2] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][2] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][2] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][2] ;
  input \CD[2].col_reg[1][2] ;
  input \CD[2].col_reg[1][2]_0 ;
  input \CD[0].col[3][2]_i_2_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][3] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][3] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][3] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][3] ;
  input \CD[2].col_reg[1][3] ;
  input \CD[2].col_reg[1][3]_0 ;
  input \CD[0].col[3][3]_i_2_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][4] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][4] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][4] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][4] ;
  input \CD[2].col_reg[1][4] ;
  input \CD[2].col_reg[1][4]_0 ;
  input \CD[0].col[3][4]_i_2_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][5] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][5] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][5] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][5] ;
  input \CD[2].col_reg[1][5] ;
  input \CD[2].col_reg[1][5]_0 ;
  input \CD[0].col[3][5]_i_2_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][6] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][6] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][6] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][6] ;
  input \CD[2].col_reg[1][6] ;
  input \CD[2].col_reg[1][6]_0 ;
  input \CD[0].col[3][6]_i_2_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][7] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][7] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][7] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][7] ;
  input \CD[2].col_reg[1][7] ;
  input \CD[2].col_reg[1][7]_0 ;
  input \CD[0].col[3][7]_i_2_0 ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][8] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][8] ;
  input \CD[1].col_reg[2][8] ;
  input \CD[1].col_reg[2][8]_0 ;
  input \CD[1].col_reg[2][8]_1 ;
  input \IV_BKP_REGISTERS[3].bkp[3][8]_i_2 ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][9] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][9] ;
  input \CD[1].col_reg[2][9] ;
  input \CD[1].col_reg[2][9]_0 ;
  input \CD[1].col_reg[2][9]_1 ;
  input \IV_BKP_REGISTERS[3].bkp[3][9]_i_2 ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][10] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][10] ;
  input \CD[1].col_reg[2][10] ;
  input \CD[1].col_reg[2][10]_0 ;
  input \CD[1].col_reg[2][10]_1 ;
  input \CD[0].col[3][10]_i_3_0 ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][11] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][11] ;
  input \CD[1].col_reg[2][11] ;
  input \CD[1].col_reg[2][11]_0 ;
  input \CD[1].col_reg[2][11]_1 ;
  input \CD[0].col[3][11]_i_3_0 ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][12] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][12] ;
  input \CD[1].col_reg[2][12] ;
  input \CD[1].col_reg[2][12]_0 ;
  input \CD[1].col_reg[2][12]_1 ;
  input \CD[0].col[3][12]_i_3_0 ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][13] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][13] ;
  input \CD[1].col_reg[2][13] ;
  input \CD[1].col_reg[2][13]_0 ;
  input \CD[1].col_reg[2][13]_1 ;
  input \CD[0].col[3][13]_i_3_0 ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][14] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][14] ;
  input \CD[1].col_reg[2][14] ;
  input \CD[1].col_reg[2][14]_0 ;
  input \CD[1].col_reg[2][14]_1 ;
  input \IV_BKP_REGISTERS[3].bkp[3][14]_i_2 ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][15] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][15] ;
  input \CD[1].col_reg[2][15] ;
  input \CD[1].col_reg[2][15]_0 ;
  input \CD[1].col_reg[2][15]_1 ;
  input \IV_BKP_REGISTERS[3].bkp[3][15]_i_4 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][16] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][16] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][16] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][16] ;
  input \CD[1].col_reg[2][16] ;
  input \CD[1].col_reg[2][16]_0 ;
  input \CD[0].col[3][16]_i_2_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][17] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][17] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][17] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][17] ;
  input \CD[1].col_reg[2][17] ;
  input \CD[1].col_reg[2][17]_0 ;
  input \CD[0].col[3][17]_i_2_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][18] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][18] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][18] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][18] ;
  input \CD[1].col_reg[2][18] ;
  input \CD[1].col_reg[2][18]_0 ;
  input \CD[0].col[3][18]_i_2_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][19] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][19] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][19] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][19] ;
  input \CD[1].col_reg[2][19] ;
  input \CD[1].col_reg[2][19]_0 ;
  input \CD[0].col[3][19]_i_2_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][20] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][20] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][20] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][20] ;
  input \CD[1].col_reg[2][20] ;
  input \CD[1].col_reg[2][20]_0 ;
  input \CD[0].col[3][20]_i_2_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][21] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][21] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][21] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][21] ;
  input \CD[1].col_reg[2][21] ;
  input \CD[1].col_reg[2][21]_0 ;
  input \CD[0].col[3][21]_i_2_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][22] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][22] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][22] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][22] ;
  input \CD[1].col_reg[2][22] ;
  input \CD[1].col_reg[2][22]_0 ;
  input \CD[0].col[3][22]_i_2_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][23] ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][23] ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][23] ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][23] ;
  input \CD[1].col_reg[2][23]_0 ;
  input \CD[1].col_reg[2][23]_1 ;
  input \CD[0].col[3][23]_i_2_0 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][24] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][24] ;
  input \CD[2].col_reg[1][24] ;
  input \CD[2].col_reg[1][24]_0 ;
  input \CD[2].col_reg[1][24]_1 ;
  input \IV_BKP_REGISTERS[2].bkp[2][24]_i_2 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][25] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][25] ;
  input \CD[2].col_reg[1][25] ;
  input \CD[2].col_reg[1][25]_0 ;
  input \CD[2].col_reg[1][25]_1 ;
  input \IV_BKP_REGISTERS[2].bkp[2][25]_i_2 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][26] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][26] ;
  input \CD[2].col_reg[1][26] ;
  input \CD[2].col_reg[1][26]_0 ;
  input \CD[2].col_reg[1][26]_1 ;
  input \IV_BKP_REGISTERS[2].bkp[2][26]_i_2 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][27] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][27] ;
  input \CD[2].col_reg[1][27] ;
  input \CD[2].col_reg[1][27]_0 ;
  input \CD[2].col_reg[1][27]_1 ;
  input \IV_BKP_REGISTERS[2].bkp[2][27]_i_2 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][28] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][28] ;
  input \CD[2].col_reg[1][28] ;
  input \CD[2].col_reg[1][28]_0 ;
  input \CD[2].col_reg[1][28]_1 ;
  input \CD[0].col[3][28]_i_2_0 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][29] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][29] ;
  input \CD[2].col_reg[1][29] ;
  input \CD[2].col_reg[1][29]_0 ;
  input \CD[2].col_reg[1][29]_1 ;
  input \IV_BKP_REGISTERS[2].bkp[2][29]_i_2 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][30] ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][30] ;
  input \CD[2].col_reg[1][30] ;
  input \CD[2].col_reg[1][30]_0 ;
  input \CD[2].col_reg[1][30]_1 ;
  input \IV_BKP_REGISTERS[2].bkp[2][30]_i_2 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 ;
  input \CD[2].col_reg[1][31]_2 ;
  input \CD[2].col_reg[1][31]_3 ;
  input \CD[2].col_reg[1][31]_4 ;
  input \IV_BKP_REGISTERS[2].bkp[2][31]_i_2 ;
  input \KR[2].key_reg[1][30] ;
  input [127:0]key_in;
  input \KR[2].key_reg[1][28] ;
  input [1:0]g_func;
  input \KR[2].key_reg[1][31]_0 ;
  input \KR[2].key_reg[1][24] ;
  input \KR[2].key_reg[1][29] ;
  input \KR[2].key_reg[1][25] ;
  input isomorphism_inv_return033_out;
  input isomorphism_inv_return03_out;
  input [5:0]sbox_out_enc;
  input isomorphism_inv_return05_out;
  input p_86_in;
  input p_93_in;
  input p_16_in;
  input isomorphism_inv_return033_out_6;
  input isomorphism_inv_return03_out_7;
  input isomorphism_inv_return05_out_8;
  input p_86_in_9;
  input p_93_in_10;
  input p_16_in_11;
  input isomorphism_inv_return033_out_12;
  input isomorphism_inv_return03_out_13;
  input isomorphism_inv_return05_out_14;
  input p_86_in_15;
  input p_93_in_16;
  input p_16_in_17;
  input [31:0]\CD[0].col[3][31]_i_5_0 ;
  input \CD[0].col[3][5]_i_2_1 ;
  input \CD[0].col[3][5]_i_2_2 ;
  input \CD[0].col[3][0]_i_2_0 ;
  input \CD[0].col[3][1]_i_2_1 ;
  input \CD[0].col[3][2]_i_2_1 ;
  input \CD[0].col[3][3]_i_2_1 ;
  input \CD[0].col[3][4]_i_2_1 ;
  input \CD[0].col[3][6]_i_2_1 ;
  input \CD[0].col[3][7]_i_2_1 ;
  input \CD[0].col[3][8]_i_3_0 ;
  input \CD[0].col[3][9]_i_3_0 ;
  input [31:0]\CD[0].col[3][31]_i_10_0 ;
  input \CD[0].col[3][10]_i_6_0 ;
  input \CD[0].col[3][14]_i_3_0 ;
  input \CD[0].col[3][15]_i_5_0 ;
  input \CD[0].col[3][16]_i_2_1 ;
  input \CD[0].col[3][17]_i_2_1 ;
  input \CD[0].col[3][18]_i_2_1 ;
  input \CD[0].col[3][19]_i_2_1 ;
  input \CD[0].col[3][20]_i_2_1 ;
  input \CD[0].col[3][21]_i_2_1 ;
  input \CD[0].col[3][22]_i_2_1 ;
  input \CD[0].col[3][23]_i_2_1 ;
  input \CD[0].col[3][24]_i_2_0 ;
  input \CD[0].col[3][25]_i_2_0 ;
  input \CD[0].col[3][26]_i_2_0 ;
  input \CD[0].col[3][27]_i_2_0 ;
  input \CD[0].col[3][29]_i_2_0 ;
  input \CD[0].col[3][30]_i_2_0 ;
  input \CD[0].col[3][31]_i_5_1 ;
  input \CD[0].col[3][0]_i_4_0 ;
  input first_block;
  input [27:0]\info_o[31]_3 ;
  input [31:0]\CD[0].col[3][31]_i_13_0 ;
  input [31:0]\CD[0].col[3][31]_i_13_1 ;
  input [3:0]\CD[0].col_reg[3][31]_1 ;
  input [3:0]col_en_host;
  input \CD[0].col[3][31]_i_22 ;
  input [1:0]\CD[3].col_reg[0][31]_2 ;
  input \CD[3].col_reg[0][31]_3 ;
  input \CD[0].col[3][10]_i_12_0 ;
  input [3:0]\KR[0].key_reg[3][31] ;
  input \KR[3].key_reg[0][31]_0 ;
  input [0:0]\info_o[31]_INST_0_i_4 ;
  input \info_o[31]_INST_0_i_4_0 ;
  input [0:0]\info_o[31]_INST_0_i_4_1 ;
  input key_sel_pp1;
  input [6:0]O;
  input [7:0]\IV_BKP_REGISTERS[3].iv_reg[3][24]_0 ;
  input [7:0]\IV_BKP_REGISTERS[3].iv_reg[3][16] ;
  input [7:0]\IV_BKP_REGISTERS[3].iv_reg[3][8]_0 ;
  input rk_out_sel_pp2;
  input \info_o[28]_INST_0_i_15 ;
  input \info_o[28]_INST_0_i_15_0 ;
  input [1:0]\CD[0].col[3][31]_i_7_0 ;
  input \info_o[31]_INST_0_i_12_0 ;
  input enc_dec;
  input \base_new_pp_reg[7] ;
  input \base_new_pp_reg[7]_0 ;
  input \base_new_pp_reg[7]_1 ;
  input \out_gf_pp[1]_i_2 ;
  input \base_new_pp_reg[7]_2 ;
  input \base_new_pp_reg[7]_3 ;
  input \base_new_pp_reg[7]_4 ;
  input \out_gf_pp[1]_i_2__0 ;
  input \base_new_pp_reg[7]_5 ;
  input \base_new_pp_reg[7]_6 ;
  input \base_new_pp_reg[7]_7 ;
  input \out_gf_pp[1]_i_2__1 ;
  input \base_new_pp_reg[7]_8 ;
  input \base_new_pp_reg[7]_9 ;
  input \base_new_pp_reg[7]_10 ;
  input \out_gf_pp[1]_i_2__2 ;
  input clk_i;
  input rst_i;
  input [0:0]\FSM_sequential_state_reg[1]_1 ;

  wire [1:0]\AES_CORE_DATAPATH/col_sel_w_bypass ;
  wire [31:0]\AES_CORE_DATAPATH/g_in ;
  wire \AES_CORE_DATAPATH/iv_mux_out1 ;
  wire \AES_CORE_DATAPATH/iv_mux_out10_out ;
  wire \AES_CORE_DATAPATH/key1_mux_cnt ;
  wire \CD[0].col[3][0]_i_10_n_0 ;
  wire \CD[0].col[3][0]_i_13_n_0 ;
  wire \CD[0].col[3][0]_i_14_n_0 ;
  wire \CD[0].col[3][0]_i_2_0 ;
  wire \CD[0].col[3][0]_i_2_n_0 ;
  wire \CD[0].col[3][0]_i_4_0 ;
  wire \CD[0].col[3][0]_i_4_n_0 ;
  wire \CD[0].col[3][0]_i_7_n_0 ;
  wire \CD[0].col[3][10]_i_12_0 ;
  wire \CD[0].col[3][10]_i_12_n_0 ;
  wire \CD[0].col[3][10]_i_3_0 ;
  wire \CD[0].col[3][10]_i_3_n_0 ;
  wire \CD[0].col[3][10]_i_6_0 ;
  wire \CD[0].col[3][10]_i_6_n_0 ;
  wire \CD[0].col[3][10]_i_9_n_0 ;
  wire \CD[0].col[3][11]_i_13_n_0 ;
  wire \CD[0].col[3][11]_i_3_0 ;
  wire \CD[0].col[3][11]_i_3_n_0 ;
  wire \CD[0].col[3][11]_i_6_n_0 ;
  wire \CD[0].col[3][11]_i_9_n_0 ;
  wire \CD[0].col[3][12]_i_14_n_0 ;
  wire \CD[0].col[3][12]_i_3_0 ;
  wire \CD[0].col[3][12]_i_3_n_0 ;
  wire \CD[0].col[3][12]_i_6_n_0 ;
  wire \CD[0].col[3][12]_i_9_n_0 ;
  wire \CD[0].col[3][13]_i_11_n_0 ;
  wire \CD[0].col[3][13]_i_3_0 ;
  wire \CD[0].col[3][13]_i_3_n_0 ;
  wire \CD[0].col[3][13]_i_6_n_0 ;
  wire \CD[0].col[3][13]_i_9_n_0 ;
  wire \CD[0].col[3][14]_i_11_n_0 ;
  wire \CD[0].col[3][14]_i_15_n_0 ;
  wire \CD[0].col[3][14]_i_3_0 ;
  wire \CD[0].col[3][14]_i_3_n_0 ;
  wire \CD[0].col[3][14]_i_6_n_0 ;
  wire \CD[0].col[3][15]_i_16_n_0 ;
  wire \CD[0].col[3][15]_i_20_n_0 ;
  wire \CD[0].col[3][15]_i_3_n_0 ;
  wire \CD[0].col[3][15]_i_5_0 ;
  wire \CD[0].col[3][15]_i_5_n_0 ;
  wire \CD[0].col[3][15]_i_9_n_0 ;
  wire \CD[0].col[3][16]_i_12_n_0 ;
  wire \CD[0].col[3][16]_i_2_0 ;
  wire \CD[0].col[3][16]_i_2_1 ;
  wire \CD[0].col[3][16]_i_2_n_0 ;
  wire \CD[0].col[3][16]_i_3_n_0 ;
  wire \CD[0].col[3][16]_i_4_n_0 ;
  wire \CD[0].col[3][16]_i_7_n_0 ;
  wire \CD[0].col[3][16]_i_8_n_0 ;
  wire \CD[0].col[3][17]_i_12_n_0 ;
  wire \CD[0].col[3][17]_i_2_0 ;
  wire \CD[0].col[3][17]_i_2_1 ;
  wire \CD[0].col[3][17]_i_2_n_0 ;
  wire \CD[0].col[3][17]_i_3_n_0 ;
  wire \CD[0].col[3][17]_i_4_n_0 ;
  wire \CD[0].col[3][17]_i_7_n_0 ;
  wire \CD[0].col[3][17]_i_8_n_0 ;
  wire \CD[0].col[3][18]_i_12_n_0 ;
  wire \CD[0].col[3][18]_i_2_0 ;
  wire \CD[0].col[3][18]_i_2_1 ;
  wire \CD[0].col[3][18]_i_2_n_0 ;
  wire \CD[0].col[3][18]_i_3_n_0 ;
  wire \CD[0].col[3][18]_i_4_n_0 ;
  wire \CD[0].col[3][18]_i_7_n_0 ;
  wire \CD[0].col[3][18]_i_8_n_0 ;
  wire \CD[0].col[3][19]_i_12_n_0 ;
  wire \CD[0].col[3][19]_i_2_0 ;
  wire \CD[0].col[3][19]_i_2_1 ;
  wire \CD[0].col[3][19]_i_2_n_0 ;
  wire \CD[0].col[3][19]_i_3_n_0 ;
  wire \CD[0].col[3][19]_i_4_n_0 ;
  wire \CD[0].col[3][19]_i_7_n_0 ;
  wire \CD[0].col[3][19]_i_8_n_0 ;
  wire \CD[0].col[3][1]_i_10_n_0 ;
  wire \CD[0].col[3][1]_i_12_n_0 ;
  wire \CD[0].col[3][1]_i_15_n_0 ;
  wire \CD[0].col[3][1]_i_2_0 ;
  wire \CD[0].col[3][1]_i_2_1 ;
  wire \CD[0].col[3][1]_i_2_n_0 ;
  wire \CD[0].col[3][1]_i_4_n_0 ;
  wire \CD[0].col[3][1]_i_7_n_0 ;
  wire \CD[0].col[3][20]_i_12_n_0 ;
  wire \CD[0].col[3][20]_i_2_0 ;
  wire \CD[0].col[3][20]_i_2_1 ;
  wire \CD[0].col[3][20]_i_2_n_0 ;
  wire \CD[0].col[3][20]_i_3_n_0 ;
  wire \CD[0].col[3][20]_i_4_n_0 ;
  wire \CD[0].col[3][20]_i_7_n_0 ;
  wire \CD[0].col[3][20]_i_8_n_0 ;
  wire \CD[0].col[3][21]_i_12_n_0 ;
  wire \CD[0].col[3][21]_i_2_0 ;
  wire \CD[0].col[3][21]_i_2_1 ;
  wire \CD[0].col[3][21]_i_2_n_0 ;
  wire \CD[0].col[3][21]_i_3_n_0 ;
  wire \CD[0].col[3][21]_i_4_n_0 ;
  wire \CD[0].col[3][21]_i_7_n_0 ;
  wire \CD[0].col[3][21]_i_8_n_0 ;
  wire \CD[0].col[3][22]_i_12_n_0 ;
  wire \CD[0].col[3][22]_i_2_0 ;
  wire \CD[0].col[3][22]_i_2_1 ;
  wire \CD[0].col[3][22]_i_2_n_0 ;
  wire \CD[0].col[3][22]_i_3_n_0 ;
  wire \CD[0].col[3][22]_i_4_n_0 ;
  wire \CD[0].col[3][22]_i_7_n_0 ;
  wire \CD[0].col[3][22]_i_8_n_0 ;
  wire \CD[0].col[3][23]_i_13_n_0 ;
  wire \CD[0].col[3][23]_i_2_0 ;
  wire \CD[0].col[3][23]_i_2_1 ;
  wire \CD[0].col[3][23]_i_2_n_0 ;
  wire \CD[0].col[3][23]_i_3_n_0 ;
  wire \CD[0].col[3][23]_i_4_n_0 ;
  wire \CD[0].col[3][23]_i_5_n_0 ;
  wire \CD[0].col[3][23]_i_8_n_0 ;
  wire \CD[0].col[3][23]_i_9_n_0 ;
  wire \CD[0].col[3][24]_i_10_n_0 ;
  wire \CD[0].col[3][24]_i_14_n_0 ;
  wire \CD[0].col[3][24]_i_2_0 ;
  wire \CD[0].col[3][24]_i_2_n_0 ;
  wire \CD[0].col[3][24]_i_4_n_0 ;
  wire \CD[0].col[3][25]_i_10_n_0 ;
  wire \CD[0].col[3][25]_i_14_n_0 ;
  wire \CD[0].col[3][25]_i_2_0 ;
  wire \CD[0].col[3][25]_i_2_n_0 ;
  wire \CD[0].col[3][25]_i_4_n_0 ;
  wire \CD[0].col[3][26]_i_10_n_0 ;
  wire \CD[0].col[3][26]_i_14_n_0 ;
  wire \CD[0].col[3][26]_i_2_0 ;
  wire \CD[0].col[3][26]_i_2_n_0 ;
  wire \CD[0].col[3][26]_i_4_n_0 ;
  wire \CD[0].col[3][27]_i_10_n_0 ;
  wire \CD[0].col[3][27]_i_14_n_0 ;
  wire \CD[0].col[3][27]_i_2_0 ;
  wire \CD[0].col[3][27]_i_2_n_0 ;
  wire \CD[0].col[3][27]_i_4_n_0 ;
  wire \CD[0].col[3][28]_i_10_n_0 ;
  wire \CD[0].col[3][28]_i_2_0 ;
  wire \CD[0].col[3][28]_i_2_n_0 ;
  wire \CD[0].col[3][28]_i_4_n_0 ;
  wire \CD[0].col[3][28]_i_7_n_0 ;
  wire \CD[0].col[3][29]_i_10_n_0 ;
  wire \CD[0].col[3][29]_i_14_n_0 ;
  wire \CD[0].col[3][29]_i_2_0 ;
  wire \CD[0].col[3][29]_i_2_n_0 ;
  wire \CD[0].col[3][29]_i_4_n_0 ;
  wire \CD[0].col[3][2]_i_10_n_0 ;
  wire \CD[0].col[3][2]_i_12_n_0 ;
  wire \CD[0].col[3][2]_i_15_n_0 ;
  wire \CD[0].col[3][2]_i_2_0 ;
  wire \CD[0].col[3][2]_i_2_1 ;
  wire \CD[0].col[3][2]_i_2_n_0 ;
  wire \CD[0].col[3][2]_i_4_n_0 ;
  wire \CD[0].col[3][2]_i_7_n_0 ;
  wire \CD[0].col[3][30]_i_10_n_0 ;
  wire \CD[0].col[3][30]_i_14_n_0 ;
  wire \CD[0].col[3][30]_i_2_0 ;
  wire \CD[0].col[3][30]_i_2_n_0 ;
  wire \CD[0].col[3][30]_i_4_n_0 ;
  wire [31:0]\CD[0].col[3][31]_i_10_0 ;
  wire \CD[0].col[3][31]_i_10_n_0 ;
  wire [31:0]\CD[0].col[3][31]_i_13_0 ;
  wire [31:0]\CD[0].col[3][31]_i_13_1 ;
  wire \CD[0].col[3][31]_i_18_n_0 ;
  wire \CD[0].col[3][31]_i_22 ;
  wire \CD[0].col[3][31]_i_27_n_0 ;
  wire \CD[0].col[3][31]_i_28_n_0 ;
  wire \CD[0].col[3][31]_i_4_n_0 ;
  wire [31:0]\CD[0].col[3][31]_i_5_0 ;
  wire \CD[0].col[3][31]_i_5_1 ;
  wire \CD[0].col[3][31]_i_5_n_0 ;
  wire [1:0]\CD[0].col[3][31]_i_7_0 ;
  wire \CD[0].col[3][31]_i_7_n_0 ;
  wire \CD[0].col[3][31]_i_8_n_0 ;
  wire \CD[0].col[3][3]_i_10_n_0 ;
  wire \CD[0].col[3][3]_i_12_n_0 ;
  wire \CD[0].col[3][3]_i_15_n_0 ;
  wire \CD[0].col[3][3]_i_2_0 ;
  wire \CD[0].col[3][3]_i_2_1 ;
  wire \CD[0].col[3][3]_i_2_n_0 ;
  wire \CD[0].col[3][3]_i_4_n_0 ;
  wire \CD[0].col[3][3]_i_7_n_0 ;
  wire \CD[0].col[3][4]_i_10_n_0 ;
  wire \CD[0].col[3][4]_i_14_n_0 ;
  wire \CD[0].col[3][4]_i_2_0 ;
  wire \CD[0].col[3][4]_i_2_1 ;
  wire \CD[0].col[3][4]_i_2_n_0 ;
  wire \CD[0].col[3][4]_i_4_n_0 ;
  wire \CD[0].col[3][4]_i_7_n_0 ;
  wire \CD[0].col[3][5]_i_10_n_0 ;
  wire \CD[0].col[3][5]_i_12_n_0 ;
  wire \CD[0].col[3][5]_i_15_n_0 ;
  wire \CD[0].col[3][5]_i_2_0 ;
  wire \CD[0].col[3][5]_i_2_1 ;
  wire \CD[0].col[3][5]_i_2_2 ;
  wire \CD[0].col[3][5]_i_2_n_0 ;
  wire \CD[0].col[3][5]_i_4_n_0 ;
  wire \CD[0].col[3][5]_i_7_n_0 ;
  wire \CD[0].col[3][6]_i_10_n_0 ;
  wire \CD[0].col[3][6]_i_14_n_0 ;
  wire \CD[0].col[3][6]_i_2_0 ;
  wire \CD[0].col[3][6]_i_2_1 ;
  wire \CD[0].col[3][6]_i_2_n_0 ;
  wire \CD[0].col[3][6]_i_4_n_0 ;
  wire \CD[0].col[3][6]_i_7_n_0 ;
  wire \CD[0].col[3][7]_i_11_n_0 ;
  wire \CD[0].col[3][7]_i_15_n_0 ;
  wire \CD[0].col[3][7]_i_2_0 ;
  wire \CD[0].col[3][7]_i_2_1 ;
  wire \CD[0].col[3][7]_i_2_n_0 ;
  wire \CD[0].col[3][7]_i_4_n_0 ;
  wire \CD[0].col[3][7]_i_5_n_0 ;
  wire \CD[0].col[3][7]_i_8_n_0 ;
  wire \CD[0].col[3][8]_i_12_n_0 ;
  wire \CD[0].col[3][8]_i_16_n_0 ;
  wire \CD[0].col[3][8]_i_3_0 ;
  wire \CD[0].col[3][8]_i_3_n_0 ;
  wire \CD[0].col[3][8]_i_6_n_0 ;
  wire \CD[0].col[3][9]_i_11_n_0 ;
  wire \CD[0].col[3][9]_i_15_n_0 ;
  wire \CD[0].col[3][9]_i_3_0 ;
  wire \CD[0].col[3][9]_i_3_n_0 ;
  wire \CD[0].col[3][9]_i_6_n_0 ;
  wire [23:0]\CD[0].col_reg[3][31] ;
  wire [31:0]\CD[0].col_reg[3][31]_0 ;
  wire [3:0]\CD[0].col_reg[3][31]_1 ;
  wire \CD[1].col[2][0]_i_2_n_0 ;
  wire \CD[1].col[2][1]_i_2_n_0 ;
  wire \CD[1].col[2][2]_i_2_n_0 ;
  wire \CD[1].col[2][3]_i_2_n_0 ;
  wire \CD[1].col[2][4]_i_2_n_0 ;
  wire \CD[1].col[2][5]_i_2_n_0 ;
  wire \CD[1].col[2][6]_i_2_n_0 ;
  wire \CD[1].col[2][7]_i_2_n_0 ;
  wire \CD[1].col_reg[2][10] ;
  wire \CD[1].col_reg[2][10]_0 ;
  wire \CD[1].col_reg[2][10]_1 ;
  wire \CD[1].col_reg[2][11] ;
  wire \CD[1].col_reg[2][11]_0 ;
  wire \CD[1].col_reg[2][11]_1 ;
  wire \CD[1].col_reg[2][12] ;
  wire \CD[1].col_reg[2][12]_0 ;
  wire \CD[1].col_reg[2][12]_1 ;
  wire \CD[1].col_reg[2][13] ;
  wire \CD[1].col_reg[2][13]_0 ;
  wire \CD[1].col_reg[2][13]_1 ;
  wire \CD[1].col_reg[2][14] ;
  wire \CD[1].col_reg[2][14]_0 ;
  wire \CD[1].col_reg[2][14]_1 ;
  wire \CD[1].col_reg[2][15] ;
  wire \CD[1].col_reg[2][15]_0 ;
  wire \CD[1].col_reg[2][15]_1 ;
  wire \CD[1].col_reg[2][16] ;
  wire \CD[1].col_reg[2][16]_0 ;
  wire \CD[1].col_reg[2][17] ;
  wire \CD[1].col_reg[2][17]_0 ;
  wire \CD[1].col_reg[2][18] ;
  wire \CD[1].col_reg[2][18]_0 ;
  wire \CD[1].col_reg[2][19] ;
  wire \CD[1].col_reg[2][19]_0 ;
  wire \CD[1].col_reg[2][20] ;
  wire \CD[1].col_reg[2][20]_0 ;
  wire \CD[1].col_reg[2][21] ;
  wire \CD[1].col_reg[2][21]_0 ;
  wire \CD[1].col_reg[2][22] ;
  wire \CD[1].col_reg[2][22]_0 ;
  wire [23:0]\CD[1].col_reg[2][23] ;
  wire \CD[1].col_reg[2][23]_0 ;
  wire \CD[1].col_reg[2][23]_1 ;
  wire [31:0]\CD[1].col_reg[2][31] ;
  wire [31:0]\CD[1].col_reg[2][31]_0 ;
  wire \CD[1].col_reg[2][8] ;
  wire \CD[1].col_reg[2][8]_0 ;
  wire \CD[1].col_reg[2][8]_1 ;
  wire \CD[1].col_reg[2][9] ;
  wire \CD[1].col_reg[2][9]_0 ;
  wire \CD[1].col_reg[2][9]_1 ;
  wire \CD[2].col_reg[1][0] ;
  wire \CD[2].col_reg[1][0]_0 ;
  wire \CD[2].col_reg[1][1] ;
  wire \CD[2].col_reg[1][1]_0 ;
  wire [23:0]\CD[2].col_reg[1][23] ;
  wire \CD[2].col_reg[1][24] ;
  wire \CD[2].col_reg[1][24]_0 ;
  wire \CD[2].col_reg[1][24]_1 ;
  wire \CD[2].col_reg[1][25] ;
  wire \CD[2].col_reg[1][25]_0 ;
  wire \CD[2].col_reg[1][25]_1 ;
  wire \CD[2].col_reg[1][26] ;
  wire \CD[2].col_reg[1][26]_0 ;
  wire \CD[2].col_reg[1][26]_1 ;
  wire \CD[2].col_reg[1][27] ;
  wire \CD[2].col_reg[1][27]_0 ;
  wire \CD[2].col_reg[1][27]_1 ;
  wire \CD[2].col_reg[1][28] ;
  wire \CD[2].col_reg[1][28]_0 ;
  wire \CD[2].col_reg[1][28]_1 ;
  wire \CD[2].col_reg[1][29] ;
  wire \CD[2].col_reg[1][29]_0 ;
  wire \CD[2].col_reg[1][29]_1 ;
  wire \CD[2].col_reg[1][2] ;
  wire \CD[2].col_reg[1][2]_0 ;
  wire \CD[2].col_reg[1][30] ;
  wire \CD[2].col_reg[1][30]_0 ;
  wire \CD[2].col_reg[1][30]_1 ;
  wire [31:0]\CD[2].col_reg[1][31] ;
  wire [31:0]\CD[2].col_reg[1][31]_0 ;
  wire \CD[2].col_reg[1][31]_1 ;
  wire \CD[2].col_reg[1][31]_2 ;
  wire \CD[2].col_reg[1][31]_3 ;
  wire \CD[2].col_reg[1][31]_4 ;
  wire \CD[2].col_reg[1][3] ;
  wire \CD[2].col_reg[1][3]_0 ;
  wire \CD[2].col_reg[1][4] ;
  wire \CD[2].col_reg[1][4]_0 ;
  wire \CD[2].col_reg[1][5] ;
  wire \CD[2].col_reg[1][5]_0 ;
  wire \CD[2].col_reg[1][6] ;
  wire \CD[2].col_reg[1][6]_0 ;
  wire \CD[2].col_reg[1][7] ;
  wire \CD[2].col_reg[1][7]_0 ;
  wire \CD[3].col_reg[0][0] ;
  wire \CD[3].col_reg[0][10] ;
  wire \CD[3].col_reg[0][11] ;
  wire \CD[3].col_reg[0][12] ;
  wire \CD[3].col_reg[0][13] ;
  wire \CD[3].col_reg[0][14] ;
  wire \CD[3].col_reg[0][15] ;
  wire \CD[3].col_reg[0][16] ;
  wire \CD[3].col_reg[0][17] ;
  wire \CD[3].col_reg[0][18] ;
  wire \CD[3].col_reg[0][19] ;
  wire \CD[3].col_reg[0][1] ;
  wire \CD[3].col_reg[0][20] ;
  wire \CD[3].col_reg[0][21] ;
  wire \CD[3].col_reg[0][22] ;
  wire \CD[3].col_reg[0][23] ;
  wire \CD[3].col_reg[0][24] ;
  wire \CD[3].col_reg[0][25] ;
  wire \CD[3].col_reg[0][26] ;
  wire \CD[3].col_reg[0][27] ;
  wire \CD[3].col_reg[0][28] ;
  wire \CD[3].col_reg[0][29] ;
  wire \CD[3].col_reg[0][2] ;
  wire \CD[3].col_reg[0][30] ;
  wire [23:0]\CD[3].col_reg[0][31] ;
  wire [31:0]\CD[3].col_reg[0][31]_0 ;
  wire \CD[3].col_reg[0][31]_1 ;
  wire [1:0]\CD[3].col_reg[0][31]_2 ;
  wire \CD[3].col_reg[0][31]_3 ;
  wire \CD[3].col_reg[0][3] ;
  wire \CD[3].col_reg[0][4] ;
  wire \CD[3].col_reg[0][5] ;
  wire \CD[3].col_reg[0][6] ;
  wire \CD[3].col_reg[0][7] ;
  wire \CD[3].col_reg[0][8] ;
  wire \CD[3].col_reg[0][9] ;
  wire [1:0]D;
  wire [0:0]E;
  wire \FSM_sequential_state[0]_i_1__0_n_0 ;
  wire \FSM_sequential_state[0]_i_2_n_0 ;
  wire \FSM_sequential_state[0]_i_3__0_n_0 ;
  wire \FSM_sequential_state[0]_i_5_n_0 ;
  wire \FSM_sequential_state[0]_i_6_n_0 ;
  wire \FSM_sequential_state[0]_i_7_n_0 ;
  wire \FSM_sequential_state[1]_i_8_n_0 ;
  wire \FSM_sequential_state[2]_i_1__0_n_0 ;
  wire \FSM_sequential_state[2]_i_2__0_n_0 ;
  wire \FSM_sequential_state[2]_i_3_n_0 ;
  wire \FSM_sequential_state[2]_i_5__0_n_0 ;
  wire \FSM_sequential_state[3]_i_1_n_0 ;
  wire \FSM_sequential_state[3]_i_2_n_0 ;
  wire \FSM_sequential_state[3]_i_4_n_0 ;
  wire \FSM_sequential_state[3]_i_5_n_0 ;
  wire \FSM_sequential_state_reg[0]_0 ;
  wire [3:0]\FSM_sequential_state_reg[0]_1 ;
  wire \FSM_sequential_state_reg[0]_2 ;
  wire \FSM_sequential_state_reg[0]_3 ;
  wire \FSM_sequential_state_reg[0]_4 ;
  wire \FSM_sequential_state_reg[0]_5 ;
  wire [1:0]\FSM_sequential_state_reg[1]_0 ;
  wire [0:0]\FSM_sequential_state_reg[1]_1 ;
  wire \FSM_sequential_state_reg[2]_0 ;
  wire \FSM_sequential_state_reg[2]_1 ;
  wire [3:0]\FSM_sequential_state_reg[2]_2 ;
  wire [1:0]\FSM_sequential_state_reg[2]_3 ;
  wire \FSM_sequential_state_reg[2]_4 ;
  wire \FSM_sequential_state_reg[2]_5 ;
  wire \FSM_sequential_state_reg[2]_6 ;
  wire \FSM_sequential_state_reg[2]_7 ;
  wire \FSM_sequential_state_reg[3]_0 ;
  wire \FSM_sequential_state_reg[3]_1 ;
  wire \FSM_sequential_state_reg[3]_10 ;
  wire \FSM_sequential_state_reg[3]_11 ;
  wire \FSM_sequential_state_reg[3]_2 ;
  wire \FSM_sequential_state_reg[3]_3 ;
  wire \FSM_sequential_state_reg[3]_4 ;
  wire [0:0]\FSM_sequential_state_reg[3]_5 ;
  wire [0:0]\FSM_sequential_state_reg[3]_6 ;
  wire \FSM_sequential_state_reg[3]_7 ;
  wire \FSM_sequential_state_reg[3]_8 ;
  wire \FSM_sequential_state_reg[3]_9 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][0]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][16]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][16]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][17]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][17]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][18]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][18]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][19]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][19]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][1]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][20]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][20]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][21]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][21]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][22]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][22]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][23]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][23]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][24]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][25]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][26]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][27]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][28]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][29]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][2]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][30]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][31]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][3]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][4]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][5]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][6]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][7]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][0] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][16] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][17] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][18] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][19] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][1] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][20] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][21] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][22] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][23] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][24] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][25] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][26] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][27] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][28] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][29] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][2] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][30] ;
  wire [31:0]\IV_BKP_REGISTERS[0].bkp_reg[0][31] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][3] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][4] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][5] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][6] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][7] ;
  wire \IV_BKP_REGISTERS[1].bkp[1][0]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][0]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][10]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][11]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][12]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][13]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][14]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][15]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][16]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][17]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][18]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][19]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][1]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][1]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][20]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][21]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][22]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][23]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][2]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][2]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][3]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][3]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][4]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][4]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][5]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][5]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][6]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][6]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][7]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][7]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][8]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][9]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][0] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][10] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][11] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][12] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][13] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][14] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][15] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][16] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][17] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][18] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][19] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][1] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][20] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][21] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][22] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][23] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][2] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][3] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][4] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][5] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][6] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][7] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][8] ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][9] ;
  wire \IV_BKP_REGISTERS[2].bkp[2][0]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][0]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][10]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][11]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][12]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][13]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][14]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][15]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][16]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][17]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][18]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][19]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][1]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][1]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][20]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][21]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][22]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][23]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][24]_i_2 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][25]_i_2 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][26]_i_2 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][27]_i_2 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][28]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][28]_i_6_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][29]_i_2 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][2]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][2]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][30]_i_2 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][31]_i_2 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][3]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][3]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][4]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][4]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][5]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][5]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][6]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][6]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][7]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][7]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][8]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][9]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][0] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][10] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][11] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][12] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][13] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][14] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][15] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][16] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][17] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][18] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][19] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][1] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][20] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][21] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][22] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][23] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][2] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][3] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][4] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][5] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][6] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][7] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][8] ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][9] ;
  wire \IV_BKP_REGISTERS[2].iv_reg[2][14] ;
  wire \IV_BKP_REGISTERS[2].iv_reg[2][15] ;
  wire \IV_BKP_REGISTERS[2].iv_reg[2][24] ;
  wire \IV_BKP_REGISTERS[2].iv_reg[2][25] ;
  wire \IV_BKP_REGISTERS[2].iv_reg[2][26] ;
  wire \IV_BKP_REGISTERS[2].iv_reg[2][27] ;
  wire \IV_BKP_REGISTERS[2].iv_reg[2][29] ;
  wire \IV_BKP_REGISTERS[2].iv_reg[2][30] ;
  wire \IV_BKP_REGISTERS[2].iv_reg[2][31] ;
  wire \IV_BKP_REGISTERS[2].iv_reg[2][8] ;
  wire \IV_BKP_REGISTERS[2].iv_reg[2][9] ;
  wire \IV_BKP_REGISTERS[3].bkp[3][0]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][10]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][10]_i_6_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][11]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][11]_i_6_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][12]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][12]_i_6_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][13]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][13]_i_6_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][14]_i_2 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][15]_i_4 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][16]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][16]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][17]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][17]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][18]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][18]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][19]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][19]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][1]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][20]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][20]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][21]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][21]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][22]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][22]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][23]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][23]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][24]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][25]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][26]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][27]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][28]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][29]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][2]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][30]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][31]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][3]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][4]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][5]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][6]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][7]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][8]_i_2 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][9]_i_2 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][0] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][16] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][17] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][18] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][19] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][1] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][20] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][21] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][22] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][23] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][24] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][25] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][26] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][27] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][28] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][29] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][2] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][30] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][31] ;
  wire [31:0]\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][3] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][4] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][5] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][6] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][7] ;
  wire \IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][14] ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][15] ;
  wire [7:0]\IV_BKP_REGISTERS[3].iv_reg[3][16] ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][24] ;
  wire [7:0]\IV_BKP_REGISTERS[3].iv_reg[3][24]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][25] ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][26] ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][27] ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][29] ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][30] ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][31] ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][8] ;
  wire [7:0]\IV_BKP_REGISTERS[3].iv_reg[3][8]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][9] ;
  wire [3:0]\KR[0].key_reg[3][31] ;
  wire \KR[2].key[1][0]_i_2_n_0 ;
  wire \KR[2].key[1][10]_i_2_n_0 ;
  wire \KR[2].key[1][11]_i_2_n_0 ;
  wire \KR[2].key[1][12]_i_2_n_0 ;
  wire \KR[2].key[1][13]_i_2_n_0 ;
  wire \KR[2].key[1][14]_i_2_n_0 ;
  wire \KR[2].key[1][15]_i_2_n_0 ;
  wire \KR[2].key[1][16]_i_2_n_0 ;
  wire \KR[2].key[1][17]_i_2_n_0 ;
  wire \KR[2].key[1][18]_i_2_n_0 ;
  wire \KR[2].key[1][19]_i_2_n_0 ;
  wire \KR[2].key[1][1]_i_2_n_0 ;
  wire \KR[2].key[1][20]_i_2_n_0 ;
  wire \KR[2].key[1][21]_i_2_n_0 ;
  wire \KR[2].key[1][22]_i_2_n_0 ;
  wire \KR[2].key[1][23]_i_2_n_0 ;
  wire \KR[2].key[1][24]_i_2_n_0 ;
  wire \KR[2].key[1][25]_i_2_n_0 ;
  wire \KR[2].key[1][26]_i_2_n_0 ;
  wire \KR[2].key[1][27]_i_2_n_0 ;
  wire \KR[2].key[1][28]_i_2_n_0 ;
  wire \KR[2].key[1][29]_i_2_n_0 ;
  wire \KR[2].key[1][2]_i_2_n_0 ;
  wire \KR[2].key[1][30]_i_2_n_0 ;
  wire \KR[2].key[1][31]_i_3_n_0 ;
  wire \KR[2].key[1][3]_i_2_n_0 ;
  wire \KR[2].key[1][4]_i_2_n_0 ;
  wire \KR[2].key[1][5]_i_2_n_0 ;
  wire \KR[2].key[1][6]_i_2_n_0 ;
  wire \KR[2].key[1][7]_i_2_n_0 ;
  wire \KR[2].key[1][8]_i_2_n_0 ;
  wire \KR[2].key[1][9]_i_2_n_0 ;
  wire \KR[2].key_reg[1][24] ;
  wire \KR[2].key_reg[1][25] ;
  wire \KR[2].key_reg[1][28] ;
  wire \KR[2].key_reg[1][29] ;
  wire \KR[2].key_reg[1][30] ;
  wire [31:0]\KR[2].key_reg[1][31] ;
  wire \KR[2].key_reg[1][31]_0 ;
  wire \KR[3].key[0][31]_i_4_n_0 ;
  wire [31:0]\KR[3].key_reg[0][31] ;
  wire \KR[3].key_reg[0][31]_0 ;
  wire [6:0]O;
  wire [3:0]Q;
  wire [15:0]add_rk_out;
  wire add_rk_sel;
  wire \aes_cr_reg[4] ;
  wire \aes_cr_reg[5] ;
  wire \aes_cr_reg[5]_0 ;
  wire \aes_cr_reg[7] ;
  wire \base_new_pp_reg[7] ;
  wire \base_new_pp_reg[7]_0 ;
  wire \base_new_pp_reg[7]_1 ;
  wire \base_new_pp_reg[7]_10 ;
  wire \base_new_pp_reg[7]_2 ;
  wire \base_new_pp_reg[7]_3 ;
  wire \base_new_pp_reg[7]_4 ;
  wire \base_new_pp_reg[7]_5 ;
  wire \base_new_pp_reg[7]_6 ;
  wire \base_new_pp_reg[7]_7 ;
  wire \base_new_pp_reg[7]_8 ;
  wire \base_new_pp_reg[7]_9 ;
  wire [31:0]bus_swap;
  wire bypass_key_en;
  wire ccf;
  wire ccf_reg;
  wire ccf_reg_0;
  wire clk_i;
  wire \col_en_cnt_unit_pp1_reg[3] ;
  wire [0:0]\col_en_cnt_unit_pp2_reg[0] ;
  wire [0:0]\col_en_cnt_unit_pp2_reg[1] ;
  wire [0:0]\col_en_cnt_unit_pp2_reg[2] ;
  wire \col_en_cnt_unit_pp2_reg[3] ;
  wire [3:0]col_en_host;
  wire [26:0]col_out;
  wire \col_sel_pp1[0]_i_2_n_0 ;
  wire \col_sel_pp1[0]_i_3_n_0 ;
  wire \col_sel_pp1[0]_i_4_n_0 ;
  wire \col_sel_pp1[0]_i_5_n_0 ;
  wire \col_sel_pp1_reg[1] ;
  wire [4:0]data_in;
  wire [31:0]enable_i;
  wire [31:0]\enable_i[31] ;
  wire enc_dec;
  wire enc_dec_sbox;
  wire first_block;
  wire first_block_reg;
  wire first_block_reg_0;
  wire first_block_reg_1;
  wire [1:0]g_func;
  wire [27:0]info_o;
  wire [4:0]\info_o[0]_0 ;
  wire \info_o[0]_INST_0_i_5_n_0 ;
  wire \info_o[10]_INST_0_i_4_n_0 ;
  wire \info_o[11]_INST_0_i_4_n_0 ;
  wire \info_o[12]_INST_0_i_4_n_0 ;
  wire \info_o[13]_INST_0_i_4_n_0 ;
  wire \info_o[14]_INST_0_i_4_n_0 ;
  wire \info_o[15]_INST_0_i_4_n_0 ;
  wire \info_o[16]_INST_0_i_5_n_0 ;
  wire \info_o[17]_INST_0_i_5_n_0 ;
  wire \info_o[18]_INST_0_i_5_n_0 ;
  wire \info_o[19]_INST_0_i_5_n_0 ;
  wire \info_o[20]_INST_0_i_5_n_0 ;
  wire \info_o[21]_INST_0_i_5_n_0 ;
  wire \info_o[22]_INST_0_i_5_n_0 ;
  wire \info_o[23]_INST_0_i_5_n_0 ;
  wire \info_o[24]_INST_0_i_6_n_0 ;
  wire \info_o[25]_INST_0_i_6_n_0 ;
  wire \info_o[26]_INST_0_i_6_n_0 ;
  wire \info_o[27]_INST_0_i_6_n_0 ;
  wire \info_o[28]_INST_0_i_15 ;
  wire \info_o[28]_INST_0_i_15_0 ;
  wire \info_o[28]_INST_0_i_8_n_0 ;
  wire \info_o[29]_INST_0_i_8_n_0 ;
  wire \info_o[30]_INST_0_i_8_n_0 ;
  wire \info_o[31] ;
  wire \info_o[31]_0 ;
  wire \info_o[31]_1 ;
  wire [31:0]\info_o[31]_2 ;
  wire [27:0]\info_o[31]_3 ;
  wire \info_o[31]_INST_0_i_12_0 ;
  wire \info_o[31]_INST_0_i_14_n_0 ;
  wire \info_o[31]_INST_0_i_16_n_0 ;
  wire \info_o[31]_INST_0_i_26_n_0 ;
  wire [0:0]\info_o[31]_INST_0_i_4 ;
  wire \info_o[31]_INST_0_i_4_0 ;
  wire [0:0]\info_o[31]_INST_0_i_4_1 ;
  wire \info_o[4]_INST_0_i_4_n_0 ;
  wire \info_o[6]_INST_0_i_4_n_0 ;
  wire \info_o[7]_INST_0_i_4_n_0 ;
  wire \info_o[8]_INST_0_i_4_n_0 ;
  wire \info_o[9]_INST_0_i_4_n_0 ;
  wire info_o_0_sn_1;
  wire info_o_10_sn_1;
  wire info_o_11_sn_1;
  wire info_o_12_sn_1;
  wire info_o_4_sn_1;
  wire info_o_6_sn_1;
  wire info_o_9_sn_1;
  wire isomorphism_inv_return033_out;
  wire isomorphism_inv_return033_out_12;
  wire isomorphism_inv_return033_out_6;
  wire isomorphism_inv_return03_out;
  wire isomorphism_inv_return03_out_13;
  wire isomorphism_inv_return03_out_7;
  wire isomorphism_inv_return05_out;
  wire isomorphism_inv_return05_out_14;
  wire isomorphism_inv_return05_out_8;
  wire isomorphism_return114_out;
  wire isomorphism_return114_out_1;
  wire isomorphism_return114_out_3;
  wire isomorphism_return114_out_5;
  wire isomorphism_return179_out;
  wire isomorphism_return179_out_0;
  wire isomorphism_return179_out_2;
  wire isomorphism_return179_out_4;
  wire iv_mux_out13_out;
  wire [31:0]iv_out;
  wire [3:0]key_en;
  wire [0:0]\key_en_pp1_reg[0] ;
  wire [0:0]\key_en_pp1_reg[1] ;
  wire [0:0]\key_en_pp1_reg[2] ;
  wire [0:0]\key_en_pp1_reg[3] ;
  wire \key_en_pp1_reg[3]_0 ;
  wire [127:0]key_in;
  wire [21:0]key_out;
  wire \key_out_sel_pp1_reg[1] ;
  wire key_sel;
  wire key_sel_mux;
  wire key_sel_pp1;
  wire last_round;
  wire \out_gf_pp[1]_i_2 ;
  wire \out_gf_pp[1]_i_2__0 ;
  wire \out_gf_pp[1]_i_2__1 ;
  wire \out_gf_pp[1]_i_2__2 ;
  wire p_16_in;
  wire p_16_in_11;
  wire p_16_in_17;
  wire p_86_in;
  wire p_86_in_15;
  wire p_86_in_9;
  wire p_93_in;
  wire p_93_in_10;
  wire p_93_in_16;
  wire \rd_count[0]_i_1_n_0 ;
  wire \rd_count[1]_i_1_n_0 ;
  wire \rd_count[1]_i_2_n_0 ;
  wire \rd_count[2]_i_1_n_0 ;
  wire \rd_count[2]_i_2_n_0 ;
  wire \rd_count[2]_i_3_n_0 ;
  wire \rd_count[3]_i_1_n_0 ;
  wire \rd_count[3]_i_2_n_0 ;
  wire \rd_count[3]_i_3_n_0 ;
  wire \rd_count[3]_i_4_n_0 ;
  wire \rd_count[3]_i_5_n_0 ;
  wire \rd_count[3]_i_6_n_0 ;
  wire \rd_count_reg[3]_0 ;
  wire [3:0]\rd_count_reg[3]_1 ;
  wire rk_out_sel_pp2;
  wire rst_i;
  wire [5:0]sbox_out_enc;
  wire [2:2]sbox_sel;

  assign info_o_0_sn_1 = info_o_0_sp_1;
  assign info_o_10_sn_1 = info_o_10_sp_1;
  assign info_o_11_sn_1 = info_o_11_sp_1;
  assign info_o_12_sn_1 = info_o_12_sp_1;
  assign info_o_4_sn_1 = info_o_4_sp_1;
  assign info_o_6_sn_1 = info_o_6_sp_1;
  assign info_o_9_sn_1 = info_o_9_sp_1;
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][0]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [0]),
        .I2(\CD[0].col[3][0]_i_2_n_0 ),
        .I3(add_rk_out[0]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [0]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][0]_i_10 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [0]),
        .O(\CD[0].col[3][0]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][0]_i_13 
       (.I0(\col_en_cnt_unit_pp2_reg[3] ),
        .I1(\info_o[31]_3 [0]),
        .O(\CD[0].col[3][0]_i_13_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][0]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[0]),
        .O(\CD[0].col[3][0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][0]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][0]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][0] ),
        .I4(\CD[2].col_reg[1][0]_0 ),
        .I5(\CD[0].col[3][0]_i_7_n_0 ),
        .O(\CD[0].col[3][0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][0]_i_4 
       (.I0(\CD[0].col[3][0]_i_10_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [0]),
        .I3(\CD[0].col[3][0]_i_2_0 ),
        .I4(\info_o[0]_INST_0_i_5_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][0]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [0]),
        .I2(\CD[0].col[3][0]_i_13_n_0 ),
        .I3(\info_o[0]_INST_0_i_5_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][0]_i_14_n_0 ),
        .O(\CD[0].col[3][0]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[0].col[3][10]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [10]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][10] ),
        .I4(\CD[0].col[3][10]_i_3_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [10]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \CD[0].col[3][10]_i_10 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [10]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [10]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [10]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][10] ));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \CD[0].col[3][10]_i_12 
       (.I0(\CD[0].col[3][31]_i_5_0 [10]),
        .I1(\CD[0].col[3][31]_i_10_0 [10]),
        .I2(\CD[0].col[3][10]_i_6_0 ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\CD[0].col[3][10]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \CD[0].col[3][10]_i_15 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[34]),
        .I5(key_in[2]),
        .O(\AES_CORE_DATAPATH/g_in [10]));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][10]_i_3 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][10]_i_6_n_0 ),
        .I3(\CD[1].col_reg[2][10]_0 ),
        .I4(\CD[1].col_reg[2][10]_1 ),
        .I5(\CD[0].col[3][10]_i_9_n_0 ),
        .O(\CD[0].col[3][10]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \CD[0].col[3][10]_i_6 
       (.I0(\CD[0].col[3][10]_i_12_n_0 ),
        .I1(\info_o[31]_INST_0_i_14_n_0 ),
        .I2(\info_o[31]_2 [10]),
        .I3(\CD[0].col[3][10]_i_3_0 ),
        .I4(\info_o[10]_INST_0_i_4_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][10]_i_9 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [10]),
        .I2(\CD[0].col[3][10]_i_3_0 ),
        .I3(\info_o[10]_INST_0_i_4_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp[3][10]_i_5_n_0 ),
        .O(\CD[0].col[3][10]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[0].col[3][11]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [11]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][11] ),
        .I4(\CD[0].col[3][11]_i_3_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [11]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \CD[0].col[3][11]_i_13 
       (.I0(\CD[0].col[3][31]_i_5_0 [11]),
        .I1(\CD[0].col[3][31]_i_10_0 [11]),
        .I2(\CD[0].col[3][10]_i_6_0 ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\CD[0].col[3][11]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][11]_i_3 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][11]_i_6_n_0 ),
        .I3(\CD[1].col_reg[2][11]_0 ),
        .I4(\CD[1].col_reg[2][11]_1 ),
        .I5(\CD[0].col[3][11]_i_9_n_0 ),
        .O(\CD[0].col[3][11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \CD[0].col[3][11]_i_6 
       (.I0(\CD[0].col[3][11]_i_13_n_0 ),
        .I1(\info_o[31]_INST_0_i_14_n_0 ),
        .I2(\info_o[31]_2 [11]),
        .I3(\CD[0].col[3][11]_i_3_0 ),
        .I4(\info_o[11]_INST_0_i_4_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][11]_i_9 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [11]),
        .I2(\CD[0].col[3][11]_i_3_0 ),
        .I3(\info_o[11]_INST_0_i_4_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp[3][11]_i_5_n_0 ),
        .O(\CD[0].col[3][11]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[0].col[3][12]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [12]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][12] ),
        .I4(\CD[0].col[3][12]_i_3_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [12]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \CD[0].col[3][12]_i_10 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [12]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [12]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [12]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][12] ));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \CD[0].col[3][12]_i_14 
       (.I0(\CD[0].col[3][31]_i_5_0 [12]),
        .I1(\CD[0].col[3][31]_i_10_0 [12]),
        .I2(\CD[0].col[3][10]_i_6_0 ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\CD[0].col[3][12]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \CD[0].col[3][12]_i_17 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[36]),
        .I5(key_in[4]),
        .O(\AES_CORE_DATAPATH/g_in [12]));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][12]_i_3 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][12]_i_6_n_0 ),
        .I3(\CD[1].col_reg[2][12]_0 ),
        .I4(\CD[1].col_reg[2][12]_1 ),
        .I5(\CD[0].col[3][12]_i_9_n_0 ),
        .O(\CD[0].col[3][12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \CD[0].col[3][12]_i_6 
       (.I0(\CD[0].col[3][12]_i_14_n_0 ),
        .I1(\info_o[31]_INST_0_i_14_n_0 ),
        .I2(\info_o[31]_2 [12]),
        .I3(\CD[0].col[3][12]_i_3_0 ),
        .I4(\info_o[12]_INST_0_i_4_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][12]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][12]_i_9 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [12]),
        .I2(\CD[0].col[3][12]_i_3_0 ),
        .I3(\info_o[12]_INST_0_i_4_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp[3][12]_i_5_n_0 ),
        .O(\CD[0].col[3][12]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[0].col[3][13]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [13]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][13] ),
        .I4(\CD[0].col[3][13]_i_3_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [13]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \CD[0].col[3][13]_i_11 
       (.I0(\CD[0].col[3][31]_i_5_0 [13]),
        .I1(\CD[0].col[3][31]_i_10_0 [13]),
        .I2(\CD[0].col[3][10]_i_6_0 ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\CD[0].col[3][13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][13]_i_3 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][13]_i_6_n_0 ),
        .I3(\CD[1].col_reg[2][13]_0 ),
        .I4(\CD[1].col_reg[2][13]_1 ),
        .I5(\CD[0].col[3][13]_i_9_n_0 ),
        .O(\CD[0].col[3][13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \CD[0].col[3][13]_i_6 
       (.I0(\CD[0].col[3][13]_i_11_n_0 ),
        .I1(\info_o[31]_INST_0_i_14_n_0 ),
        .I2(\info_o[31]_2 [13]),
        .I3(\CD[0].col[3][13]_i_3_0 ),
        .I4(\info_o[13]_INST_0_i_4_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][13]_i_9 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [13]),
        .I2(\CD[0].col[3][13]_i_3_0 ),
        .I3(\info_o[13]_INST_0_i_4_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp[3][13]_i_5_n_0 ),
        .O(\CD[0].col[3][13]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[0].col[3][14]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [14]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][14] ),
        .I4(\CD[0].col[3][14]_i_3_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [14]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][14]_i_11 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [14]),
        .O(\CD[0].col[3][14]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][14]_i_15 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[14]),
        .O(\CD[0].col[3][14]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][14]_i_3 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][14]_i_6_n_0 ),
        .I3(\CD[1].col_reg[2][14]_0 ),
        .I4(\CD[1].col_reg[2][14]_1 ),
        .I5(\IV_BKP_REGISTERS[2].iv_reg[2][14] ),
        .O(\CD[0].col[3][14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][14]_i_6 
       (.I0(\CD[0].col[3][14]_i_11_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [14]),
        .I3(\CD[0].col[3][14]_i_3_0 ),
        .I4(\info_o[14]_INST_0_i_4_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][14]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][14]_i_9 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [14]),
        .I2(\IV_BKP_REGISTERS[3].bkp[3][14]_i_2 ),
        .I3(\info_o[14]_INST_0_i_4_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][14]_i_15_n_0 ),
        .O(\IV_BKP_REGISTERS[2].iv_reg[2][14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[0].col[3][15]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [15]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][15] ),
        .I4(\CD[0].col[3][15]_i_5_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][15]_i_12 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [15]),
        .I2(\IV_BKP_REGISTERS[3].bkp[3][15]_i_4 ),
        .I3(\info_o[15]_INST_0_i_4_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][15]_i_20_n_0 ),
        .O(\IV_BKP_REGISTERS[2].iv_reg[2][15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \CD[0].col[3][15]_i_13 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [15]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [15]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [15]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][15] ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][15]_i_16 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [15]),
        .O(\CD[0].col[3][15]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \CD[0].col[3][15]_i_2 
       (.I0(\AES_CORE_DATAPATH/col_sel_w_bypass [0]),
        .I1(\AES_CORE_DATAPATH/col_sel_w_bypass [1]),
        .O(\FSM_sequential_state_reg[0]_2 ));
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][15]_i_20 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[15]),
        .O(\CD[0].col[3][15]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \CD[0].col[3][15]_i_21 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[39]),
        .I5(key_in[7]),
        .O(\AES_CORE_DATAPATH/g_in [15]));
  LUT6 #(
    .INIT(64'h00000000EEEEEE2E)) 
    \CD[0].col[3][15]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_0 [0]),
        .I1(\FSM_sequential_state_reg[2]_5 ),
        .I2(Q[0]),
        .I3(\col_sel_pp1[0]_i_3_n_0 ),
        .I4(\col_sel_pp1[0]_i_2_n_0 ),
        .I5(\AES_CORE_DATAPATH/col_sel_w_bypass [1]),
        .O(\CD[0].col[3][15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][15]_i_5 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][15]_i_9_n_0 ),
        .I3(\CD[1].col_reg[2][15]_0 ),
        .I4(\CD[1].col_reg[2][15]_1 ),
        .I5(\IV_BKP_REGISTERS[2].iv_reg[2][15] ),
        .O(\CD[0].col[3][15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEF000000EF)) 
    \CD[0].col[3][15]_i_6 
       (.I0(\col_sel_pp1[0]_i_2_n_0 ),
        .I1(\col_sel_pp1[0]_i_3_n_0 ),
        .I2(Q[0]),
        .I3(Q[2]),
        .I4(Q[3]),
        .I5(\CD[0].col[3][31]_i_7_0 [0]),
        .O(\AES_CORE_DATAPATH/col_sel_w_bypass [0]));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][15]_i_9 
       (.I0(\CD[0].col[3][15]_i_16_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [15]),
        .I3(\CD[0].col[3][15]_i_5_0 ),
        .I4(\info_o[15]_INST_0_i_4_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][15]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[0].col[3][16]_i_1 
       (.I0(\CD[0].col[3][16]_i_2_n_0 ),
        .I1(\CD[0].col[3][16]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [16]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [16]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [16]));
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][16]_i_12 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[16]),
        .O(\CD[0].col[3][16]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][16]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][16]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][16] ),
        .I4(\CD[1].col_reg[2][16]_0 ),
        .I5(\CD[0].col[3][16]_i_7_n_0 ),
        .O(\CD[0].col[3][16]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][16]_i_3 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[8]),
        .O(\CD[0].col[3][16]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][16]_i_4 
       (.I0(\CD[0].col[3][16]_i_8_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [16]),
        .I3(\CD[0].col[3][16]_i_2_1 ),
        .I4(\info_o[16]_INST_0_i_5_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][16]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][16]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [16]),
        .I2(\CD[0].col[3][16]_i_2_0 ),
        .I3(\info_o[16]_INST_0_i_5_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][16]_i_12_n_0 ),
        .O(\CD[0].col[3][16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][16]_i_8 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [16]),
        .O(\CD[0].col[3][16]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[0].col[3][17]_i_1 
       (.I0(\CD[0].col[3][17]_i_2_n_0 ),
        .I1(\CD[0].col[3][17]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [17]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [17]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [17]));
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][17]_i_12 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[17]),
        .O(\CD[0].col[3][17]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][17]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][17]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][17] ),
        .I4(\CD[1].col_reg[2][17]_0 ),
        .I5(\CD[0].col[3][17]_i_7_n_0 ),
        .O(\CD[0].col[3][17]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][17]_i_3 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[9]),
        .O(\CD[0].col[3][17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][17]_i_4 
       (.I0(\CD[0].col[3][17]_i_8_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [17]),
        .I3(\CD[0].col[3][17]_i_2_1 ),
        .I4(\info_o[17]_INST_0_i_5_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][17]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [17]),
        .I2(\CD[0].col[3][17]_i_2_0 ),
        .I3(\info_o[17]_INST_0_i_5_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][17]_i_12_n_0 ),
        .O(\CD[0].col[3][17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][17]_i_8 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [17]),
        .O(\CD[0].col[3][17]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[0].col[3][18]_i_1 
       (.I0(\CD[0].col[3][18]_i_2_n_0 ),
        .I1(\CD[0].col[3][18]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [18]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [18]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [18]));
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][18]_i_12 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[18]),
        .O(\CD[0].col[3][18]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][18]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][18]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][18] ),
        .I4(\CD[1].col_reg[2][18]_0 ),
        .I5(\CD[0].col[3][18]_i_7_n_0 ),
        .O(\CD[0].col[3][18]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][18]_i_3 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[10]),
        .O(\CD[0].col[3][18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][18]_i_4 
       (.I0(\CD[0].col[3][18]_i_8_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [18]),
        .I3(\CD[0].col[3][18]_i_2_1 ),
        .I4(\info_o[18]_INST_0_i_5_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][18]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][18]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [18]),
        .I2(\CD[0].col[3][18]_i_2_0 ),
        .I3(\info_o[18]_INST_0_i_5_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][18]_i_12_n_0 ),
        .O(\CD[0].col[3][18]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][18]_i_8 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [18]),
        .O(\CD[0].col[3][18]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[0].col[3][19]_i_1 
       (.I0(\CD[0].col[3][19]_i_2_n_0 ),
        .I1(\CD[0].col[3][19]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [19]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [19]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [19]));
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][19]_i_12 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[19]),
        .O(\CD[0].col[3][19]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][19]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][19]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][19] ),
        .I4(\CD[1].col_reg[2][19]_0 ),
        .I5(\CD[0].col[3][19]_i_7_n_0 ),
        .O(\CD[0].col[3][19]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][19]_i_3 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[11]),
        .O(\CD[0].col[3][19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][19]_i_4 
       (.I0(\CD[0].col[3][19]_i_8_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [19]),
        .I3(\CD[0].col[3][19]_i_2_1 ),
        .I4(\info_o[19]_INST_0_i_5_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][19]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][19]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [19]),
        .I2(\CD[0].col[3][19]_i_2_0 ),
        .I3(\info_o[19]_INST_0_i_5_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][19]_i_12_n_0 ),
        .O(\CD[0].col[3][19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][19]_i_8 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [19]),
        .O(\CD[0].col[3][19]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][1]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [1]),
        .I2(\CD[0].col[3][1]_i_2_n_0 ),
        .I3(add_rk_out[1]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [1]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][1]_i_10 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [1]),
        .O(\CD[0].col[3][1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \CD[0].col[3][1]_i_12 
       (.I0(\CD[0].col[3][31]_i_13_0 [1]),
        .I1(\CD[0].col[3][31]_i_13_1 [1]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\CD[0].col[3][1]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][1]_i_15 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[1]),
        .O(\CD[0].col[3][1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][1]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][1]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][1] ),
        .I4(\CD[2].col_reg[1][1]_0 ),
        .I5(\CD[0].col[3][1]_i_7_n_0 ),
        .O(\CD[0].col[3][1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][1]_i_4 
       (.I0(\CD[0].col[3][1]_i_10_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [1]),
        .I3(\CD[0].col[3][1]_i_2_1 ),
        .I4(\CD[0].col[3][1]_i_12_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][1]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [1]),
        .I2(\CD[0].col[3][1]_i_2_0 ),
        .I3(\CD[0].col[3][1]_i_12_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][1]_i_15_n_0 ),
        .O(\CD[0].col[3][1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[0].col[3][20]_i_1 
       (.I0(\CD[0].col[3][20]_i_2_n_0 ),
        .I1(\CD[0].col[3][20]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [20]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [20]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [20]));
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][20]_i_12 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[20]),
        .O(\CD[0].col[3][20]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][20]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][20]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][20] ),
        .I4(\CD[1].col_reg[2][20]_0 ),
        .I5(\CD[0].col[3][20]_i_7_n_0 ),
        .O(\CD[0].col[3][20]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][20]_i_3 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[12]),
        .O(\CD[0].col[3][20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][20]_i_4 
       (.I0(\CD[0].col[3][20]_i_8_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [20]),
        .I3(\CD[0].col[3][20]_i_2_1 ),
        .I4(\info_o[20]_INST_0_i_5_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][20]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][20]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [20]),
        .I2(\CD[0].col[3][20]_i_2_0 ),
        .I3(\info_o[20]_INST_0_i_5_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][20]_i_12_n_0 ),
        .O(\CD[0].col[3][20]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][20]_i_8 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [20]),
        .O(\CD[0].col[3][20]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[0].col[3][21]_i_1 
       (.I0(\CD[0].col[3][21]_i_2_n_0 ),
        .I1(\CD[0].col[3][21]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [21]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [21]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [21]));
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][21]_i_12 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[21]),
        .O(\CD[0].col[3][21]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][21]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][21]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][21] ),
        .I4(\CD[1].col_reg[2][21]_0 ),
        .I5(\CD[0].col[3][21]_i_7_n_0 ),
        .O(\CD[0].col[3][21]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][21]_i_3 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[13]),
        .O(\CD[0].col[3][21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][21]_i_4 
       (.I0(\CD[0].col[3][21]_i_8_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [21]),
        .I3(\CD[0].col[3][21]_i_2_1 ),
        .I4(\info_o[21]_INST_0_i_5_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][21]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [21]),
        .I2(\CD[0].col[3][21]_i_2_0 ),
        .I3(\info_o[21]_INST_0_i_5_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][21]_i_12_n_0 ),
        .O(\CD[0].col[3][21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][21]_i_8 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [21]),
        .O(\CD[0].col[3][21]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[0].col[3][22]_i_1 
       (.I0(\CD[0].col[3][22]_i_2_n_0 ),
        .I1(\CD[0].col[3][22]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [22]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [22]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [22]));
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][22]_i_12 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[22]),
        .O(\CD[0].col[3][22]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][22]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][22]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][22] ),
        .I4(\CD[1].col_reg[2][22]_0 ),
        .I5(\CD[0].col[3][22]_i_7_n_0 ),
        .O(\CD[0].col[3][22]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][22]_i_3 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[14]),
        .O(\CD[0].col[3][22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][22]_i_4 
       (.I0(\CD[0].col[3][22]_i_8_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [22]),
        .I3(\CD[0].col[3][22]_i_2_1 ),
        .I4(\info_o[22]_INST_0_i_5_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][22]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][22]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [22]),
        .I2(\CD[0].col[3][22]_i_2_0 ),
        .I3(\info_o[22]_INST_0_i_5_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][22]_i_12_n_0 ),
        .O(\CD[0].col[3][22]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][22]_i_8 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [22]),
        .O(\CD[0].col[3][22]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[0].col[3][23]_i_1 
       (.I0(\CD[0].col[3][23]_i_2_n_0 ),
        .I1(\CD[0].col[3][23]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [23]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [23]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [23]));
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][23]_i_13 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[23]),
        .O(\CD[0].col[3][23]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][23]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][23]_i_5_n_0 ),
        .I3(\CD[1].col_reg[2][23]_0 ),
        .I4(\CD[1].col_reg[2][23]_1 ),
        .I5(\CD[0].col[3][23]_i_8_n_0 ),
        .O(\CD[0].col[3][23]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][23]_i_3 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[15]),
        .O(\CD[0].col[3][23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA08AA08AA08AA)) 
    \CD[0].col[3][23]_i_4 
       (.I0(\FSM_sequential_state_reg[0]_2 ),
        .I1(\info_o[0]_0 [3]),
        .I2(\info_o[0]_0 [2]),
        .I3(\info_o[0]_0 [1]),
        .I4(Q[1]),
        .I5(Q[2]),
        .O(\CD[0].col[3][23]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][23]_i_5 
       (.I0(\CD[0].col[3][23]_i_9_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [23]),
        .I3(\CD[0].col[3][23]_i_2_1 ),
        .I4(\info_o[23]_INST_0_i_5_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][23]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][23]_i_8 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [23]),
        .I2(\CD[0].col[3][23]_i_2_0 ),
        .I3(\info_o[23]_INST_0_i_5_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][23]_i_13_n_0 ),
        .O(\CD[0].col[3][23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][23]_i_9 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [23]),
        .O(\CD[0].col[3][23]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][24]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [24]),
        .I2(\CD[0].col[3][24]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][24] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [24]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][24]_i_10 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [24]),
        .O(\CD[0].col[3][24]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][24]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[24]),
        .O(\CD[0].col[3][24]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][24]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][24]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][24]_0 ),
        .I4(\CD[2].col_reg[1][24]_1 ),
        .I5(\IV_BKP_REGISTERS[2].iv_reg[2][24] ),
        .O(\CD[0].col[3][24]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][24]_i_4 
       (.I0(\CD[0].col[3][24]_i_10_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [24]),
        .I3(\CD[0].col[3][24]_i_2_0 ),
        .I4(\info_o[24]_INST_0_i_6_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][24]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][24]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [24]),
        .I2(\IV_BKP_REGISTERS[2].bkp[2][24]_i_2 ),
        .I3(\info_o[24]_INST_0_i_6_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][24]_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[2].iv_reg[2][24] ));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][25]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [25]),
        .I2(\CD[0].col[3][25]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][25] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [25]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][25]_i_10 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [25]),
        .O(\CD[0].col[3][25]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][25]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[25]),
        .O(\CD[0].col[3][25]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][25]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][25]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][25]_0 ),
        .I4(\CD[2].col_reg[1][25]_1 ),
        .I5(\IV_BKP_REGISTERS[2].iv_reg[2][25] ),
        .O(\CD[0].col[3][25]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][25]_i_4 
       (.I0(\CD[0].col[3][25]_i_10_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [25]),
        .I3(\CD[0].col[3][25]_i_2_0 ),
        .I4(\info_o[25]_INST_0_i_6_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][25]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][25]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [25]),
        .I2(\IV_BKP_REGISTERS[2].bkp[2][25]_i_2 ),
        .I3(\info_o[25]_INST_0_i_6_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][25]_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[2].iv_reg[2][25] ));
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][26]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [26]),
        .I2(\CD[0].col[3][26]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][26] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [26]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][26]_i_10 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [26]),
        .O(\CD[0].col[3][26]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][26]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[26]),
        .O(\CD[0].col[3][26]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \CD[0].col[3][26]_i_15 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [26]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [26]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [26]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][26] ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][26]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][26]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][26]_0 ),
        .I4(\CD[2].col_reg[1][26]_1 ),
        .I5(\IV_BKP_REGISTERS[2].iv_reg[2][26] ),
        .O(\CD[0].col[3][26]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \CD[0].col[3][26]_i_20 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[50]),
        .I5(key_in[18]),
        .O(\AES_CORE_DATAPATH/g_in [26]));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][26]_i_4 
       (.I0(\CD[0].col[3][26]_i_10_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [26]),
        .I3(\CD[0].col[3][26]_i_2_0 ),
        .I4(\info_o[26]_INST_0_i_6_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][26]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][26]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [26]),
        .I2(\IV_BKP_REGISTERS[2].bkp[2][26]_i_2 ),
        .I3(\info_o[26]_INST_0_i_6_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][26]_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[2].iv_reg[2][26] ));
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][27]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [27]),
        .I2(\CD[0].col[3][27]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][27] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [27]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][27]_i_10 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [27]),
        .O(\CD[0].col[3][27]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][27]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[27]),
        .O(\CD[0].col[3][27]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][27]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][27]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][27]_0 ),
        .I4(\CD[2].col_reg[1][27]_1 ),
        .I5(\IV_BKP_REGISTERS[2].iv_reg[2][27] ),
        .O(\CD[0].col[3][27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][27]_i_4 
       (.I0(\CD[0].col[3][27]_i_10_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [27]),
        .I3(\CD[0].col[3][27]_i_2_0 ),
        .I4(\info_o[27]_INST_0_i_6_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][27]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][27]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [27]),
        .I2(\IV_BKP_REGISTERS[2].bkp[2][27]_i_2 ),
        .I3(\info_o[27]_INST_0_i_6_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][27]_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[2].iv_reg[2][27] ));
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][28]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [28]),
        .I2(\CD[0].col[3][28]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][28] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [28]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \CD[0].col[3][28]_i_10 
       (.I0(\CD[0].col[3][31]_i_5_0 [28]),
        .I1(\CD[0].col[3][31]_i_10_0 [28]),
        .I2(\CD[0].col[3][10]_i_6_0 ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\CD[0].col[3][28]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \CD[0].col[3][28]_i_13 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [28]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [28]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [28]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][28] ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][28]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][28]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][28]_0 ),
        .I4(\CD[2].col_reg[1][28]_1 ),
        .I5(\CD[0].col[3][28]_i_7_n_0 ),
        .O(\CD[0].col[3][28]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \CD[0].col[3][28]_i_20 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[52]),
        .I5(key_in[20]),
        .O(\AES_CORE_DATAPATH/g_in [28]));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \CD[0].col[3][28]_i_4 
       (.I0(\CD[0].col[3][28]_i_10_n_0 ),
        .I1(\info_o[31]_INST_0_i_14_n_0 ),
        .I2(\info_o[31]_2 [28]),
        .I3(\CD[0].col[3][28]_i_2_0 ),
        .I4(\info_o[28]_INST_0_i_8_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][28]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][28]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [28]),
        .I2(\CD[0].col[3][28]_i_2_0 ),
        .I3(\info_o[28]_INST_0_i_8_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\IV_BKP_REGISTERS[2].bkp[2][28]_i_5_n_0 ),
        .O(\CD[0].col[3][28]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][29]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [29]),
        .I2(\CD[0].col[3][29]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][29] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [29]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][29]_i_10 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [29]),
        .O(\CD[0].col[3][29]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][29]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[29]),
        .O(\CD[0].col[3][29]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][29]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][29]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][29]_0 ),
        .I4(\CD[2].col_reg[1][29]_1 ),
        .I5(\IV_BKP_REGISTERS[2].iv_reg[2][29] ),
        .O(\CD[0].col[3][29]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][29]_i_4 
       (.I0(\CD[0].col[3][29]_i_10_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [29]),
        .I3(\CD[0].col[3][29]_i_2_0 ),
        .I4(\info_o[29]_INST_0_i_8_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][29]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][29]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [29]),
        .I2(\IV_BKP_REGISTERS[2].bkp[2][29]_i_2 ),
        .I3(\info_o[29]_INST_0_i_8_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][29]_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[2].iv_reg[2][29] ));
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][2]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [2]),
        .I2(\CD[0].col[3][2]_i_2_n_0 ),
        .I3(add_rk_out[2]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [2]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][2]_i_10 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [2]),
        .O(\CD[0].col[3][2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \CD[0].col[3][2]_i_12 
       (.I0(\CD[0].col[3][31]_i_13_0 [2]),
        .I1(\CD[0].col[3][31]_i_13_1 [2]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\CD[0].col[3][2]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][2]_i_15 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[2]),
        .O(\CD[0].col[3][2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \CD[0].col[3][2]_i_16 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [2]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [2]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [2]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][2] ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][2]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][2]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][2] ),
        .I4(\CD[2].col_reg[1][2]_0 ),
        .I5(\CD[0].col[3][2]_i_7_n_0 ),
        .O(\CD[0].col[3][2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \CD[0].col[3][2]_i_20 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[58]),
        .I5(key_in[26]),
        .O(\AES_CORE_DATAPATH/g_in [2]));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][2]_i_4 
       (.I0(\CD[0].col[3][2]_i_10_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [2]),
        .I3(\CD[0].col[3][2]_i_2_1 ),
        .I4(\CD[0].col[3][2]_i_12_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][2]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [2]),
        .I2(\CD[0].col[3][2]_i_2_0 ),
        .I3(\CD[0].col[3][2]_i_12_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][2]_i_15_n_0 ),
        .O(\CD[0].col[3][2]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][30]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [30]),
        .I2(\CD[0].col[3][30]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][30] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [30]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][30]_i_10 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [30]),
        .O(\CD[0].col[3][30]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][30]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[30]),
        .O(\CD[0].col[3][30]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][30]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][30]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][30]_0 ),
        .I4(\CD[2].col_reg[1][30]_1 ),
        .I5(\IV_BKP_REGISTERS[2].iv_reg[2][30] ),
        .O(\CD[0].col[3][30]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][30]_i_4 
       (.I0(\CD[0].col[3][30]_i_10_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [30]),
        .I3(\CD[0].col[3][30]_i_2_0 ),
        .I4(\info_o[30]_INST_0_i_8_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][30]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][30]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [30]),
        .I2(\IV_BKP_REGISTERS[2].bkp[2][30]_i_2 ),
        .I3(\info_o[30]_INST_0_i_8_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][30]_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[2].iv_reg[2][30] ));
  LUT6 #(
    .INIT(64'hFFE2E2E2E2E2E2E2)) 
    \CD[0].col[3][31]_i_1 
       (.I0(\CD[0].col_reg[3][31]_1 [3]),
        .I1(\FSM_sequential_state_reg[2]_5 ),
        .I2(\FSM_sequential_state_reg[2]_2 [3]),
        .I3(\CD[3].col_reg[0][31]_2 [0]),
        .I4(\CD[3].col_reg[0][31]_2 [1]),
        .I5(\CD[3].col_reg[0][31]_3 ),
        .O(E));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][31]_i_10 
       (.I0(\CD[0].col[3][31]_i_18_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [31]),
        .I3(\CD[0].col[3][31]_i_5_1 ),
        .I4(\info_o[31]_INST_0_i_16_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][31]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][31]_i_13 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [31]),
        .I2(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2 ),
        .I3(\info_o[31]_INST_0_i_16_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][31]_i_28_n_0 ),
        .O(\IV_BKP_REGISTERS[2].iv_reg[2][31] ));
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \CD[0].col[3][31]_i_15 
       (.I0(rk_out_sel_pp2),
        .I1(Q[3]),
        .I2(Q[2]),
        .O(add_rk_sel));
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \CD[0].col[3][31]_i_17 
       (.I0(D[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(\CD[0].col[3][31]_i_7_0 [1]),
        .O(\AES_CORE_DATAPATH/col_sel_w_bypass [1]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][31]_i_18 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [31]),
        .O(\CD[0].col[3][31]_i_18_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT5 #(
    .INIT(32'h00150000)) 
    \CD[0].col[3][31]_i_19 
       (.I0(\col_en_cnt_unit_pp2_reg[3] ),
        .I1(\key_en_pp1_reg[3]_0 ),
        .I2(first_block),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .O(first_block_reg));
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][31]_i_2 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [31]),
        .I2(\CD[0].col[3][31]_i_5_n_0 ),
        .I3(\CD[2].col_reg[1][31]_2 ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [31]));
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT4 #(
    .INIT(16'h002A)) 
    \CD[0].col[3][31]_i_23 
       (.I0(iv_mux_out13_out),
        .I1(first_block),
        .I2(\key_en_pp1_reg[3]_0 ),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .O(first_block_reg_1));
  LUT5 #(
    .INIT(32'h0000DF00)) 
    \CD[0].col[3][31]_i_27 
       (.I0(\rd_count_reg[3]_1 [3]),
        .I1(\rd_count_reg[3]_1 [2]),
        .I2(\rd_count_reg[3]_1 [1]),
        .I3(\info_o[0]_0 [3]),
        .I4(\info_o[0]_0 [2]),
        .O(\CD[0].col[3][31]_i_27_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][31]_i_28 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[31]),
        .O(\CD[0].col[3][31]_i_28_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \CD[0].col[3][31]_i_3 
       (.I0(Q[2]),
        .I1(Q[3]),
        .O(\FSM_sequential_state_reg[2]_5 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \CD[0].col[3][31]_i_30 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [31]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [31]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [31]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][31]_1 ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \CD[0].col[3][31]_i_38 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[55]),
        .I5(key_in[23]),
        .O(\AES_CORE_DATAPATH/g_in [31]));
  LUT6 #(
    .INIT(64'h0000A200A200A200)) 
    \CD[0].col[3][31]_i_4 
       (.I0(\FSM_sequential_state_reg[0]_2 ),
        .I1(\info_o[0]_0 [3]),
        .I2(\info_o[0]_0 [2]),
        .I3(\info_o[0]_0 [1]),
        .I4(Q[1]),
        .I5(Q[2]),
        .O(\CD[0].col[3][31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][31]_i_5 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][31]_i_10_n_0 ),
        .I3(\CD[2].col_reg[1][31]_3 ),
        .I4(\CD[2].col_reg[1][31]_4 ),
        .I5(\IV_BKP_REGISTERS[2].iv_reg[2][31] ),
        .O(\CD[0].col[3][31]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF40555555)) 
    \CD[0].col[3][31]_i_7 
       (.I0(\AES_CORE_DATAPATH/col_sel_w_bypass [1]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(\info_o[0]_0 [1]),
        .I4(\key_en_pp1_reg[3]_0 ),
        .I5(\CD[0].col[3][15]_i_3_n_0 ),
        .O(\CD[0].col[3][31]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \CD[0].col[3][31]_i_8 
       (.I0(\AES_CORE_DATAPATH/col_sel_w_bypass [1]),
        .I1(\AES_CORE_DATAPATH/col_sel_w_bypass [0]),
        .O(\CD[0].col[3][31]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][3]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [3]),
        .I2(\CD[0].col[3][3]_i_2_n_0 ),
        .I3(add_rk_out[3]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [3]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][3]_i_10 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [3]),
        .O(\CD[0].col[3][3]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \CD[0].col[3][3]_i_12 
       (.I0(\CD[0].col[3][31]_i_13_0 [3]),
        .I1(\CD[0].col[3][31]_i_13_1 [3]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\CD[0].col[3][3]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][3]_i_15 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[3]),
        .O(\CD[0].col[3][3]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][3]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][3]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][3] ),
        .I4(\CD[2].col_reg[1][3]_0 ),
        .I5(\CD[0].col[3][3]_i_7_n_0 ),
        .O(\CD[0].col[3][3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][3]_i_4 
       (.I0(\CD[0].col[3][3]_i_10_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [3]),
        .I3(\CD[0].col[3][3]_i_2_1 ),
        .I4(\CD[0].col[3][3]_i_12_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][3]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [3]),
        .I2(\CD[0].col[3][3]_i_2_0 ),
        .I3(\CD[0].col[3][3]_i_12_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][3]_i_15_n_0 ),
        .O(\CD[0].col[3][3]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][4]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [4]),
        .I2(\CD[0].col[3][4]_i_2_n_0 ),
        .I3(add_rk_out[4]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [4]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][4]_i_10 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [4]),
        .O(\CD[0].col[3][4]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][4]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[4]),
        .O(\CD[0].col[3][4]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \CD[0].col[3][4]_i_15 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [4]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [4]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [4]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][4] ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \CD[0].col[3][4]_i_18 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[60]),
        .I5(key_in[28]),
        .O(\AES_CORE_DATAPATH/g_in [4]));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][4]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][4]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][4] ),
        .I4(\CD[2].col_reg[1][4]_0 ),
        .I5(\CD[0].col[3][4]_i_7_n_0 ),
        .O(\CD[0].col[3][4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][4]_i_4 
       (.I0(\CD[0].col[3][4]_i_10_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [4]),
        .I3(\CD[0].col[3][4]_i_2_1 ),
        .I4(\info_o[4]_INST_0_i_4_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][4]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [4]),
        .I2(\CD[0].col[3][4]_i_2_0 ),
        .I3(\info_o[4]_INST_0_i_4_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][4]_i_14_n_0 ),
        .O(\CD[0].col[3][4]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][5]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [5]),
        .I2(\CD[0].col[3][5]_i_2_n_0 ),
        .I3(add_rk_out[5]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [5]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][5]_i_10 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [5]),
        .O(\CD[0].col[3][5]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \CD[0].col[3][5]_i_12 
       (.I0(\CD[0].col[3][31]_i_13_0 [5]),
        .I1(\CD[0].col[3][31]_i_13_1 [5]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\CD[0].col[3][5]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][5]_i_15 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[5]),
        .O(\CD[0].col[3][5]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][5]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][5]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][5] ),
        .I4(\CD[2].col_reg[1][5]_0 ),
        .I5(\CD[0].col[3][5]_i_7_n_0 ),
        .O(\CD[0].col[3][5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][5]_i_4 
       (.I0(\CD[0].col[3][5]_i_10_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [5]),
        .I3(\CD[0].col[3][5]_i_2_1 ),
        .I4(\CD[0].col[3][5]_i_12_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][5]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [5]),
        .I2(\CD[0].col[3][5]_i_2_0 ),
        .I3(\CD[0].col[3][5]_i_12_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][5]_i_15_n_0 ),
        .O(\CD[0].col[3][5]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][6]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [6]),
        .I2(\CD[0].col[3][6]_i_2_n_0 ),
        .I3(add_rk_out[6]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [6]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][6]_i_10 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [6]),
        .O(\CD[0].col[3][6]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][6]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[6]),
        .O(\CD[0].col[3][6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][6]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][6]_i_4_n_0 ),
        .I3(\CD[2].col_reg[1][6] ),
        .I4(\CD[2].col_reg[1][6]_0 ),
        .I5(\CD[0].col[3][6]_i_7_n_0 ),
        .O(\CD[0].col[3][6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][6]_i_4 
       (.I0(\CD[0].col[3][6]_i_10_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [6]),
        .I3(\CD[0].col[3][6]_i_2_1 ),
        .I4(\info_o[6]_INST_0_i_4_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][6]_i_7 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [6]),
        .I2(\CD[0].col[3][6]_i_2_0 ),
        .I3(\info_o[6]_INST_0_i_4_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][6]_i_14_n_0 ),
        .O(\CD[0].col[3][6]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[0].col[3][7]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [7]),
        .I2(\CD[0].col[3][7]_i_2_n_0 ),
        .I3(add_rk_out[7]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [7]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][7]_i_11 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [7]),
        .O(\CD[0].col[3][7]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][7]_i_15 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[7]),
        .O(\CD[0].col[3][7]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \CD[0].col[3][7]_i_16 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [7]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [7]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [7]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][7] ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][7]_i_2 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][7]_i_5_n_0 ),
        .I3(\CD[2].col_reg[1][7] ),
        .I4(\CD[2].col_reg[1][7]_0 ),
        .I5(\CD[0].col[3][7]_i_8_n_0 ),
        .O(\CD[0].col[3][7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \CD[0].col[3][7]_i_20 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[63]),
        .I5(key_in[31]),
        .O(\AES_CORE_DATAPATH/g_in [7]));
  LUT6 #(
    .INIT(64'hFFFFFFFF00007000)) 
    \CD[0].col[3][7]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\AES_CORE_DATAPATH/col_sel_w_bypass [1]),
        .I5(\CD[0].col[3][15]_i_3_n_0 ),
        .O(\CD[0].col[3][7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][7]_i_5 
       (.I0(\CD[0].col[3][7]_i_11_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [7]),
        .I3(\CD[0].col[3][7]_i_2_1 ),
        .I4(\info_o[7]_INST_0_i_4_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][7]_i_8 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [7]),
        .I2(\CD[0].col[3][7]_i_2_0 ),
        .I3(\info_o[7]_INST_0_i_4_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][7]_i_15_n_0 ),
        .O(\CD[0].col[3][7]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[0].col[3][8]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [8]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][8] ),
        .I4(\CD[0].col[3][8]_i_3_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [8]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][8]_i_12 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [8]),
        .O(\CD[0].col[3][8]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][8]_i_16 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[8]),
        .O(\CD[0].col[3][8]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][8]_i_3 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][8]_i_6_n_0 ),
        .I3(\CD[1].col_reg[2][8]_0 ),
        .I4(\CD[1].col_reg[2][8]_1 ),
        .I5(\IV_BKP_REGISTERS[2].iv_reg[2][8] ),
        .O(\CD[0].col[3][8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][8]_i_6 
       (.I0(\CD[0].col[3][8]_i_12_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [8]),
        .I3(\CD[0].col[3][8]_i_3_0 ),
        .I4(\info_o[8]_INST_0_i_4_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][8]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][8]_i_9 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [8]),
        .I2(\IV_BKP_REGISTERS[3].bkp[3][8]_i_2 ),
        .I3(\info_o[8]_INST_0_i_4_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][8]_i_16_n_0 ),
        .O(\IV_BKP_REGISTERS[2].iv_reg[2][8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[0].col[3][9]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [9]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][9] ),
        .I4(\CD[0].col[3][9]_i_3_n_0 ),
        .O(\CD[0].col_reg[3][31]_0 [9]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \CD[0].col[3][9]_i_11 
       (.I0(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .I1(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][0]_i_4_0 ),
        .I4(\col_en_cnt_unit_pp2_reg[3] ),
        .I5(\CD[0].col[3][31]_i_10_0 [9]),
        .O(\CD[0].col[3][9]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][9]_i_15 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[9]),
        .O(\CD[0].col[3][9]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88800008)) 
    \CD[0].col[3][9]_i_3 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\CD[2].col_reg[1][31]_1 ),
        .I2(\CD[0].col[3][9]_i_6_n_0 ),
        .I3(\CD[1].col_reg[2][9]_0 ),
        .I4(\CD[1].col_reg[2][9]_1 ),
        .I5(\IV_BKP_REGISTERS[2].iv_reg[2][9] ),
        .O(\CD[0].col[3][9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAEAEAEAEA)) 
    \CD[0].col[3][9]_i_6 
       (.I0(\CD[0].col[3][9]_i_11_n_0 ),
        .I1(first_block_reg),
        .I2(\CD[0].col[3][31]_i_5_0 [9]),
        .I3(\CD[0].col[3][9]_i_3_0 ),
        .I4(\info_o[9]_INST_0_i_4_n_0 ),
        .I5(\CD[0].col[3][5]_i_2_2 ),
        .O(\CD[0].col[3][9]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF80000)) 
    \CD[0].col[3][9]_i_9 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [9]),
        .I2(\IV_BKP_REGISTERS[3].bkp[3][9]_i_2 ),
        .I3(\info_o[9]_INST_0_i_4_n_0 ),
        .I4(\CD[0].col[3][31]_i_27_n_0 ),
        .I5(\CD[0].col[3][9]_i_15_n_0 ),
        .O(\IV_BKP_REGISTERS[2].iv_reg[2][9] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[1].col[2][0]_i_1 
       (.I0(\CD[0].col[3][0]_i_2_n_0 ),
        .I1(\CD[1].col[2][0]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [0]),
        .I4(\CD[2].col_reg[1][31]_0 [0]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [0]));
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[1].col[2][0]_i_2 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[0]),
        .O(\CD[1].col[2][0]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][10]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [10]),
        .I2(\CD[0].col[3][10]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][10] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [10]));
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][11]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [11]),
        .I2(\CD[0].col[3][11]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][11] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [11]));
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][12]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [12]),
        .I2(\CD[0].col[3][12]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][12] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [12]));
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][13]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [13]),
        .I2(\CD[0].col[3][13]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][13] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [13]));
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][14]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [14]),
        .I2(\CD[0].col[3][14]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][14] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [14]));
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][15]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [15]),
        .I2(\CD[0].col[3][15]_i_5_n_0 ),
        .I3(\CD[1].col_reg[2][15] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [15]));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][16]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [16]),
        .I2(\CD[0].col[3][16]_i_2_n_0 ),
        .I3(add_rk_out[8]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[1].col_reg[2][31] [16]));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][17]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [17]),
        .I2(\CD[0].col[3][17]_i_2_n_0 ),
        .I3(add_rk_out[9]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[1].col_reg[2][31] [17]));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][18]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [18]),
        .I2(\CD[0].col[3][18]_i_2_n_0 ),
        .I3(add_rk_out[10]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[1].col_reg[2][31] [18]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \CD[1].col[2][18]_i_5 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [18]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [18]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [18]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][18] ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \CD[1].col[2][18]_i_7 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[42]),
        .I5(key_in[10]),
        .O(\AES_CORE_DATAPATH/g_in [18]));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][19]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [19]),
        .I2(\CD[0].col[3][19]_i_2_n_0 ),
        .I3(add_rk_out[11]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[1].col_reg[2][31] [19]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[1].col[2][1]_i_1 
       (.I0(\CD[0].col[3][1]_i_2_n_0 ),
        .I1(\CD[1].col[2][1]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [1]),
        .I4(\CD[2].col_reg[1][31]_0 [1]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [1]));
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[1].col[2][1]_i_2 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[1]),
        .O(\CD[1].col[2][1]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][20]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [20]),
        .I2(\CD[0].col[3][20]_i_2_n_0 ),
        .I3(add_rk_out[12]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[1].col_reg[2][31] [20]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \CD[1].col[2][20]_i_5 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [20]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [20]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [20]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][20] ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \CD[1].col[2][20]_i_9 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[44]),
        .I5(key_in[12]),
        .O(\AES_CORE_DATAPATH/g_in [20]));
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][21]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [21]),
        .I2(\CD[0].col[3][21]_i_2_n_0 ),
        .I3(add_rk_out[13]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[1].col_reg[2][31] [21]));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][22]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [22]),
        .I2(\CD[0].col[3][22]_i_2_n_0 ),
        .I3(add_rk_out[14]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[1].col_reg[2][31] [22]));
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][23]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [23]),
        .I2(\CD[0].col[3][23]_i_2_n_0 ),
        .I3(add_rk_out[15]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[1].col_reg[2][31] [23]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \CD[1].col[2][23]_i_5 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [23]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [23]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [23]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][23] ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \CD[1].col[2][23]_i_7 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[47]),
        .I5(key_in[15]),
        .O(\AES_CORE_DATAPATH/g_in [23]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[1].col[2][24]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [24]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][24] ),
        .I4(\CD[0].col[3][24]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [24]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[1].col[2][25]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [25]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][25] ),
        .I4(\CD[0].col[3][25]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [25]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[1].col[2][26]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [26]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][26] ),
        .I4(\CD[0].col[3][26]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [26]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[1].col[2][27]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [27]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][27] ),
        .I4(\CD[0].col[3][27]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [27]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[1].col[2][28]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [28]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][28] ),
        .I4(\CD[0].col[3][28]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [28]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[1].col[2][29]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [29]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][29] ),
        .I4(\CD[0].col[3][29]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [29]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[1].col[2][2]_i_1 
       (.I0(\CD[0].col[3][2]_i_2_n_0 ),
        .I1(\CD[1].col[2][2]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [2]),
        .I4(\CD[2].col_reg[1][31]_0 [2]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [2]));
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[1].col[2][2]_i_2 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[2]),
        .O(\CD[1].col[2][2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[1].col[2][30]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [30]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][30] ),
        .I4(\CD[0].col[3][30]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [30]));
  LUT6 #(
    .INIT(64'hE2E2E2E2FFE2E2E2)) 
    \CD[1].col[2][31]_i_1 
       (.I0(\CD[0].col_reg[3][31]_1 [2]),
        .I1(\FSM_sequential_state_reg[2]_5 ),
        .I2(\FSM_sequential_state_reg[2]_2 [2]),
        .I3(\CD[3].col_reg[0][31]_3 ),
        .I4(\CD[3].col_reg[0][31]_2 [1]),
        .I5(\CD[3].col_reg[0][31]_2 [0]),
        .O(\col_en_cnt_unit_pp2_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[1].col[2][31]_i_2 
       (.I0(\CD[1].col_reg[2][31]_0 [31]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][31]_2 ),
        .I4(\CD[0].col[3][31]_i_5_n_0 ),
        .O(\CD[1].col_reg[2][31] [31]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[1].col[2][3]_i_1 
       (.I0(\CD[0].col[3][3]_i_2_n_0 ),
        .I1(\CD[1].col[2][3]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [3]),
        .I4(\CD[2].col_reg[1][31]_0 [3]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [3]));
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[1].col[2][3]_i_2 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[3]),
        .O(\CD[1].col[2][3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[1].col[2][4]_i_1 
       (.I0(\CD[0].col[3][4]_i_2_n_0 ),
        .I1(\CD[1].col[2][4]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [4]),
        .I4(\CD[2].col_reg[1][31]_0 [4]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [4]));
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[1].col[2][4]_i_2 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[4]),
        .O(\CD[1].col[2][4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[1].col[2][5]_i_1 
       (.I0(\CD[0].col[3][5]_i_2_n_0 ),
        .I1(\CD[1].col[2][5]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [5]),
        .I4(\CD[2].col_reg[1][31]_0 [5]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [5]));
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[1].col[2][5]_i_2 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[5]),
        .O(\CD[1].col[2][5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[1].col[2][6]_i_1 
       (.I0(\CD[0].col[3][6]_i_2_n_0 ),
        .I1(\CD[1].col[2][6]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [6]),
        .I4(\CD[2].col_reg[1][31]_0 [6]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [6]));
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[1].col[2][6]_i_2 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[6]),
        .O(\CD[1].col[2][6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[1].col[2][7]_i_1 
       (.I0(\CD[0].col[3][7]_i_2_n_0 ),
        .I1(\CD[1].col[2][7]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [7]),
        .I4(\CD[2].col_reg[1][31]_0 [7]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [7]));
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[1].col[2][7]_i_2 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(add_rk_out[7]),
        .O(\CD[1].col[2][7]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][8]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [8]),
        .I2(\CD[0].col[3][8]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][8] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [8]));
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[1].col[2][9]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [9]),
        .I2(\CD[0].col[3][9]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][9] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[1].col_reg[2][31] [9]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[2].col[1][0]_i_1 
       (.I0(\CD[0].col[3][0]_i_2_n_0 ),
        .I1(\CD[1].col[2][0]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [0]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [0]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [0]));
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][10]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [10]),
        .I2(\CD[0].col[3][10]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][10] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[2].col_reg[1][31] [10]));
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][11]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [11]),
        .I2(\CD[0].col[3][11]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][11] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[2].col_reg[1][31] [11]));
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][12]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [12]),
        .I2(\CD[0].col[3][12]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][12] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[2].col_reg[1][31] [12]));
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][13]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [13]),
        .I2(\CD[0].col[3][13]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][13] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[2].col_reg[1][31] [13]));
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][14]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [14]),
        .I2(\CD[0].col[3][14]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][14] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[2].col_reg[1][31] [14]));
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][15]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [15]),
        .I2(\CD[0].col[3][15]_i_5_n_0 ),
        .I3(\CD[1].col_reg[2][15] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[2].col_reg[1][31] [15]));
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][16]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [16]),
        .I2(\CD[0].col[3][16]_i_2_n_0 ),
        .I3(add_rk_out[8]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [16]));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][17]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [17]),
        .I2(\CD[0].col[3][17]_i_2_n_0 ),
        .I3(add_rk_out[9]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [17]));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][18]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [18]),
        .I2(\CD[0].col[3][18]_i_2_n_0 ),
        .I3(add_rk_out[10]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [18]));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][19]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [19]),
        .I2(\CD[0].col[3][19]_i_2_n_0 ),
        .I3(add_rk_out[11]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [19]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[2].col[1][1]_i_1 
       (.I0(\CD[0].col[3][1]_i_2_n_0 ),
        .I1(\CD[1].col[2][1]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [1]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [1]));
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][20]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [20]),
        .I2(\CD[0].col[3][20]_i_2_n_0 ),
        .I3(add_rk_out[12]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [20]));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][21]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [21]),
        .I2(\CD[0].col[3][21]_i_2_n_0 ),
        .I3(add_rk_out[13]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [21]));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][22]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [22]),
        .I2(\CD[0].col[3][22]_i_2_n_0 ),
        .I3(add_rk_out[14]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [22]));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][23]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][31]_0 [23]),
        .I2(\CD[0].col[3][23]_i_2_n_0 ),
        .I3(add_rk_out[15]),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [23]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[2].col[1][24]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [24]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][24] ),
        .I4(\CD[0].col[3][24]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][31] [24]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[2].col[1][25]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [25]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][25] ),
        .I4(\CD[0].col[3][25]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][31] [25]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[2].col[1][26]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [26]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][26] ),
        .I4(\CD[0].col[3][26]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][31] [26]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[2].col[1][27]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [27]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][27] ),
        .I4(\CD[0].col[3][27]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][31] [27]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[2].col[1][28]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [28]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][28] ),
        .I4(\CD[0].col[3][28]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][31] [28]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[2].col[1][29]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [29]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][29] ),
        .I4(\CD[0].col[3][29]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][31] [29]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[2].col[1][2]_i_1 
       (.I0(\CD[0].col[3][2]_i_2_n_0 ),
        .I1(\CD[1].col[2][2]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [2]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [2]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [2]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[2].col[1][30]_i_1 
       (.I0(\CD[2].col_reg[1][31]_0 [30]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][30] ),
        .I4(\CD[0].col[3][30]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][31] [30]));
  LUT6 #(
    .INIT(64'hE2E2E2E2FFE2E2E2)) 
    \CD[2].col[1][31]_i_1 
       (.I0(\CD[0].col_reg[3][31]_1 [1]),
        .I1(\FSM_sequential_state_reg[2]_5 ),
        .I2(\FSM_sequential_state_reg[2]_2 [1]),
        .I3(\CD[3].col_reg[0][31]_3 ),
        .I4(\CD[3].col_reg[0][31]_2 [0]),
        .I5(\CD[3].col_reg[0][31]_2 [1]),
        .O(\col_en_cnt_unit_pp2_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[2].col[1][31]_i_2 
       (.I0(\CD[2].col_reg[1][31]_0 [31]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[2].col_reg[1][31]_2 ),
        .I4(\CD[0].col[3][31]_i_5_n_0 ),
        .O(\CD[2].col_reg[1][31] [31]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[2].col[1][3]_i_1 
       (.I0(\CD[0].col[3][3]_i_2_n_0 ),
        .I1(\CD[1].col[2][3]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [3]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [3]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [3]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[2].col[1][4]_i_1 
       (.I0(\CD[0].col[3][4]_i_2_n_0 ),
        .I1(\CD[1].col[2][4]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [4]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [4]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [4]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[2].col[1][5]_i_1 
       (.I0(\CD[0].col[3][5]_i_2_n_0 ),
        .I1(\CD[1].col[2][5]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [5]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [5]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [5]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[2].col[1][6]_i_1 
       (.I0(\CD[0].col[3][6]_i_2_n_0 ),
        .I1(\CD[1].col[2][6]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [6]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [6]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [6]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[2].col[1][7]_i_1 
       (.I0(\CD[0].col[3][7]_i_2_n_0 ),
        .I1(\CD[1].col[2][7]_i_2_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\CD[1].col_reg[2][31]_0 [7]),
        .I4(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [7]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [7]));
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][8]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [8]),
        .I2(\CD[0].col[3][8]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][8] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[2].col_reg[1][31] [8]));
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[2].col[1][9]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [9]),
        .I2(\CD[0].col[3][9]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][9] ),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[2].col_reg[1][31] [9]));
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][0]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [0]),
        .I2(\CD[0].col[3][0]_i_2_n_0 ),
        .I3(add_rk_out[0]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [0]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[3].col[0][10]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [10]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][10] ),
        .I4(\CD[0].col[3][10]_i_3_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [10]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[3].col[0][11]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [11]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][11] ),
        .I4(\CD[0].col[3][11]_i_3_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [11]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[3].col[0][12]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [12]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][12] ),
        .I4(\CD[0].col[3][12]_i_3_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [12]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[3].col[0][13]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [13]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][13] ),
        .I4(\CD[0].col[3][13]_i_3_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [13]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[3].col[0][14]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [14]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][14] ),
        .I4(\CD[0].col[3][14]_i_3_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [14]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[3].col[0][15]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [15]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][15] ),
        .I4(\CD[0].col[3][15]_i_5_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [15]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[3].col[0][16]_i_1 
       (.I0(\CD[0].col[3][16]_i_2_n_0 ),
        .I1(\CD[0].col[3][16]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [16]),
        .I4(\CD[2].col_reg[1][31]_0 [16]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [16]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[3].col[0][17]_i_1 
       (.I0(\CD[0].col[3][17]_i_2_n_0 ),
        .I1(\CD[0].col[3][17]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [17]),
        .I4(\CD[2].col_reg[1][31]_0 [17]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [17]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[3].col[0][18]_i_1 
       (.I0(\CD[0].col[3][18]_i_2_n_0 ),
        .I1(\CD[0].col[3][18]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [18]),
        .I4(\CD[2].col_reg[1][31]_0 [18]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [18]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[3].col[0][19]_i_1 
       (.I0(\CD[0].col[3][19]_i_2_n_0 ),
        .I1(\CD[0].col[3][19]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [19]),
        .I4(\CD[2].col_reg[1][31]_0 [19]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [19]));
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][1]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [1]),
        .I2(\CD[0].col[3][1]_i_2_n_0 ),
        .I3(add_rk_out[1]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [1]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[3].col[0][20]_i_1 
       (.I0(\CD[0].col[3][20]_i_2_n_0 ),
        .I1(\CD[0].col[3][20]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [20]),
        .I4(\CD[2].col_reg[1][31]_0 [20]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [20]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[3].col[0][21]_i_1 
       (.I0(\CD[0].col[3][21]_i_2_n_0 ),
        .I1(\CD[0].col[3][21]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [21]),
        .I4(\CD[2].col_reg[1][31]_0 [21]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [21]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[3].col[0][22]_i_1 
       (.I0(\CD[0].col[3][22]_i_2_n_0 ),
        .I1(\CD[0].col[3][22]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [22]),
        .I4(\CD[2].col_reg[1][31]_0 [22]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [22]));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \CD[3].col[0][23]_i_1 
       (.I0(\CD[0].col[3][23]_i_2_n_0 ),
        .I1(\CD[0].col[3][23]_i_3_n_0 ),
        .I2(\CD[0].col[3][31]_i_4_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [23]),
        .I4(\CD[2].col_reg[1][31]_0 [23]),
        .I5(\CD[0].col[3][23]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [23]));
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][24]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [24]),
        .I2(\CD[0].col[3][24]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][24] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [24]));
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][25]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [25]),
        .I2(\CD[0].col[3][25]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][25] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [25]));
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][26]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [26]),
        .I2(\CD[0].col[3][26]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][26] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [26]));
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][27]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [27]),
        .I2(\CD[0].col[3][27]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][27] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [27]));
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][28]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [28]),
        .I2(\CD[0].col[3][28]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][28] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [28]));
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][29]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [29]),
        .I2(\CD[0].col[3][29]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][29] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [29]));
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][2]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [2]),
        .I2(\CD[0].col[3][2]_i_2_n_0 ),
        .I3(add_rk_out[2]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [2]));
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][30]_i_1 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [30]),
        .I2(\CD[0].col[3][30]_i_2_n_0 ),
        .I3(\CD[2].col_reg[1][30] ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [30]));
  LUT6 #(
    .INIT(64'hE2E2E2E2E2E2FFE2)) 
    \CD[3].col[0][31]_i_1 
       (.I0(\CD[0].col_reg[3][31]_1 [0]),
        .I1(\FSM_sequential_state_reg[2]_5 ),
        .I2(\FSM_sequential_state_reg[2]_2 [0]),
        .I3(\CD[3].col_reg[0][31]_3 ),
        .I4(\CD[3].col_reg[0][31]_2 [0]),
        .I5(\CD[3].col_reg[0][31]_2 [1]),
        .O(\col_en_cnt_unit_pp2_reg[0] ));
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][31]_i_2 
       (.I0(\CD[0].col[3][23]_i_4_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [31]),
        .I2(\CD[0].col[3][31]_i_5_n_0 ),
        .I3(\CD[2].col_reg[1][31]_2 ),
        .I4(\CD[0].col[3][7]_i_4_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [31]));
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][3]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [3]),
        .I2(\CD[0].col[3][3]_i_2_n_0 ),
        .I3(add_rk_out[3]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [3]));
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][4]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [4]),
        .I2(\CD[0].col[3][4]_i_2_n_0 ),
        .I3(add_rk_out[4]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [4]));
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][5]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [5]),
        .I2(\CD[0].col[3][5]_i_2_n_0 ),
        .I3(add_rk_out[5]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [5]));
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][6]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [6]),
        .I2(\CD[0].col[3][6]_i_2_n_0 ),
        .I3(add_rk_out[6]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [6]));
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \CD[3].col[0][7]_i_1 
       (.I0(\CD[0].col[3][31]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_0 [7]),
        .I2(\CD[0].col[3][7]_i_2_n_0 ),
        .I3(add_rk_out[7]),
        .I4(\CD[0].col[3][31]_i_7_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [7]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[3].col[0][8]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [8]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][8] ),
        .I4(\CD[0].col[3][8]_i_3_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [8]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \CD[3].col[0][9]_i_1 
       (.I0(\CD[1].col_reg[2][31]_0 [9]),
        .I1(\FSM_sequential_state_reg[0]_2 ),
        .I2(\CD[0].col[3][15]_i_3_n_0 ),
        .I3(\CD[1].col_reg[2][9] ),
        .I4(\CD[0].col[3][9]_i_3_n_0 ),
        .O(\CD[3].col_reg[0][31]_0 [9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \FSM_sequential_state[0]_i_1__0 
       (.I0(\FSM_sequential_state[0]_i_2_n_0 ),
        .I1(\FSM_sequential_state[0]_i_3__0_n_0 ),
        .I2(\FSM_sequential_state_reg[0]_3 ),
        .I3(\FSM_sequential_state[0]_i_5_n_0 ),
        .I4(\FSM_sequential_state[0]_i_6_n_0 ),
        .I5(\FSM_sequential_state[0]_i_7_n_0 ),
        .O(\FSM_sequential_state[0]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hF2F2F2F2FEFFFEFE)) 
    \FSM_sequential_state[0]_i_2 
       (.I0(\FSM_sequential_state_reg[0]_4 ),
        .I1(Q[1]),
        .I2(\FSM_sequential_state[2]_i_3_n_0 ),
        .I3(\info_o[0]_0 [0]),
        .I4(Q[0]),
        .I5(\FSM_sequential_state_reg[3]_2 ),
        .O(\FSM_sequential_state[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h000000000C808080)) 
    \FSM_sequential_state[0]_i_3__0 
       (.I0(Q[3]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(\info_o[0]_0 [1]),
        .I4(\key_en_pp1_reg[3]_0 ),
        .I5(Q[2]),
        .O(\FSM_sequential_state[0]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000444F)) 
    \FSM_sequential_state[0]_i_5 
       (.I0(\key_en_pp1_reg[3]_0 ),
        .I1(Q[2]),
        .I2(\FSM_sequential_state_reg[0]_0 ),
        .I3(\info_o[0]_0 [1]),
        .I4(Q[3]),
        .I5(\rd_count_reg[3]_1 [1]),
        .O(\FSM_sequential_state[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h003000000030B000)) 
    \FSM_sequential_state[0]_i_6 
       (.I0(\FSM_sequential_state_reg[0]_5 ),
        .I1(\key_en_pp1_reg[3]_0 ),
        .I2(Q[2]),
        .I3(Q[1]),
        .I4(Q[0]),
        .I5(\rd_count_reg[3]_0 ),
        .O(\FSM_sequential_state[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000010130000303)) 
    \FSM_sequential_state[0]_i_7 
       (.I0(\key_en_pp1_reg[3]_0 ),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(Q[3]),
        .I4(Q[2]),
        .I5(\info_o[0]_0 [1]),
        .O(\FSM_sequential_state[0]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT5 #(
    .INIT(32'h00F0F808)) 
    \FSM_sequential_state[1]_i_3__0 
       (.I0(Q[2]),
        .I1(\FSM_sequential_state[1]_i_8_n_0 ),
        .I2(Q[0]),
        .I3(Q[1]),
        .I4(Q[3]),
        .O(\FSM_sequential_state_reg[2]_4 ));
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT5 #(
    .INIT(32'hFB000000)) 
    \FSM_sequential_state[1]_i_4__0 
       (.I0(\rd_count_reg[3]_0 ),
        .I1(Q[3]),
        .I2(Q[0]),
        .I3(Q[1]),
        .I4(Q[2]),
        .O(\FSM_sequential_state_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h000000F000008000)) 
    \FSM_sequential_state[1]_i_7 
       (.I0(\key_en_pp1_reg[3]_0 ),
        .I1(\info_o[0]_0 [1]),
        .I2(Q[3]),
        .I3(Q[2]),
        .I4(Q[1]),
        .I5(Q[0]),
        .O(\aes_cr_reg[4] ));
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \FSM_sequential_state[1]_i_8 
       (.I0(\rd_count_reg[3]_1 [2]),
        .I1(\rd_count_reg[3]_1 [1]),
        .I2(\rd_count_reg[3]_1 [3]),
        .I3(\rd_count_reg[3]_1 [0]),
        .O(\FSM_sequential_state[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAAFFBAAAABAABAAA)) 
    \FSM_sequential_state[2]_i_1__0 
       (.I0(\FSM_sequential_state[2]_i_2__0_n_0 ),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(\col_en_cnt_unit_pp1_reg[3] ),
        .I4(Q[0]),
        .I5(Q[1]),
        .O(\FSM_sequential_state[2]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    \FSM_sequential_state[2]_i_2__0 
       (.I0(\FSM_sequential_state_reg[0]_3 ),
        .I1(\FSM_sequential_state[2]_i_3_n_0 ),
        .I2(\FSM_sequential_state_reg[2]_7 ),
        .I3(\FSM_sequential_state_reg[2]_0 ),
        .I4(\FSM_sequential_state_reg[3]_0 ),
        .I5(\FSM_sequential_state[2]_i_5__0_n_0 ),
        .O(\FSM_sequential_state[2]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h01011110FFFFFFFF)) 
    \FSM_sequential_state[2]_i_3 
       (.I0(\FSM_sequential_state_reg[3]_2 ),
        .I1(Q[0]),
        .I2(\rd_count_reg[3]_1 [1]),
        .I3(\rd_count_reg[3]_1 [0]),
        .I4(\rd_count_reg[3]_1 [3]),
        .I5(\FSM_sequential_state_reg[3]_9 ),
        .O(\FSM_sequential_state[2]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT4 #(
    .INIT(16'hFFFB)) 
    \FSM_sequential_state[2]_i_3__0 
       (.I0(Q[2]),
        .I1(Q[3]),
        .I2(Q[0]),
        .I3(Q[1]),
        .O(\FSM_sequential_state_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0800080008030800)) 
    \FSM_sequential_state[2]_i_5__0 
       (.I0(\rd_count_reg[3]_0 ),
        .I1(\col_en_cnt_unit_pp1_reg[3] ),
        .I2(Q[0]),
        .I3(Q[3]),
        .I4(Q[2]),
        .I5(\rd_count_reg[3]_1 [1]),
        .O(\FSM_sequential_state[2]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF4004400)) 
    \FSM_sequential_state[3]_i_1 
       (.I0(\FSM_sequential_state[3]_i_2_n_0 ),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(\FSM_sequential_state_reg[3]_9 ),
        .I4(\FSM_sequential_state_reg[3]_10 ),
        .I5(\FSM_sequential_state[3]_i_4_n_0 ),
        .O(\FSM_sequential_state[3]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \FSM_sequential_state[3]_i_2 
       (.I0(Q[0]),
        .I1(Q[1]),
        .O(\FSM_sequential_state[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hCFDCCCCCCCDCCCCC)) 
    \FSM_sequential_state[3]_i_4 
       (.I0(\FSM_sequential_state_reg[0]_0 ),
        .I1(\FSM_sequential_state[3]_i_5_n_0 ),
        .I2(Q[2]),
        .I3(Q[3]),
        .I4(\FSM_sequential_state_reg[3]_9 ),
        .I5(\FSM_sequential_state_reg[3]_11 ),
        .O(\FSM_sequential_state[3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000800080)) 
    \FSM_sequential_state[3]_i_5 
       (.I0(Q[2]),
        .I1(Q[3]),
        .I2(\FSM_sequential_state_reg[3]_9 ),
        .I3(Q[1]),
        .I4(\col_en_cnt_unit_pp1_reg[3] ),
        .I5(\rd_count_reg[3]_0 ),
        .O(\FSM_sequential_state[3]_i_5_n_0 ));
  (* FSM_ENCODED_STATES = "ROUND0_COL3:0001,ROUND0_COL2:0000,GEN_KEY2:1111,ROUND0_COL1:0010,GEN_KEY1:0111,GEN_KEY0:0110,READY:1000,ROUND0_COL0:0011,IDLE:0101,ROUND_COL1:1001,ROUND_COL3:1100,ROUND_COL2:1010,ROUND_COL0:1011,NOP:1101,GEN_KEY3:1110,ROUND_KEY0:0100" *) 
  FDPE #(
    .INIT(1'b1)) 
    \FSM_sequential_state_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\FSM_sequential_state[0]_i_1__0_n_0 ),
        .PRE(rst_i),
        .Q(Q[0]));
  (* FSM_ENCODED_STATES = "ROUND0_COL3:0001,ROUND0_COL2:0000,GEN_KEY2:1111,ROUND0_COL1:0010,GEN_KEY1:0111,GEN_KEY0:0110,READY:1000,ROUND0_COL0:0011,IDLE:0101,ROUND_COL1:1001,ROUND_COL3:1100,ROUND_COL2:1010,ROUND_COL0:1011,NOP:1101,GEN_KEY3:1110,ROUND_KEY0:0100" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_state_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\FSM_sequential_state_reg[1]_1 ),
        .Q(Q[1]));
  (* FSM_ENCODED_STATES = "ROUND0_COL3:0001,ROUND0_COL2:0000,GEN_KEY2:1111,ROUND0_COL1:0010,GEN_KEY1:0111,GEN_KEY0:0110,READY:1000,ROUND0_COL0:0011,IDLE:0101,ROUND_COL1:1001,ROUND_COL3:1100,ROUND_COL2:1010,ROUND_COL0:1011,NOP:1101,GEN_KEY3:1110,ROUND_KEY0:0100" *) 
  FDPE #(
    .INIT(1'b1)) 
    \FSM_sequential_state_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\FSM_sequential_state[2]_i_1__0_n_0 ),
        .PRE(rst_i),
        .Q(Q[2]));
  (* FSM_ENCODED_STATES = "ROUND0_COL3:0001,ROUND0_COL2:0000,GEN_KEY2:1111,ROUND0_COL1:0010,GEN_KEY1:0111,GEN_KEY0:0110,READY:1000,ROUND0_COL0:0011,IDLE:0101,ROUND_COL1:1001,ROUND_COL3:1100,ROUND_COL2:1010,ROUND_COL0:1011,NOP:1101,GEN_KEY3:1110,ROUND_KEY0:0100" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_state_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\FSM_sequential_state[3]_i_1_n_0 ),
        .Q(Q[3]));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][0]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][0] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [0]),
        .I3(\CD[0].col[3][0]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][0]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [0]));
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][0]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[0]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][16]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][16] ),
        .I1(\CD[0].col[3][16]_i_2_n_0 ),
        .I2(\CD[0].col[3][16]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp[0][16]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][16]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [8]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][16]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [16]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][16]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][16]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [16]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][16]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][17]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][17] ),
        .I1(\CD[0].col[3][17]_i_2_n_0 ),
        .I2(\CD[0].col[3][17]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp[0][17]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][17]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [9]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][17]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [17]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][17]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [17]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][18]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][18] ),
        .I1(\CD[0].col[3][18]_i_2_n_0 ),
        .I2(\CD[0].col[3][18]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp[0][18]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][18]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [10]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][18]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [18]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][18]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [18]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][18]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][19]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][19] ),
        .I1(\CD[0].col[3][19]_i_2_n_0 ),
        .I2(\CD[0].col[3][19]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp[0][19]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][19]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [11]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][19]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [19]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][19]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [19]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][19]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][1]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][1] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [1]),
        .I3(\CD[0].col[3][1]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][1]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [1]));
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][1]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[1]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][20]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][20] ),
        .I1(\CD[0].col[3][20]_i_2_n_0 ),
        .I2(\CD[0].col[3][20]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp[0][20]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][20]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [12]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][20]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [20]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][20]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [20]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][20]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][21]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][21] ),
        .I1(\CD[0].col[3][21]_i_2_n_0 ),
        .I2(\CD[0].col[3][21]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp[0][21]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][21]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [13]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][21]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [21]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][21]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [21]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][22]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][22] ),
        .I1(\CD[0].col[3][22]_i_2_n_0 ),
        .I2(\CD[0].col[3][22]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp[0][22]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][22]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [14]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][22]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [22]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][22]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [22]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][22]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][23]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][23] ),
        .I1(\CD[0].col[3][23]_i_2_n_0 ),
        .I2(\CD[0].col[3][23]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[0].bkp[0][23]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][23]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [15]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][23]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [23]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[0].bkp[0][23]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [23]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][23]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][24]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][24] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [24]),
        .I3(\CD[0].col[3][24]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][24]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [16]));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][24]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[2].col_reg[1][24] ),
        .O(\IV_BKP_REGISTERS[0].bkp[0][24]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][25]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][25] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [25]),
        .I3(\CD[0].col[3][25]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][25]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [17]));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][25]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[2].col_reg[1][25] ),
        .O(\IV_BKP_REGISTERS[0].bkp[0][25]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][26]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][26] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [26]),
        .I3(\CD[0].col[3][26]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][26]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [18]));
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][26]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[2].col_reg[1][26] ),
        .O(\IV_BKP_REGISTERS[0].bkp[0][26]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][27]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][27] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [27]),
        .I3(\CD[0].col[3][27]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][27]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [19]));
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][27]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[2].col_reg[1][27] ),
        .O(\IV_BKP_REGISTERS[0].bkp[0][27]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][28]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][28] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [28]),
        .I3(\CD[0].col[3][28]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][28]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [20]));
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][28]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[2].col_reg[1][28] ),
        .O(\IV_BKP_REGISTERS[0].bkp[0][28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][29]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][29] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [29]),
        .I3(\CD[0].col[3][29]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][29]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [21]));
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][29]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[2].col_reg[1][29] ),
        .O(\IV_BKP_REGISTERS[0].bkp[0][29]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][2]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][2] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [2]),
        .I3(\CD[0].col[3][2]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][2]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [2]));
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][2]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[2]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][30]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][30] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [30]),
        .I3(\CD[0].col[3][30]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][30]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [22]));
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][30]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[2].col_reg[1][30] ),
        .O(\IV_BKP_REGISTERS[0].bkp[0][30]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][31]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [31]),
        .I3(\CD[0].col[3][31]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][31]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [23]));
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][31]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[2].col_reg[1][31]_2 ),
        .O(\IV_BKP_REGISTERS[0].bkp[0][31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][3]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][3] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [3]),
        .I3(\CD[0].col[3][3]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][3]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [3]));
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][3]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[3]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][4]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][4] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [4]),
        .I3(\CD[0].col[3][4]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][4]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [4]));
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][4]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[4]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][5]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][5] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [5]),
        .I3(\CD[0].col[3][5]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][5]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [5]));
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][5]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[5]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][6]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][6] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [6]),
        .I3(\CD[0].col[3][6]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][6]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [6]));
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][6]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[6]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[0].bkp[0][7]_i_1 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][7] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [7]),
        .I3(\CD[0].col[3][7]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp[0][7]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[0].col_reg[3][31] [7]));
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][7]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[7]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][0]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][0] ),
        .I1(\CD[0].col[3][0]_i_2_n_0 ),
        .I2(\CD[1].col[2][0]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[1].bkp[1][0]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][0]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [0]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][0]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [0]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][0]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [0]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][10]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][10] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [10]),
        .I3(\CD[0].col[3][10]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][10]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [10]));
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][10]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][10] ),
        .O(\IV_BKP_REGISTERS[1].bkp[1][10]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][11]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][11] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [11]),
        .I3(\CD[0].col[3][11]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][11]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [11]));
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][11]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][11] ),
        .O(\IV_BKP_REGISTERS[1].bkp[1][11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][12]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][12] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [12]),
        .I3(\CD[0].col[3][12]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][12]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [12]));
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][12]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][12] ),
        .O(\IV_BKP_REGISTERS[1].bkp[1][12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][13]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][13] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [13]),
        .I3(\CD[0].col[3][13]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][13]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [13]));
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][13]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][13] ),
        .O(\IV_BKP_REGISTERS[1].bkp[1][13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][14]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][14] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [14]),
        .I3(\CD[0].col[3][14]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][14]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [14]));
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][14]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][14] ),
        .O(\IV_BKP_REGISTERS[1].bkp[1][14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][15]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][15] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [15]),
        .I3(\CD[0].col[3][15]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][15]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [15]));
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][15]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][15] ),
        .O(\IV_BKP_REGISTERS[1].bkp[1][15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][16]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][16] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [16]),
        .I3(\CD[0].col[3][16]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][16]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [16]));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][16]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[8]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][16]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][17]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][17] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [17]),
        .I3(\CD[0].col[3][17]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][17]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [17]));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][17]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[9]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][18]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][18] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [18]),
        .I3(\CD[0].col[3][18]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][18]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [18]));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][18]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[10]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][19]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][19] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [19]),
        .I3(\CD[0].col[3][19]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][19]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [19]));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][19]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[11]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][1]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][1] ),
        .I1(\CD[0].col[3][1]_i_2_n_0 ),
        .I2(\CD[1].col[2][1]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[1].bkp[1][1]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][1]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [1]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][1]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [1]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][1]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [1]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][20]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][20] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [20]),
        .I3(\CD[0].col[3][20]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][20]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [20]));
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][20]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[12]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][21]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][21] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [21]),
        .I3(\CD[0].col[3][21]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][21]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [21]));
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][21]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[13]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][22]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][22] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [22]),
        .I3(\CD[0].col[3][22]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][22]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [22]));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][22]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[14]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][23]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][23] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [23]),
        .I3(\CD[0].col[3][23]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][23]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [23]));
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][23]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[15]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][2]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][2] ),
        .I1(\CD[0].col[3][2]_i_2_n_0 ),
        .I2(\CD[1].col[2][2]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[1].bkp[1][2]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][2]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [2]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][2]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [2]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][2]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [2]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][3]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][3] ),
        .I1(\CD[0].col[3][3]_i_2_n_0 ),
        .I2(\CD[1].col[2][3]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[1].bkp[1][3]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][3]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [3]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][3]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [3]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][3]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [3]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][4]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][4] ),
        .I1(\CD[0].col[3][4]_i_2_n_0 ),
        .I2(\CD[1].col[2][4]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[1].bkp[1][4]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][4]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [4]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][4]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [4]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][4]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [4]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][5]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][5] ),
        .I1(\CD[0].col[3][5]_i_2_n_0 ),
        .I2(\CD[1].col[2][5]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[1].bkp[1][5]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][5]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [5]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][5]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [5]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][5]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [5]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][6]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][6] ),
        .I1(\CD[0].col[3][6]_i_2_n_0 ),
        .I2(\CD[1].col[2][6]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[1].bkp[1][6]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][6]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [6]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][6]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [6]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][6]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [6]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][7]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][7] ),
        .I1(\CD[0].col[3][7]_i_2_n_0 ),
        .I2(\CD[1].col[2][7]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[1].bkp[1][7]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][7]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [7]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][7]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [7]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[1].bkp[1][7]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [7]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][8]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][8] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [8]),
        .I3(\CD[0].col[3][8]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][8]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [8]));
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][8]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][8] ),
        .O(\IV_BKP_REGISTERS[1].bkp[1][8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[1].bkp[1][9]_i_1 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][9] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [9]),
        .I3(\CD[0].col[3][9]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp[1][9]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[2].col_reg[1][23] [9]));
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][9]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[1].col_reg[2][9] ),
        .O(\IV_BKP_REGISTERS[1].bkp[1][9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][0]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][0] ),
        .I1(\CD[0].col[3][0]_i_2_n_0 ),
        .I2(\CD[1].col[2][0]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][0]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][0]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [0]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][0]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [0]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][0]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [0]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][10]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][10] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [10]),
        .I3(\CD[0].col[3][10]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][10]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [10]));
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][10]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[1].col_reg[2][10] ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][10]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][11]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][11] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [11]),
        .I3(\CD[0].col[3][11]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][11]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [11]));
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][11]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[1].col_reg[2][11] ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][12]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][12] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [12]),
        .I3(\CD[0].col[3][12]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][12]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [12]));
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][12]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[1].col_reg[2][12] ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][13]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][13] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [13]),
        .I3(\CD[0].col[3][13]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][13]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [13]));
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][13]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[1].col_reg[2][13] ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][14]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][14] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [14]),
        .I3(\CD[0].col[3][14]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][14]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [14]));
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][14]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[1].col_reg[2][14] ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][15]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][15] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [15]),
        .I3(\CD[0].col[3][15]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][15]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [15]));
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][15]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[1].col_reg[2][15] ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][16]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][16] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [16]),
        .I3(\CD[0].col[3][16]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][16]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [16]));
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][16]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[8]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][16]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][17]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][17] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [17]),
        .I3(\CD[0].col[3][17]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][17]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [17]));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][17]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[9]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][18]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][18] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [18]),
        .I3(\CD[0].col[3][18]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][18]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [18]));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][18]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[10]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][19]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][19] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [19]),
        .I3(\CD[0].col[3][19]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][19]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [19]));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][19]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[11]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][1]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][1] ),
        .I1(\CD[0].col[3][1]_i_2_n_0 ),
        .I2(\CD[1].col[2][1]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][1]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][1]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [1]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][1]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [1]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][1]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [1]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][20]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][20] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [20]),
        .I3(\CD[0].col[3][20]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][20]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [20]));
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][20]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[12]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][21]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][21] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [21]),
        .I3(\CD[0].col[3][21]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][21]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [21]));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][21]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[13]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][22]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][22] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [22]),
        .I3(\CD[0].col[3][22]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][22]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [22]));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][22]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[14]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][23]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][23] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\CD[1].col_reg[2][31]_0 [23]),
        .I3(\CD[0].col[3][23]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][23]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [23]));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][23]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(add_rk_out[15]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[2].bkp[2][24]_i_6 
       (.I0(\CD[0].col[3][5]_i_2_2 ),
        .I1(\info_o[24]_INST_0_i_6_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [20]),
        .I4(\info_o[31]_2 [24]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][24] ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[2].bkp[2][25]_i_6 
       (.I0(\CD[0].col[3][5]_i_2_2 ),
        .I1(\info_o[25]_INST_0_i_6_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [21]),
        .I4(\info_o[31]_2 [25]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][25] ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[2].bkp[2][26]_i_6 
       (.I0(\CD[0].col[3][5]_i_2_2 ),
        .I1(\info_o[26]_INST_0_i_6_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [22]),
        .I4(\info_o[31]_2 [26]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][26] ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[2].bkp[2][27]_i_6 
       (.I0(\CD[0].col[3][5]_i_2_2 ),
        .I1(\info_o[27]_INST_0_i_6_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [23]),
        .I4(\info_o[31]_2 [27]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][27] ));
  LUT6 #(
    .INIT(64'hFEFEFEEFEEEEEEEE)) 
    \IV_BKP_REGISTERS[2].bkp[2][28]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp[2][28]_i_5_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp[2][28]_i_6_n_0 ),
        .I2(\CD[2].col_reg[1][28]_1 ),
        .I3(\CD[2].col_reg[1][28]_0 ),
        .I4(\CD[0].col[3][28]_i_4_n_0 ),
        .I5(\CD[2].col_reg[1][31]_1 ),
        .O(data_in[4]));
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][28]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[28]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][28]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[2].bkp[2][28]_i_6 
       (.I0(\CD[0].col[3][31]_i_27_n_0 ),
        .I1(\info_o[28]_INST_0_i_8_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [24]),
        .I4(\info_o[31]_2 [28]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][28]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[2].bkp[2][29]_i_6 
       (.I0(\CD[0].col[3][5]_i_2_2 ),
        .I1(\info_o[29]_INST_0_i_8_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [25]),
        .I4(\info_o[31]_2 [29]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][29] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][2]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][2] ),
        .I1(\CD[0].col[3][2]_i_2_n_0 ),
        .I2(\CD[1].col[2][2]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][2]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][2]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [2]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][2]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [2]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][2]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [2]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[2].bkp[2][30]_i_6 
       (.I0(\CD[0].col[3][5]_i_2_2 ),
        .I1(\info_o[30]_INST_0_i_8_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [26]),
        .I4(\info_o[31]_2 [30]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][30] ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[2].bkp[2][31]_i_6 
       (.I0(\CD[0].col[3][5]_i_2_2 ),
        .I1(\info_o[31]_INST_0_i_16_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [27]),
        .I4(\info_o[31]_2 [31]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][31] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][3]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][3] ),
        .I1(\CD[0].col[3][3]_i_2_n_0 ),
        .I2(\CD[1].col[2][3]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][3]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][3]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [3]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][3]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [3]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][3]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [3]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][4]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][4] ),
        .I1(\CD[0].col[3][4]_i_2_n_0 ),
        .I2(\CD[1].col[2][4]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][4]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][4]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [4]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][4]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [4]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][4]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [4]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][5]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][5] ),
        .I1(\CD[0].col[3][5]_i_2_n_0 ),
        .I2(\CD[1].col[2][5]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][5]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][5]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [5]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][5]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [5]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][5]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [5]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][6]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][6] ),
        .I1(\CD[0].col[3][6]_i_2_n_0 ),
        .I2(\CD[1].col[2][6]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][6]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][6]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [6]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][6]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [6]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][6]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [6]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][7]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][7] ),
        .I1(\CD[0].col[3][7]_i_2_n_0 ),
        .I2(\CD[1].col[2][7]_i_2_n_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][7]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][7]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [7]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][7]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[1].col_reg[2][31]_0 [7]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[2].bkp[2][7]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [7]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][8]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][8] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [8]),
        .I3(\CD[0].col[3][8]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][8]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [8]));
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][8]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[1].col_reg[2][8] ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][9]_i_1 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][9] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [9]),
        .I3(\CD[0].col[3][9]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][9]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[1].col_reg[2][23] [9]));
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][9]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(\CD[1].col_reg[2][9] ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][0]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][0] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [0]),
        .I3(\CD[0].col[3][0]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][0]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [0]));
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][0]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[0]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEEFEEEEEEEE)) 
    \IV_BKP_REGISTERS[3].bkp[3][10]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][10]_i_5_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][10]_i_6_n_0 ),
        .I2(\CD[1].col_reg[2][10]_1 ),
        .I3(\CD[1].col_reg[2][10]_0 ),
        .I4(\CD[0].col[3][10]_i_6_n_0 ),
        .I5(\CD[2].col_reg[1][31]_1 ),
        .O(data_in[0]));
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][10]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[10]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][10]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[3].bkp[3][10]_i_6 
       (.I0(\CD[0].col[3][31]_i_27_n_0 ),
        .I1(\info_o[10]_INST_0_i_4_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [6]),
        .I4(\info_o[31]_2 [10]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEEFEEEEEEEE)) 
    \IV_BKP_REGISTERS[3].bkp[3][11]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][11]_i_5_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][11]_i_6_n_0 ),
        .I2(\CD[1].col_reg[2][11]_1 ),
        .I3(\CD[1].col_reg[2][11]_0 ),
        .I4(\CD[0].col[3][11]_i_6_n_0 ),
        .I5(\CD[2].col_reg[1][31]_1 ),
        .O(data_in[1]));
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][11]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[11]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[3].bkp[3][11]_i_6 
       (.I0(\CD[0].col[3][31]_i_27_n_0 ),
        .I1(\info_o[11]_INST_0_i_4_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [7]),
        .I4(\info_o[31]_2 [11]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEEFEEEEEEEE)) 
    \IV_BKP_REGISTERS[3].bkp[3][12]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][12]_i_5_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][12]_i_6_n_0 ),
        .I2(\CD[1].col_reg[2][12]_1 ),
        .I3(\CD[1].col_reg[2][12]_0 ),
        .I4(\CD[0].col[3][12]_i_6_n_0 ),
        .I5(\CD[2].col_reg[1][31]_1 ),
        .O(data_in[2]));
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][12]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[12]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][12]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[3].bkp[3][12]_i_6 
       (.I0(\CD[0].col[3][31]_i_27_n_0 ),
        .I1(\info_o[12]_INST_0_i_4_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [8]),
        .I4(\info_o[31]_2 [12]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][12]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEEFEEEEEEEE)) 
    \IV_BKP_REGISTERS[3].bkp[3][13]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_5_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][13]_i_6_n_0 ),
        .I2(\CD[1].col_reg[2][13]_1 ),
        .I3(\CD[1].col_reg[2][13]_0 ),
        .I4(\CD[0].col[3][13]_i_6_n_0 ),
        .I5(\CD[2].col_reg[1][31]_1 ),
        .O(data_in[3]));
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][13]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ),
        .I1(bus_swap[13]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][13]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[3].bkp[3][13]_i_6 
       (.I0(\CD[0].col[3][31]_i_27_n_0 ),
        .I1(\info_o[13]_INST_0_i_4_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [9]),
        .I4(\info_o[31]_2 [13]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00002A00FFFF)) 
    \IV_BKP_REGISTERS[3].bkp[3][13]_i_8 
       (.I0(\rd_count_reg[3]_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(\info_o[0]_0 [1]),
        .I4(\info_o[0]_0 [2]),
        .I5(\info_o[0]_0 [3]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[3].bkp[3][14]_i_6 
       (.I0(\CD[0].col[3][5]_i_2_2 ),
        .I1(\info_o[14]_INST_0_i_4_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [10]),
        .I4(\info_o[31]_2 [14]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][14] ));
  LUT6 #(
    .INIT(64'h0000001500000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][15]_i_11 
       (.I0(\col_en_cnt_unit_pp2_reg[3] ),
        .I1(\key_en_pp1_reg[3]_0 ),
        .I2(first_block),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(first_block_reg_0));
  LUT6 #(
    .INIT(64'h0808000800080008)) 
    \IV_BKP_REGISTERS[3].bkp[3][15]_i_3 
       (.I0(\CD[0].col[3][31]_i_8_n_0 ),
        .I1(\info_o[0]_0 [2]),
        .I2(\info_o[0]_0 [3]),
        .I3(\info_o[0]_0 [1]),
        .I4(Q[1]),
        .I5(Q[2]),
        .O(\aes_cr_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[3].bkp[3][15]_i_8 
       (.I0(\CD[0].col[3][5]_i_2_2 ),
        .I1(\info_o[15]_INST_0_i_4_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [11]),
        .I4(\info_o[31]_2 [15]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][15] ));
  LUT6 #(
    .INIT(64'h0808000800080008)) 
    \IV_BKP_REGISTERS[3].bkp[3][15]_i_9 
       (.I0(\CD[0].col[3][15]_i_3_n_0 ),
        .I1(\info_o[0]_0 [2]),
        .I2(\info_o[0]_0 [3]),
        .I3(\info_o[0]_0 [1]),
        .I4(Q[1]),
        .I5(Q[2]),
        .O(\aes_cr_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][16]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][16] ),
        .I1(\CD[0].col[3][16]_i_2_n_0 ),
        .I2(\CD[0].col[3][16]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][16]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][16]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [8]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][16]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [16]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][16]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][16]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [16]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][16]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][17]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][17] ),
        .I1(\CD[0].col[3][17]_i_2_n_0 ),
        .I2(\CD[0].col[3][17]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][17]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][17]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [9]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][17]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [17]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][17]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [17]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][18]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][18] ),
        .I1(\CD[0].col[3][18]_i_2_n_0 ),
        .I2(\CD[0].col[3][18]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][18]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][18]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [10]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][18]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [18]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][18]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [18]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][18]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][19]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][19] ),
        .I1(\CD[0].col[3][19]_i_2_n_0 ),
        .I2(\CD[0].col[3][19]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][19]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][19]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [11]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][19]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [19]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][19]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [19]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][19]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][1]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][1] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [1]),
        .I3(\CD[0].col[3][1]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][1]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [1]));
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][1]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[1]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][20]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][20] ),
        .I1(\CD[0].col[3][20]_i_2_n_0 ),
        .I2(\CD[0].col[3][20]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][20]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][20]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [12]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][20]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [20]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][20]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [20]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][20]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][21]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][21] ),
        .I1(\CD[0].col[3][21]_i_2_n_0 ),
        .I2(\CD[0].col[3][21]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][21]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][21]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [13]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][21]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [21]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][21]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [21]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][22]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][22] ),
        .I1(\CD[0].col[3][22]_i_2_n_0 ),
        .I2(\CD[0].col[3][22]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][22]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][22]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [14]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][22]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [22]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][22]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [22]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][22]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][23]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][23] ),
        .I1(\CD[0].col[3][23]_i_2_n_0 ),
        .I2(\CD[0].col[3][23]_i_3_n_0 ),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][23]_i_3_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][23]_i_4_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [15]));
  LUT6 #(
    .INIT(64'h7000000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][23]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [23]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF000000000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][23]_i_4 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(\info_o[0]_0 [1]),
        .I3(\key_en_pp1_reg[3]_0 ),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(\CD[2].col_reg[1][31]_0 [23]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][23]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][24]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][24] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [24]),
        .I3(\CD[0].col[3][24]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][24]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [16]));
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][24]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][24] ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][24]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][25]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][25] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [25]),
        .I3(\CD[0].col[3][25]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][25]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [17]));
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][25]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][25] ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][25]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][26]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][26] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [26]),
        .I3(\CD[0].col[3][26]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][26]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [18]));
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][26]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][26] ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][26]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][27]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][27] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [27]),
        .I3(\CD[0].col[3][27]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][27]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [19]));
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][27]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][27] ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][27]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][28]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][28] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [28]),
        .I3(\CD[0].col[3][28]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][28]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [20]));
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][28]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][28] ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][29]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][29] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [29]),
        .I3(\CD[0].col[3][29]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][29]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [21]));
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][29]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][29] ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][29]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][2]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][2] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [2]),
        .I3(\CD[0].col[3][2]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][2]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [2]));
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][2]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[2]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][30]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][30] ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [30]),
        .I3(\CD[0].col[3][30]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][30]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [22]));
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][30]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][30] ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][30]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][31]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 ),
        .I1(\CD[0].col[3][23]_i_4_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [31]),
        .I3(\CD[0].col[3][31]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [23]));
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][31]_i_3 
       (.I0(\CD[0].col[3][7]_i_4_n_0 ),
        .I1(\CD[2].col_reg[1][31]_2 ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][3]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][3] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [3]),
        .I3(\CD[0].col[3][3]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][3]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [3]));
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][3]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[3]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][4]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][4] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [4]),
        .I3(\CD[0].col[3][4]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][4]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [4]));
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][4]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[4]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][5]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][5] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [5]),
        .I3(\CD[0].col[3][5]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][5]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [5]));
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][5]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[5]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][6]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][6] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [6]),
        .I3(\CD[0].col[3][6]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][6]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [6]));
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][6]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[6]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][7]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][7] ),
        .I1(\CD[0].col[3][31]_i_4_n_0 ),
        .I2(\CD[2].col_reg[1][31]_0 [7]),
        .I3(\CD[0].col[3][7]_i_2_n_0 ),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][7]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_reg[3][31] ),
        .O(\CD[3].col_reg[0][31] [7]));
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][7]_i_3 
       (.I0(\CD[0].col[3][31]_i_7_n_0 ),
        .I1(add_rk_out[7]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[3].bkp[3][8]_i_6 
       (.I0(\CD[0].col[3][5]_i_2_2 ),
        .I1(\info_o[8]_INST_0_i_4_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [4]),
        .I4(\info_o[31]_2 [8]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][8] ));
  LUT6 #(
    .INIT(64'hAAAAA888A888A888)) 
    \IV_BKP_REGISTERS[3].bkp[3][9]_i_6 
       (.I0(\CD[0].col[3][5]_i_2_2 ),
        .I1(\info_o[9]_INST_0_i_4_n_0 ),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [5]),
        .I4(\info_o[31]_2 [9]),
        .I5(\info_o[31]_INST_0_i_14_n_0 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][9] ));
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'h8B)) 
    \IV_BKP_REGISTERS[3].iv[3][0]_i_1 
       (.I0(enable_i[0]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\info_o[31]_3 [0]),
        .O(\enable_i[31] [0]));
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][10]_i_1 
       (.I0(enable_i[10]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][16] [1]),
        .O(\enable_i[31] [10]));
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][11]_i_1 
       (.I0(enable_i[11]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][16] [2]),
        .O(\enable_i[31] [11]));
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][12]_i_1 
       (.I0(enable_i[12]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][16] [3]),
        .O(\enable_i[31] [12]));
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][13]_i_1 
       (.I0(enable_i[13]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][16] [4]),
        .O(\enable_i[31] [13]));
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][14]_i_1 
       (.I0(enable_i[14]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][16] [5]),
        .O(\enable_i[31] [14]));
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][15]_i_1 
       (.I0(enable_i[15]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][16] [6]),
        .O(\enable_i[31] [15]));
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][16]_i_1 
       (.I0(enable_i[16]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][16] [7]),
        .O(\enable_i[31] [16]));
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][17]_i_1 
       (.I0(enable_i[17]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][24]_0 [0]),
        .O(\enable_i[31] [17]));
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][18]_i_1 
       (.I0(enable_i[18]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][24]_0 [1]),
        .O(\enable_i[31] [18]));
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][19]_i_1 
       (.I0(enable_i[19]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][24]_0 [2]),
        .O(\enable_i[31] [19]));
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][1]_i_1 
       (.I0(enable_i[1]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][8]_0 [0]),
        .O(\enable_i[31] [1]));
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][20]_i_1 
       (.I0(enable_i[20]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][24]_0 [3]),
        .O(\enable_i[31] [20]));
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][21]_i_1 
       (.I0(enable_i[21]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][24]_0 [4]),
        .O(\enable_i[31] [21]));
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][22]_i_1 
       (.I0(enable_i[22]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][24]_0 [5]),
        .O(\enable_i[31] [22]));
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][23]_i_1 
       (.I0(enable_i[23]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][24]_0 [6]),
        .O(\enable_i[31] [23]));
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][24]_i_1 
       (.I0(enable_i[24]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][24]_0 [7]),
        .O(\enable_i[31] [24]));
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][25]_i_1 
       (.I0(enable_i[25]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(O[0]),
        .O(\enable_i[31] [25]));
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][26]_i_1 
       (.I0(enable_i[26]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(O[1]),
        .O(\enable_i[31] [26]));
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][27]_i_1 
       (.I0(enable_i[27]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(O[2]),
        .O(\enable_i[31] [27]));
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][28]_i_1 
       (.I0(enable_i[28]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(O[3]),
        .O(\enable_i[31] [28]));
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][29]_i_1 
       (.I0(enable_i[29]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(O[4]),
        .O(\enable_i[31] [29]));
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][2]_i_1 
       (.I0(enable_i[2]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][8]_0 [1]),
        .O(\enable_i[31] [2]));
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][30]_i_1 
       (.I0(enable_i[30]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(O[5]),
        .O(\enable_i[31] [30]));
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][31]_i_2 
       (.I0(enable_i[31]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(O[6]),
        .O(\enable_i[31] [31]));
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \IV_BKP_REGISTERS[3].iv[3][31]_i_5 
       (.I0(Q[3]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(\FSM_sequential_state_reg[3]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF7)) 
    \IV_BKP_REGISTERS[3].iv[3][31]_i_6 
       (.I0(Q[3]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\rd_count_reg[3]_0 ),
        .I5(\key_en_pp1_reg[3]_0 ),
        .O(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][3]_i_1 
       (.I0(enable_i[3]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][8]_0 [2]),
        .O(\enable_i[31] [3]));
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][4]_i_1 
       (.I0(enable_i[4]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][8]_0 [3]),
        .O(\enable_i[31] [4]));
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][5]_i_1 
       (.I0(enable_i[5]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][8]_0 [4]),
        .O(\enable_i[31] [5]));
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][6]_i_1 
       (.I0(enable_i[6]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][8]_0 [5]),
        .O(\enable_i[31] [6]));
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][7]_i_1 
       (.I0(enable_i[7]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][8]_0 [6]),
        .O(\enable_i[31] [7]));
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][8]_i_1 
       (.I0(enable_i[8]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][8]_0 [7]),
        .O(\enable_i[31] [8]));
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \IV_BKP_REGISTERS[3].iv[3][9]_i_1 
       (.I0(enable_i[9]),
        .I1(\IV_BKP_REGISTERS[3].iv[3][31]_i_6_n_0 ),
        .I2(\IV_BKP_REGISTERS[3].iv_reg[3][16] [0]),
        .O(\enable_i[31] [9]));
  LUT5 #(
    .INIT(32'hFFFFE2FF)) 
    \KR[0].key[3][31]_i_1 
       (.I0(\KR[0].key_reg[3][31] [3]),
        .I1(bypass_key_en),
        .I2(\FSM_sequential_state_reg[0]_1 [3]),
        .I3(\KR[3].key_reg[0][31]_0 ),
        .I4(key_en[3]),
        .O(\key_en_pp1_reg[3] ));
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT4 #(
    .INIT(16'hC08F)) 
    \KR[0].key[3][31]_i_3 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(Q[3]),
        .O(bypass_key_en));
  LUT6 #(
    .INIT(64'hFFFFFF15F000C015)) 
    \KR[0].key[3][31]_i_5 
       (.I0(\col_en_cnt_unit_pp1_reg[3] ),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(Q[3]),
        .I5(key_sel_pp1),
        .O(key_sel_mux));
  LUT5 #(
    .INIT(32'hFFFFE2FF)) 
    \KR[1].key[2][31]_i_1 
       (.I0(\KR[0].key_reg[3][31] [2]),
        .I1(bypass_key_en),
        .I2(\FSM_sequential_state_reg[0]_1 [2]),
        .I3(\KR[3].key_reg[0][31]_0 ),
        .I4(key_en[2]),
        .O(\key_en_pp1_reg[2] ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][0]_i_1 
       (.I0(\KR[2].key[1][0]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(p_86_in_15),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[96]),
        .I5(key_in[64]),
        .O(\KR[3].key_reg[0][31] [0]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][0]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[0]),
        .I3(\KR[2].key_reg[1][31] [0]),
        .O(\KR[2].key[1][0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][10]_i_1 
       (.I0(\KR[2].key[1][10]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(sbox_out_enc[2]),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[106]),
        .I5(key_in[74]),
        .O(\KR[3].key_reg[0][31] [10]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][10]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[10]),
        .I3(\KR[2].key_reg[1][31] [10]),
        .O(\KR[2].key[1][10]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][11]_i_1 
       (.I0(\KR[2].key[1][11]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(sbox_out_enc[3]),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[107]),
        .I5(key_in[75]),
        .O(\KR[3].key_reg[0][31] [11]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][11]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[11]),
        .I3(\KR[2].key_reg[1][31] [11]),
        .O(\KR[2].key[1][11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][12]_i_1 
       (.I0(\KR[2].key[1][12]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(isomorphism_inv_return03_out_7),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[108]),
        .I5(key_in[76]),
        .O(\KR[3].key_reg[0][31] [12]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][12]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[12]),
        .I3(\KR[2].key_reg[1][31] [12]),
        .O(\KR[2].key[1][12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][13]_i_1 
       (.I0(\KR[2].key[1][13]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(p_93_in_10),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[109]),
        .I5(key_in[77]),
        .O(\KR[3].key_reg[0][31] [13]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][13]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[13]),
        .I3(\KR[2].key_reg[1][31] [13]),
        .O(\KR[2].key[1][13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][14]_i_1 
       (.I0(\KR[2].key[1][14]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(isomorphism_inv_return033_out_6),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[110]),
        .I5(key_in[78]),
        .O(\KR[3].key_reg[0][31] [14]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][14]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[14]),
        .I3(\KR[2].key_reg[1][31] [14]),
        .O(\KR[2].key[1][14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][15]_i_1 
       (.I0(\KR[2].key[1][15]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(isomorphism_inv_return05_out_8),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[111]),
        .I5(key_in[79]),
        .O(\KR[3].key_reg[0][31] [15]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][15]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[15]),
        .I3(\KR[2].key_reg[1][31] [15]),
        .O(\KR[2].key[1][15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][16]_i_1 
       (.I0(\KR[2].key[1][16]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(p_86_in),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[112]),
        .I5(key_in[80]),
        .O(\KR[3].key_reg[0][31] [16]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][16]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[16]),
        .I3(\KR[2].key_reg[1][31] [16]),
        .O(\KR[2].key[1][16]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][17]_i_1 
       (.I0(\KR[2].key[1][17]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(p_16_in),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[113]),
        .I5(key_in[81]),
        .O(\KR[3].key_reg[0][31] [17]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][17]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[17]),
        .I3(\KR[2].key_reg[1][31] [17]),
        .O(\KR[2].key[1][17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][18]_i_1 
       (.I0(\KR[2].key[1][18]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(sbox_out_enc[4]),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[114]),
        .I5(key_in[82]),
        .O(\KR[3].key_reg[0][31] [18]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][18]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[18]),
        .I3(\KR[2].key_reg[1][31] [18]),
        .O(\KR[2].key[1][18]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][19]_i_1 
       (.I0(\KR[2].key[1][19]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(sbox_out_enc[5]),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[115]),
        .I5(key_in[83]),
        .O(\KR[3].key_reg[0][31] [19]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][19]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[19]),
        .I3(\KR[2].key_reg[1][31] [19]),
        .O(\KR[2].key[1][19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][1]_i_1 
       (.I0(\KR[2].key[1][1]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(p_16_in_17),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[97]),
        .I5(key_in[65]),
        .O(\KR[3].key_reg[0][31] [1]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][1]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[1]),
        .I3(\KR[2].key_reg[1][31] [1]),
        .O(\KR[2].key[1][1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][20]_i_1 
       (.I0(\KR[2].key[1][20]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(isomorphism_inv_return03_out),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[116]),
        .I5(key_in[84]),
        .O(\KR[3].key_reg[0][31] [20]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][20]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[20]),
        .I3(\KR[2].key_reg[1][31] [20]),
        .O(\KR[2].key[1][20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][21]_i_1 
       (.I0(\KR[2].key[1][21]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(p_93_in),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[117]),
        .I5(key_in[85]),
        .O(\KR[3].key_reg[0][31] [21]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][21]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[21]),
        .I3(\KR[2].key_reg[1][31] [21]),
        .O(\KR[2].key[1][21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][22]_i_1 
       (.I0(\KR[2].key[1][22]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(isomorphism_inv_return033_out),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[118]),
        .I5(key_in[86]),
        .O(\KR[3].key_reg[0][31] [22]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][22]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[22]),
        .I3(\KR[2].key_reg[1][31] [22]),
        .O(\KR[2].key[1][22]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][23]_i_1 
       (.I0(\KR[2].key[1][23]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(isomorphism_inv_return05_out),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[119]),
        .I5(key_in[87]),
        .O(\KR[3].key_reg[0][31] [23]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][23]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[23]),
        .I3(\KR[2].key_reg[1][31] [23]),
        .O(\KR[2].key[1][23]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][24]_i_1 
       (.I0(\KR[2].key[1][24]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(\KR[2].key_reg[1][24] ),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[120]),
        .I5(key_in[88]),
        .O(\KR[3].key_reg[0][31] [24]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][24]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[24]),
        .I3(\KR[2].key_reg[1][31] [24]),
        .O(\KR[2].key[1][24]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][25]_i_1 
       (.I0(\KR[2].key[1][25]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(\KR[2].key_reg[1][25] ),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[121]),
        .I5(key_in[89]),
        .O(\KR[3].key_reg[0][31] [25]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][25]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[25]),
        .I3(\KR[2].key_reg[1][31] [25]),
        .O(\KR[2].key[1][25]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][26]_i_1 
       (.I0(\KR[2].key[1][26]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(g_func[0]),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[122]),
        .I5(key_in[90]),
        .O(\KR[3].key_reg[0][31] [26]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][26]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[26]),
        .I3(\KR[2].key_reg[1][31] [26]),
        .O(\KR[2].key[1][26]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][27]_i_1 
       (.I0(\KR[2].key[1][27]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(g_func[1]),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[123]),
        .I5(key_in[91]),
        .O(\KR[3].key_reg[0][31] [27]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][27]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[27]),
        .I3(\KR[2].key_reg[1][31] [27]),
        .O(\KR[2].key[1][27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][28]_i_1 
       (.I0(\KR[2].key[1][28]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(\KR[2].key_reg[1][28] ),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[124]),
        .I5(key_in[92]),
        .O(\KR[3].key_reg[0][31] [28]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][28]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[28]),
        .I3(\KR[2].key_reg[1][31] [28]),
        .O(\KR[2].key[1][28]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][29]_i_1 
       (.I0(\KR[2].key[1][29]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(\KR[2].key_reg[1][29] ),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[125]),
        .I5(key_in[93]),
        .O(\KR[3].key_reg[0][31] [29]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][29]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[29]),
        .I3(\KR[2].key_reg[1][31] [29]),
        .O(\KR[2].key[1][29]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][2]_i_1 
       (.I0(\KR[2].key[1][2]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(sbox_out_enc[0]),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[98]),
        .I5(key_in[66]),
        .O(\KR[3].key_reg[0][31] [2]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][2]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[2]),
        .I3(\KR[2].key_reg[1][31] [2]),
        .O(\KR[2].key[1][2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][30]_i_1 
       (.I0(\KR[2].key[1][30]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(\KR[2].key_reg[1][30] ),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[126]),
        .I5(key_in[94]),
        .O(\KR[3].key_reg[0][31] [30]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][30]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[30]),
        .I3(\KR[2].key_reg[1][31] [30]),
        .O(\KR[2].key[1][30]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFE2FF)) 
    \KR[2].key[1][31]_i_1 
       (.I0(\KR[0].key_reg[3][31] [1]),
        .I1(bypass_key_en),
        .I2(\FSM_sequential_state_reg[0]_1 [1]),
        .I3(\KR[3].key_reg[0][31]_0 ),
        .I4(key_en[1]),
        .O(\key_en_pp1_reg[1] ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][31]_i_2 
       (.I0(\KR[2].key[1][31]_i_3_n_0 ),
        .I1(key_sel_mux),
        .I2(\KR[2].key_reg[1][31]_0 ),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[127]),
        .I5(key_in[95]),
        .O(\KR[3].key_reg[0][31] [31]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][31]_i_3 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[31]),
        .I3(\KR[2].key_reg[1][31] [31]),
        .O(\KR[2].key[1][31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEEEE000005550555)) 
    \KR[2].key[1][31]_i_5 
       (.I0(Q[3]),
        .I1(Q[0]),
        .I2(\key_en_pp1_reg[3]_0 ),
        .I3(\info_o[0]_0 [1]),
        .I4(Q[1]),
        .I5(Q[2]),
        .O(\AES_CORE_DATAPATH/key1_mux_cnt ));
  LUT6 #(
    .INIT(64'hEAAAAEEEAEEEEAAA)) 
    \KR[2].key[1][3]_i_1 
       (.I0(\KR[2].key[1][3]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(sbox_out_enc[1]),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[99]),
        .I5(key_in[67]),
        .O(\KR[3].key_reg[0][31] [3]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][3]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[3]),
        .I3(\KR[2].key_reg[1][31] [3]),
        .O(\KR[2].key[1][3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][4]_i_1 
       (.I0(\KR[2].key[1][4]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(isomorphism_inv_return03_out_13),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[100]),
        .I5(key_in[68]),
        .O(\KR[3].key_reg[0][31] [4]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][4]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[4]),
        .I3(\KR[2].key_reg[1][31] [4]),
        .O(\KR[2].key[1][4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][5]_i_1 
       (.I0(\KR[2].key[1][5]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(p_93_in_16),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[101]),
        .I5(key_in[69]),
        .O(\KR[3].key_reg[0][31] [5]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][5]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[5]),
        .I3(\KR[2].key_reg[1][31] [5]),
        .O(\KR[2].key[1][5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][6]_i_1 
       (.I0(\KR[2].key[1][6]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(isomorphism_inv_return033_out_12),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[102]),
        .I5(key_in[70]),
        .O(\KR[3].key_reg[0][31] [6]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][6]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[6]),
        .I3(\KR[2].key_reg[1][31] [6]),
        .O(\KR[2].key[1][6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][7]_i_1 
       (.I0(\KR[2].key[1][7]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(isomorphism_inv_return05_out_14),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[103]),
        .I5(key_in[71]),
        .O(\KR[3].key_reg[0][31] [7]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][7]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[7]),
        .I3(\KR[2].key_reg[1][31] [7]),
        .O(\KR[2].key[1][7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][8]_i_1 
       (.I0(\KR[2].key[1][8]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(p_86_in_9),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[104]),
        .I5(key_in[72]),
        .O(\KR[3].key_reg[0][31] [8]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][8]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[8]),
        .I3(\KR[2].key_reg[1][31] [8]),
        .O(\KR[2].key[1][8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAEAEEEAEEAEAA)) 
    \KR[2].key[1][9]_i_1 
       (.I0(\KR[2].key[1][9]_i_2_n_0 ),
        .I1(key_sel_mux),
        .I2(p_16_in_11),
        .I3(\AES_CORE_DATAPATH/key1_mux_cnt ),
        .I4(key_in[105]),
        .I5(key_in[73]),
        .O(\KR[3].key_reg[0][31] [9]));
  LUT4 #(
    .INIT(16'h5140)) 
    \KR[2].key[1][9]_i_2 
       (.I0(key_sel_mux),
        .I1(key_en[1]),
        .I2(enable_i[9]),
        .I3(\KR[2].key_reg[1][31] [9]),
        .O(\KR[2].key[1][9]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF2E22FFFF)) 
    \KR[3].key[0][31]_i_1 
       (.I0(\KR[0].key_reg[3][31] [0]),
        .I1(bypass_key_en),
        .I2(\FSM_sequential_state_reg[3]_2 ),
        .I3(\KR[3].key[0][31]_i_4_n_0 ),
        .I4(\KR[3].key_reg[0][31]_0 ),
        .I5(key_en[0]),
        .O(\key_en_pp1_reg[0] ));
  LUT2 #(
    .INIT(4'hB)) 
    \KR[3].key[0][31]_i_3 
       (.I0(Q[3]),
        .I1(Q[2]),
        .O(\FSM_sequential_state_reg[3]_2 ));
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \KR[3].key[0][31]_i_4 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(\KR[3].key[0][31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[3]_i_3 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [3]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [3]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [3]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][3] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[3]_i_3__0 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [11]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [11]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [11]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][11] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[3]_i_3__1 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [27]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [27]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [27]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][27] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[3]_i_3__2 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [19]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [19]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [19]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][19] ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[3]_i_4 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[59]),
        .I5(key_in[27]),
        .O(\AES_CORE_DATAPATH/g_in [3]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[3]_i_4__0 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[35]),
        .I5(key_in[3]),
        .O(\AES_CORE_DATAPATH/g_in [11]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[3]_i_4__1 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[51]),
        .I5(key_in[19]),
        .O(\AES_CORE_DATAPATH/g_in [27]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[3]_i_4__2 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[43]),
        .I5(key_in[11]),
        .O(\AES_CORE_DATAPATH/g_in [19]));
  LUT6 #(
    .INIT(64'hEEE1EEE1EEE1111E)) 
    \base_new_pp[7]_i_2 
       (.I0(\CD[3].col_reg[0][22] ),
        .I1(\base_new_pp_reg[7]_2 ),
        .I2(\CD[3].col_reg[0][16] ),
        .I3(\base_new_pp_reg[7]_3 ),
        .I4(\base_new_pp_reg[7]_4 ),
        .I5(\CD[3].col_reg[0][17] ),
        .O(isomorphism_return179_out_0));
  LUT6 #(
    .INIT(64'hEEE1EEE1EEE1111E)) 
    \base_new_pp[7]_i_2__0 
       (.I0(\CD[3].col_reg[0][14] ),
        .I1(\base_new_pp_reg[7]_5 ),
        .I2(\CD[3].col_reg[0][8] ),
        .I3(\base_new_pp_reg[7]_6 ),
        .I4(\base_new_pp_reg[7]_7 ),
        .I5(\CD[3].col_reg[0][9] ),
        .O(isomorphism_return179_out_2));
  LUT6 #(
    .INIT(64'hEEE1EEE1EEE1111E)) 
    \base_new_pp[7]_i_2__1 
       (.I0(\CD[3].col_reg[0][6] ),
        .I1(\base_new_pp_reg[7]_8 ),
        .I2(\CD[3].col_reg[0][0] ),
        .I3(\base_new_pp_reg[7]_9 ),
        .I4(\base_new_pp_reg[7]_10 ),
        .I5(\CD[3].col_reg[0][1] ),
        .O(isomorphism_return179_out_4));
  LUT6 #(
    .INIT(64'hFF77FF7F77777777)) 
    \base_new_pp[7]_i_2__2 
       (.I0(\key_en_pp1_reg[3]_0 ),
        .I1(\info_o[0]_0 [1]),
        .I2(Q[0]),
        .I3(Q[1]),
        .I4(Q[3]),
        .I5(Q[2]),
        .O(enc_dec_sbox));
  LUT6 #(
    .INIT(64'hEEE1EEE1EEE1111E)) 
    \base_new_pp[7]_i_3 
       (.I0(\CD[3].col_reg[0][30] ),
        .I1(\base_new_pp_reg[7] ),
        .I2(\CD[3].col_reg[0][24] ),
        .I3(\base_new_pp_reg[7]_0 ),
        .I4(\base_new_pp_reg[7]_1 ),
        .I5(\CD[3].col_reg[0][25] ),
        .O(isomorphism_return179_out));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[7]_i_3__0 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [6]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [6]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [6]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][6] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[7]_i_3__1 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [14]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [14]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [14]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][14] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[7]_i_3__2 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [22]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [22]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [22]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][22] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[7]_i_4 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [0]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [0]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [0]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][0] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[7]_i_4__0 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [30]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [30]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [30]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][30] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[7]_i_4__1 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [8]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [8]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [8]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][8] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[7]_i_4__2 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [16]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [16]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [16]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][16] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[7]_i_5 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [1]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [1]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [1]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][1] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[7]_i_5__0 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [9]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [9]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [9]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][9] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[7]_i_5__1 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [24]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [24]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [24]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][24] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[7]_i_5__2 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [17]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [17]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [17]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][17] ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[7]_i_6 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[62]),
        .I5(key_in[30]),
        .O(\AES_CORE_DATAPATH/g_in [6]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[7]_i_6__0 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[38]),
        .I5(key_in[6]),
        .O(\AES_CORE_DATAPATH/g_in [14]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[7]_i_6__1 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[46]),
        .I5(key_in[14]),
        .O(\AES_CORE_DATAPATH/g_in [22]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \base_new_pp[7]_i_6__2 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [25]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [25]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [25]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][25] ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[7]_i_7 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[56]),
        .I5(key_in[24]),
        .O(\AES_CORE_DATAPATH/g_in [0]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[7]_i_7__0 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[54]),
        .I5(key_in[22]),
        .O(\AES_CORE_DATAPATH/g_in [30]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[7]_i_7__1 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[32]),
        .I5(key_in[0]),
        .O(\AES_CORE_DATAPATH/g_in [8]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[7]_i_7__2 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[40]),
        .I5(key_in[8]),
        .O(\AES_CORE_DATAPATH/g_in [16]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[7]_i_8 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[57]),
        .I5(key_in[25]),
        .O(\AES_CORE_DATAPATH/g_in [1]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[7]_i_8__0 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[33]),
        .I5(key_in[1]),
        .O(\AES_CORE_DATAPATH/g_in [9]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[7]_i_8__1 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[48]),
        .I5(key_in[16]),
        .O(\AES_CORE_DATAPATH/g_in [24]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[7]_i_8__2 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[41]),
        .I5(key_in[9]),
        .O(\AES_CORE_DATAPATH/g_in [17]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \base_new_pp[7]_i_9 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[49]),
        .I5(key_in[17]),
        .O(\AES_CORE_DATAPATH/g_in [25]));
  LUT6 #(
    .INIT(64'hFFFF040404FF0404)) 
    ccf_i_1
       (.I0(Q[2]),
        .I1(Q[3]),
        .I2(\FSM_sequential_state_reg[0]_0 ),
        .I3(enable_i[7]),
        .I4(ccf),
        .I5(ccf_reg_0),
        .O(\FSM_sequential_state_reg[2]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT2 #(
    .INIT(4'hE)) 
    ccf_i_2
       (.I0(Q[0]),
        .I1(Q[1]),
        .O(\FSM_sequential_state_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0F0300800F000000)) 
    \col_en_cnt_unit_pp1[0]_i_1 
       (.I0(\rd_count_reg[3]_0 ),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(Q[1]),
        .I4(Q[0]),
        .I5(\col_en_cnt_unit_pp1_reg[3] ),
        .O(\FSM_sequential_state_reg[2]_2 [0]));
  LUT6 #(
    .INIT(64'h04050F0A000F8000)) 
    \col_en_cnt_unit_pp1[1]_i_1 
       (.I0(\col_en_cnt_unit_pp1_reg[3] ),
        .I1(\rd_count_reg[3]_0 ),
        .I2(Q[2]),
        .I3(Q[3]),
        .I4(Q[1]),
        .I5(Q[0]),
        .O(\FSM_sequential_state_reg[2]_2 [1]));
  LUT6 #(
    .INIT(64'h1102308301023003)) 
    \col_en_cnt_unit_pp1[2]_i_1 
       (.I0(\col_en_cnt_unit_pp1_reg[3] ),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[1]),
        .I4(Q[0]),
        .I5(\rd_count_reg[3]_0 ),
        .O(\FSM_sequential_state_reg[2]_2 [2]));
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \col_en_cnt_unit_pp1[3]_i_1 
       (.I0(Q[3]),
        .I1(Q[2]),
        .O(\FSM_sequential_state_reg[3]_6 ));
  LUT6 #(
    .INIT(64'h1100010003C003C0)) 
    \col_en_cnt_unit_pp1[3]_i_2 
       (.I0(\col_en_cnt_unit_pp1_reg[3] ),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(\rd_count_reg[3]_0 ),
        .I5(Q[1]),
        .O(\FSM_sequential_state_reg[2]_2 [3]));
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \col_en_cnt_unit_pp1[3]_i_4 
       (.I0(\rd_count_reg[3]_1 [3]),
        .I1(\rd_count_reg[3]_1 [2]),
        .I2(\rd_count_reg[3]_1 [1]),
        .O(\rd_count_reg[3]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT5 #(
    .INIT(32'hEEEEEEEF)) 
    \col_sel_pp1[0]_i_1 
       (.I0(\col_sel_pp1[0]_i_2_n_0 ),
        .I1(\col_sel_pp1[0]_i_3_n_0 ),
        .I2(Q[3]),
        .I3(Q[2]),
        .I4(Q[0]),
        .O(D[0]));
  LUT6 #(
    .INIT(64'h2231334102010201)) 
    \col_sel_pp1[0]_i_2 
       (.I0(\col_en_cnt_unit_pp1_reg[3] ),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(Q[1]),
        .I4(Q[0]),
        .I5(\rd_count_reg[3]_0 ),
        .O(\col_sel_pp1[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h080808080202FF02)) 
    \col_sel_pp1[0]_i_3 
       (.I0(\col_sel_pp1[0]_i_4_n_0 ),
        .I1(\info_o[0]_0 [2]),
        .I2(\rd_count_reg[3]_0 ),
        .I3(\col_sel_pp1[0]_i_5_n_0 ),
        .I4(\info_o[0]_0 [1]),
        .I5(\info_o[0]_0 [3]),
        .O(\col_sel_pp1[0]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT4 #(
    .INIT(16'h4448)) 
    \col_sel_pp1[0]_i_4 
       (.I0(Q[2]),
        .I1(Q[3]),
        .I2(Q[0]),
        .I3(Q[1]),
        .O(\col_sel_pp1[0]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT5 #(
    .INIT(32'h0F1C0C0C)) 
    \col_sel_pp1[0]_i_5 
       (.I0(\rd_count_reg[3]_0 ),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(Q[0]),
        .I4(Q[3]),
        .O(\col_sel_pp1[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFF4FFFF444F0000)) 
    \col_sel_pp1[1]_i_1 
       (.I0(\rd_count_reg[3]_0 ),
        .I1(\col_sel_pp1_reg[1] ),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[3]),
        .I5(Q[2]),
        .O(D[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8880000)) 
    \info_o[0]_INST_0 
       (.I0(\info_o[31] ),
        .I1(iv_out[0]),
        .I2(key_out[0]),
        .I3(\info_o[31]_0 ),
        .I4(\aes_cr_reg[7] ),
        .I5(info_o_0_sn_1),
        .O(info_o[0]));
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[0]_INST_0_i_1 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [0]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(\info_o[31]_3 [0]),
        .I4(\info_o[0]_INST_0_i_5_n_0 ),
        .O(iv_out[0]));
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT5 #(
    .INIT(32'h00000200)) 
    \info_o[0]_INST_0_i_3 
       (.I0(\info_o[0]_0 [4]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(Q[3]),
        .I4(Q[2]),
        .O(\aes_cr_reg[7] ));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[0]_INST_0_i_5 
       (.I0(\CD[0].col[3][31]_i_13_0 [0]),
        .I1(\CD[0].col[3][31]_i_13_1 [0]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[0]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[10]_INST_0 
       (.I0(iv_out[10]),
        .I1(\info_o[31] ),
        .I2(ccf_reg),
        .I3(col_out[5]),
        .I4(info_o_10_sn_1),
        .O(info_o[6]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[10]_INST_0_i_1 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [10]),
        .I2(\info_o[31]_3 [6]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[10]_INST_0_i_4_n_0 ),
        .O(iv_out[10]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[10]_INST_0_i_4 
       (.I0(\CD[0].col[3][31]_i_13_0 [10]),
        .I1(\CD[0].col[3][31]_i_13_1 [10]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[10]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[11]_INST_0 
       (.I0(iv_out[11]),
        .I1(\info_o[31] ),
        .I2(ccf_reg),
        .I3(col_out[6]),
        .I4(info_o_11_sn_1),
        .O(info_o[7]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[11]_INST_0_i_1 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [11]),
        .I2(\info_o[31]_3 [7]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[11]_INST_0_i_4_n_0 ),
        .O(iv_out[11]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[11]_INST_0_i_4 
       (.I0(\CD[0].col[3][31]_i_13_0 [11]),
        .I1(\CD[0].col[3][31]_i_13_1 [11]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[11]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[12]_INST_0 
       (.I0(iv_out[12]),
        .I1(\info_o[31] ),
        .I2(ccf_reg),
        .I3(col_out[7]),
        .I4(info_o_12_sn_1),
        .O(info_o[8]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[12]_INST_0_i_1 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [12]),
        .I2(\info_o[31]_3 [8]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[12]_INST_0_i_4_n_0 ),
        .O(iv_out[12]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[12]_INST_0_i_4 
       (.I0(\CD[0].col[3][31]_i_13_0 [12]),
        .I1(\CD[0].col[3][31]_i_13_1 [12]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[12]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[13]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[8]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[3]),
        .I4(iv_out[13]),
        .I5(\info_o[31] ),
        .O(info_o[9]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[13]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [13]),
        .I2(\info_o[31]_3 [9]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[13]_INST_0_i_4_n_0 ),
        .O(iv_out[13]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[13]_INST_0_i_4 
       (.I0(\CD[0].col[3][31]_i_13_0 [13]),
        .I1(\CD[0].col[3][31]_i_13_1 [13]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[13]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[14]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[9]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[4]),
        .I4(iv_out[14]),
        .I5(\info_o[31] ),
        .O(info_o[10]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[14]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [14]),
        .I2(\info_o[31]_3 [10]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[14]_INST_0_i_4_n_0 ),
        .O(iv_out[14]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[14]_INST_0_i_4 
       (.I0(\CD[0].col[3][31]_i_13_0 [14]),
        .I1(\CD[0].col[3][31]_i_13_1 [14]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[14]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[15]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[10]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[5]),
        .I4(iv_out[15]),
        .I5(\info_o[31] ),
        .O(info_o[11]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[15]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [15]),
        .I2(\info_o[31]_3 [11]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[15]_INST_0_i_4_n_0 ),
        .O(iv_out[15]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[15]_INST_0_i_4 
       (.I0(\CD[0].col[3][31]_i_13_0 [15]),
        .I1(\CD[0].col[3][31]_i_13_1 [15]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[15]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[16]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[11]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[6]),
        .I4(iv_out[16]),
        .I5(\info_o[31] ),
        .O(info_o[12]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[16]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [16]),
        .I2(\info_o[31]_3 [12]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[16]_INST_0_i_5_n_0 ),
        .O(iv_out[16]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[16]_INST_0_i_5 
       (.I0(\CD[0].col[3][31]_i_13_0 [16]),
        .I1(\CD[0].col[3][31]_i_13_1 [16]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[16]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[17]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[12]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[7]),
        .I4(iv_out[17]),
        .I5(\info_o[31] ),
        .O(info_o[13]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[17]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [17]),
        .I2(\info_o[31]_3 [13]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[17]_INST_0_i_5_n_0 ),
        .O(iv_out[17]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[17]_INST_0_i_5 
       (.I0(\CD[0].col[3][31]_i_13_0 [17]),
        .I1(\CD[0].col[3][31]_i_13_1 [17]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[17]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[18]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[13]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[8]),
        .I4(iv_out[18]),
        .I5(\info_o[31] ),
        .O(info_o[14]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[18]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [18]),
        .I2(\info_o[31]_3 [14]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[18]_INST_0_i_5_n_0 ),
        .O(iv_out[18]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[18]_INST_0_i_5 
       (.I0(\CD[0].col[3][31]_i_13_0 [18]),
        .I1(\CD[0].col[3][31]_i_13_1 [18]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[18]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[19]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[14]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[9]),
        .I4(iv_out[19]),
        .I5(\info_o[31] ),
        .O(info_o[15]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[19]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [19]),
        .I2(\info_o[31]_3 [15]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[19]_INST_0_i_5_n_0 ),
        .O(iv_out[19]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[19]_INST_0_i_5 
       (.I0(\CD[0].col[3][31]_i_13_0 [19]),
        .I1(\CD[0].col[3][31]_i_13_1 [19]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[19]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[20]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[15]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[10]),
        .I4(iv_out[20]),
        .I5(\info_o[31] ),
        .O(info_o[16]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[20]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [20]),
        .I2(\info_o[31]_3 [16]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[20]_INST_0_i_5_n_0 ),
        .O(iv_out[20]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[20]_INST_0_i_5 
       (.I0(\CD[0].col[3][31]_i_13_0 [20]),
        .I1(\CD[0].col[3][31]_i_13_1 [20]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[20]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[21]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[16]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[11]),
        .I4(iv_out[21]),
        .I5(\info_o[31] ),
        .O(info_o[17]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[21]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [21]),
        .I2(\info_o[31]_3 [17]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[21]_INST_0_i_5_n_0 ),
        .O(iv_out[21]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[21]_INST_0_i_5 
       (.I0(\CD[0].col[3][31]_i_13_0 [21]),
        .I1(\CD[0].col[3][31]_i_13_1 [21]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[21]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[22]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[17]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[12]),
        .I4(iv_out[22]),
        .I5(\info_o[31] ),
        .O(info_o[18]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[22]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [22]),
        .I2(\info_o[31]_3 [18]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[22]_INST_0_i_5_n_0 ),
        .O(iv_out[22]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[22]_INST_0_i_5 
       (.I0(\CD[0].col[3][31]_i_13_0 [22]),
        .I1(\CD[0].col[3][31]_i_13_1 [22]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[22]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[23]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[18]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[13]),
        .I4(iv_out[23]),
        .I5(\info_o[31] ),
        .O(info_o[19]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[23]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [23]),
        .I2(\info_o[31]_3 [19]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[23]_INST_0_i_5_n_0 ),
        .O(iv_out[23]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[23]_INST_0_i_5 
       (.I0(\CD[0].col[3][31]_i_13_0 [23]),
        .I1(\CD[0].col[3][31]_i_13_1 [23]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[23]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[24]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[19]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[14]),
        .I4(iv_out[24]),
        .I5(\info_o[31] ),
        .O(info_o[20]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[24]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [24]),
        .I2(\info_o[31]_3 [20]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[24]_INST_0_i_6_n_0 ),
        .O(iv_out[24]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[24]_INST_0_i_6 
       (.I0(\CD[0].col[3][31]_i_13_0 [24]),
        .I1(\CD[0].col[3][31]_i_13_1 [24]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[24]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[25]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[20]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[15]),
        .I4(iv_out[25]),
        .I5(\info_o[31] ),
        .O(info_o[21]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[25]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [25]),
        .I2(\info_o[31]_3 [21]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[25]_INST_0_i_6_n_0 ),
        .O(iv_out[25]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[25]_INST_0_i_6 
       (.I0(\CD[0].col[3][31]_i_13_0 [25]),
        .I1(\CD[0].col[3][31]_i_13_1 [25]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[25]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[26]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[21]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[16]),
        .I4(iv_out[26]),
        .I5(\info_o[31] ),
        .O(info_o[22]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[26]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [26]),
        .I2(\info_o[31]_3 [22]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[26]_INST_0_i_6_n_0 ),
        .O(iv_out[26]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[26]_INST_0_i_6 
       (.I0(\CD[0].col[3][31]_i_13_0 [26]),
        .I1(\CD[0].col[3][31]_i_13_1 [26]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[26]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[27]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[22]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[17]),
        .I4(iv_out[27]),
        .I5(\info_o[31] ),
        .O(info_o[23]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[27]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [27]),
        .I2(\info_o[31]_3 [23]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[27]_INST_0_i_6_n_0 ),
        .O(iv_out[27]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[27]_INST_0_i_6 
       (.I0(\CD[0].col[3][31]_i_13_0 [27]),
        .I1(\CD[0].col[3][31]_i_13_1 [27]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[27]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[28]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[23]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[18]),
        .I4(iv_out[28]),
        .I5(\info_o[31] ),
        .O(info_o[24]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[28]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [28]),
        .I2(\info_o[31]_3 [24]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[28]_INST_0_i_8_n_0 ),
        .O(iv_out[28]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[28]_INST_0_i_8 
       (.I0(\CD[0].col[3][31]_i_13_0 [28]),
        .I1(\CD[0].col[3][31]_i_13_1 [28]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[28]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[29]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[24]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[19]),
        .I4(iv_out[29]),
        .I5(\info_o[31] ),
        .O(info_o[25]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[29]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [29]),
        .I2(\info_o[31]_3 [25]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[29]_INST_0_i_8_n_0 ),
        .O(iv_out[29]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[29]_INST_0_i_8 
       (.I0(\CD[0].col[3][31]_i_13_0 [29]),
        .I1(\CD[0].col[3][31]_i_13_1 [29]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[29]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[30]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[25]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[20]),
        .I4(iv_out[30]),
        .I5(\info_o[31] ),
        .O(info_o[26]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[30]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [30]),
        .I2(\info_o[31]_3 [26]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[30]_INST_0_i_8_n_0 ),
        .O(iv_out[30]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[30]_INST_0_i_8 
       (.I0(\CD[0].col[3][31]_i_13_0 [30]),
        .I1(\CD[0].col[3][31]_i_13_1 [30]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[30]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[31]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[26]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[21]),
        .I4(iv_out[31]),
        .I5(\info_o[31] ),
        .O(info_o[27]));
  LUT6 #(
    .INIT(64'h00000000AAAAABAA)) 
    \info_o[31]_INST_0_i_1 
       (.I0(ccf),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(Q[3]),
        .I4(Q[2]),
        .I5(\info_o[31]_1 ),
        .O(ccf_reg));
  LUT5 #(
    .INIT(32'hFFFF5404)) 
    \info_o[31]_INST_0_i_12 
       (.I0(bypass_key_en),
        .I1(\info_o[31]_INST_0_i_4 ),
        .I2(\info_o[31]_INST_0_i_4_0 ),
        .I3(\info_o[31]_INST_0_i_4_1 ),
        .I4(\info_o[31]_INST_0_i_26_n_0 ),
        .O(\key_out_sel_pp1_reg[1] ));
  LUT2 #(
    .INIT(4'h2)) 
    \info_o[31]_INST_0_i_14 
       (.I0(iv_mux_out13_out),
        .I1(\col_en_cnt_unit_pp2_reg[3] ),
        .O(\info_o[31]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB8FFB8)) 
    \info_o[31]_INST_0_i_15 
       (.I0(\FSM_sequential_state_reg[2]_2 [3]),
        .I1(\FSM_sequential_state_reg[2]_5 ),
        .I2(\CD[0].col_reg[3][31]_1 [3]),
        .I3(col_en_host[3]),
        .I4(enable_i[0]),
        .I5(\CD[0].col[3][31]_i_22 ),
        .O(\col_en_cnt_unit_pp2_reg[3] ));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[31]_INST_0_i_16 
       (.I0(\CD[0].col[3][31]_i_13_0 [31]),
        .I1(\CD[0].col[3][31]_i_13_1 [31]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[31]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0A0A0E0E00000E00)) 
    \info_o[31]_INST_0_i_17 
       (.I0(\FSM_sequential_state_reg[2]_3 [0]),
        .I1(\info_o[28]_INST_0_i_15 ),
        .I2(sbox_sel),
        .I3(\info_o[28]_INST_0_i_15_0 ),
        .I4(\info_o[31]_1 ),
        .I5(\FSM_sequential_state_reg[2]_3 [1]),
        .O(\FSM_sequential_state_reg[3]_4 ));
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT5 #(
    .INIT(32'hFF010101)) 
    \info_o[31]_INST_0_i_26 
       (.I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(enable_i[2]),
        .I4(\info_o[31]_INST_0_i_12_0 ),
        .O(\info_o[31]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \info_o[31]_INST_0_i_28 
       (.I0(\FSM_sequential_state_reg[2]_2 [2]),
        .I1(\FSM_sequential_state_reg[2]_5 ),
        .I2(\CD[0].col_reg[3][31]_1 [2]),
        .I3(col_en_host[2]),
        .I4(enable_i[0]),
        .I5(\CD[0].col[3][31]_i_22 ),
        .O(iv_mux_out13_out));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB8FFB8)) 
    \info_o[31]_INST_0_i_30 
       (.I0(\FSM_sequential_state_reg[2]_2 [1]),
        .I1(\FSM_sequential_state_reg[2]_5 ),
        .I2(\CD[0].col_reg[3][31]_1 [1]),
        .I3(col_en_host[1]),
        .I4(enable_i[0]),
        .I5(\CD[0].col[3][10]_i_12_0 ),
        .O(\AES_CORE_DATAPATH/iv_mux_out10_out ));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \info_o[31]_INST_0_i_31 
       (.I0(\FSM_sequential_state_reg[2]_2 [0]),
        .I1(\FSM_sequential_state_reg[2]_5 ),
        .I2(\CD[0].col_reg[3][31]_1 [0]),
        .I3(col_en_host[0]),
        .I4(enable_i[0]),
        .I5(\CD[0].col[3][10]_i_12_0 ),
        .O(\AES_CORE_DATAPATH/iv_mux_out1 ));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \info_o[31]_INST_0_i_33 
       (.I0(Q[2]),
        .I1(Q[3]),
        .I2(Q[0]),
        .O(sbox_sel));
  LUT6 #(
    .INIT(64'h0000000005050001)) 
    \info_o[31]_INST_0_i_35 
       (.I0(\FSM_sequential_state_reg[2]_3 [0]),
        .I1(\info_o[28]_INST_0_i_15 ),
        .I2(sbox_sel),
        .I3(\info_o[28]_INST_0_i_15_0 ),
        .I4(\info_o[31]_1 ),
        .I5(\FSM_sequential_state_reg[2]_3 [1]),
        .O(\FSM_sequential_state_reg[3]_3 ));
  LUT6 #(
    .INIT(64'h000000000A0A0002)) 
    \info_o[31]_INST_0_i_36 
       (.I0(sbox_sel),
        .I1(\info_o[28]_INST_0_i_15 ),
        .I2(\FSM_sequential_state_reg[2]_3 [0]),
        .I3(\info_o[28]_INST_0_i_15_0 ),
        .I4(\info_o[31]_1 ),
        .I5(\FSM_sequential_state_reg[2]_3 [1]),
        .O(\FSM_sequential_state_reg[2]_6 ));
  LUT6 #(
    .INIT(64'h000000000A0A000E)) 
    \info_o[31]_INST_0_i_37 
       (.I0(\FSM_sequential_state_reg[2]_3 [0]),
        .I1(\info_o[28]_INST_0_i_15 ),
        .I2(sbox_sel),
        .I3(\info_o[28]_INST_0_i_15_0 ),
        .I4(\info_o[31]_1 ),
        .I5(\FSM_sequential_state_reg[2]_3 [1]),
        .O(\FSM_sequential_state_reg[3]_7 ));
  LUT6 #(
    .INIT(64'h0505010100000100)) 
    \info_o[31]_INST_0_i_38 
       (.I0(\FSM_sequential_state_reg[2]_3 [0]),
        .I1(\info_o[28]_INST_0_i_15 ),
        .I2(sbox_sel),
        .I3(\info_o[28]_INST_0_i_15_0 ),
        .I4(\info_o[31]_1 ),
        .I5(\FSM_sequential_state_reg[2]_3 [1]),
        .O(\FSM_sequential_state_reg[3]_8 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[31]_INST_0_i_5 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [31]),
        .I2(\info_o[31]_3 [27]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[31]_INST_0_i_16_n_0 ),
        .O(iv_out[31]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[4]_INST_0 
       (.I0(iv_out[4]),
        .I1(\info_o[31] ),
        .I2(ccf_reg),
        .I3(col_out[0]),
        .I4(info_o_4_sn_1),
        .O(info_o[1]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[4]_INST_0_i_1 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [4]),
        .I2(\info_o[31]_3 [1]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[4]_INST_0_i_4_n_0 ),
        .O(iv_out[4]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[4]_INST_0_i_4 
       (.I0(\CD[0].col[3][31]_i_13_0 [4]),
        .I1(\CD[0].col[3][31]_i_13_1 [4]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[4]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[6]_INST_0 
       (.I0(iv_out[6]),
        .I1(\info_o[31] ),
        .I2(ccf_reg),
        .I3(col_out[1]),
        .I4(info_o_6_sn_1),
        .O(info_o[2]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[6]_INST_0_i_1 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [6]),
        .I2(\info_o[31]_3 [2]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[6]_INST_0_i_4_n_0 ),
        .O(iv_out[6]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[6]_INST_0_i_4 
       (.I0(\CD[0].col[3][31]_i_13_0 [6]),
        .I1(\CD[0].col[3][31]_i_13_1 [6]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[6]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[7]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[2]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[1]),
        .I4(iv_out[7]),
        .I5(\info_o[31] ),
        .O(info_o[3]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[7]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [7]),
        .I2(\info_o[31]_3 [3]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[7]_INST_0_i_4_n_0 ),
        .O(iv_out[7]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[7]_INST_0_i_4 
       (.I0(\CD[0].col[3][31]_i_13_0 [7]),
        .I1(\CD[0].col[3][31]_i_13_1 [7]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[7]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \info_o[8]_INST_0 
       (.I0(ccf_reg),
        .I1(col_out[3]),
        .I2(\info_o[31]_0 ),
        .I3(key_out[2]),
        .I4(iv_out[8]),
        .I5(\info_o[31] ),
        .O(info_o[4]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[8]_INST_0_i_3 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [8]),
        .I2(\info_o[31]_3 [4]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[8]_INST_0_i_4_n_0 ),
        .O(iv_out[8]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[8]_INST_0_i_4 
       (.I0(\CD[0].col[3][31]_i_13_0 [8]),
        .I1(\CD[0].col[3][31]_i_13_1 [8]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[8]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[9]_INST_0 
       (.I0(iv_out[9]),
        .I1(\info_o[31] ),
        .I2(ccf_reg),
        .I3(col_out[4]),
        .I4(info_o_9_sn_1),
        .O(info_o[5]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \info_o[9]_INST_0_i_1 
       (.I0(\info_o[31]_INST_0_i_14_n_0 ),
        .I1(\info_o[31]_2 [9]),
        .I2(\info_o[31]_3 [5]),
        .I3(\col_en_cnt_unit_pp2_reg[3] ),
        .I4(\info_o[9]_INST_0_i_4_n_0 ),
        .O(iv_out[9]));
  LUT6 #(
    .INIT(64'h000A000C000A0000)) 
    \info_o[9]_INST_0_i_4 
       (.I0(\CD[0].col[3][31]_i_13_0 [9]),
        .I1(\CD[0].col[3][31]_i_13_1 [9]),
        .I2(\col_en_cnt_unit_pp2_reg[3] ),
        .I3(iv_mux_out13_out),
        .I4(\AES_CORE_DATAPATH/iv_mux_out10_out ),
        .I5(\AES_CORE_DATAPATH/iv_mux_out1 ),
        .O(\info_o[9]_INST_0_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT4 #(
    .INIT(16'h0090)) 
    \key_en_pp1[0]_i_1 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(Q[3]),
        .O(\FSM_sequential_state_reg[0]_1 [0]));
  LUT6 #(
    .INIT(64'h2666400010000000)) 
    \key_en_pp1[1]_i_1 
       (.I0(Q[2]),
        .I1(Q[3]),
        .I2(\key_en_pp1_reg[3]_0 ),
        .I3(\info_o[0]_0 [1]),
        .I4(Q[1]),
        .I5(Q[0]),
        .O(\FSM_sequential_state_reg[0]_1 [1]));
  LUT6 #(
    .INIT(64'h8888400004441000)) 
    \key_en_pp1[2]_i_1 
       (.I0(Q[2]),
        .I1(Q[3]),
        .I2(\key_en_pp1_reg[3]_0 ),
        .I3(\info_o[0]_0 [1]),
        .I4(Q[0]),
        .I5(Q[1]),
        .O(\FSM_sequential_state_reg[0]_1 [2]));
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT4 #(
    .INIT(16'h2E6E)) 
    \key_en_pp1[3]_i_1 
       (.I0(Q[3]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(\FSM_sequential_state_reg[3]_5 ));
  LUT6 #(
    .INIT(64'h4050505042000000)) 
    \key_en_pp1[3]_i_2 
       (.I0(Q[0]),
        .I1(Q[2]),
        .I2(Q[3]),
        .I3(\info_o[0]_0 [1]),
        .I4(\key_en_pp1_reg[3]_0 ),
        .I5(Q[1]),
        .O(\FSM_sequential_state_reg[0]_1 [3]));
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT4 #(
    .INIT(16'h0318)) 
    \key_out_sel_pp1[0]_i_1 
       (.I0(Q[3]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(\FSM_sequential_state_reg[2]_3 [0]));
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT4 #(
    .INIT(16'h0149)) 
    \key_out_sel_pp1[1]_i_1 
       (.I0(Q[2]),
        .I1(Q[3]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(\FSM_sequential_state_reg[2]_3 [1]));
  LUT6 #(
    .INIT(64'hFFF000F8F0F8FF08)) 
    key_sel_pp1_i_1
       (.I0(\key_en_pp1_reg[3]_0 ),
        .I1(\info_o[0]_0 [1]),
        .I2(Q[3]),
        .I3(Q[2]),
        .I4(Q[1]),
        .I5(Q[0]),
        .O(key_sel));
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'h20)) 
    last_round_pp1_i_1
       (.I0(\rd_count_reg[3]_1 [1]),
        .I1(\rd_count_reg[3]_1 [2]),
        .I2(\rd_count_reg[3]_1 [3]),
        .O(last_round));
  LUT6 #(
    .INIT(64'h111E111E111EEEE1)) 
    \out_gf_pp[1]_i_5 
       (.I0(\CD[3].col_reg[0][30] ),
        .I1(\base_new_pp_reg[7] ),
        .I2(\CD[3].col_reg[0][24] ),
        .I3(\base_new_pp_reg[7]_0 ),
        .I4(\out_gf_pp[1]_i_2 ),
        .I5(\CD[3].col_reg[0][29] ),
        .O(isomorphism_return114_out));
  LUT6 #(
    .INIT(64'h111E111E111EEEE1)) 
    \out_gf_pp[1]_i_5__0 
       (.I0(\CD[3].col_reg[0][22] ),
        .I1(\base_new_pp_reg[7]_2 ),
        .I2(\CD[3].col_reg[0][16] ),
        .I3(\base_new_pp_reg[7]_3 ),
        .I4(\out_gf_pp[1]_i_2__0 ),
        .I5(\CD[3].col_reg[0][21] ),
        .O(isomorphism_return114_out_1));
  LUT6 #(
    .INIT(64'h111E111E111EEEE1)) 
    \out_gf_pp[1]_i_5__1 
       (.I0(\CD[3].col_reg[0][14] ),
        .I1(\base_new_pp_reg[7]_5 ),
        .I2(\CD[3].col_reg[0][8] ),
        .I3(\base_new_pp_reg[7]_6 ),
        .I4(\out_gf_pp[1]_i_2__1 ),
        .I5(\CD[3].col_reg[0][13] ),
        .O(isomorphism_return114_out_3));
  LUT6 #(
    .INIT(64'h111E111E111EEEE1)) 
    \out_gf_pp[1]_i_5__2 
       (.I0(\CD[3].col_reg[0][6] ),
        .I1(\base_new_pp_reg[7]_8 ),
        .I2(\CD[3].col_reg[0][0] ),
        .I3(\base_new_pp_reg[7]_9 ),
        .I4(\out_gf_pp[1]_i_2__2 ),
        .I5(\CD[3].col_reg[0][5] ),
        .O(isomorphism_return114_out_5));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \out_gf_pp[1]_i_6 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [5]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [5]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [5]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][5] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \out_gf_pp[1]_i_6__0 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [13]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [13]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [13]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][13] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \out_gf_pp[1]_i_6__1 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [29]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [29]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [29]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][29] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \out_gf_pp[1]_i_6__2 
       (.I0(\FSM_sequential_state_reg[2]_6 ),
        .I1(\AES_CORE_DATAPATH/g_in [21]),
        .I2(\FSM_sequential_state_reg[3]_3 ),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 [21]),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [21]),
        .I5(\FSM_sequential_state_reg[3]_4 ),
        .O(\CD[3].col_reg[0][21] ));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \out_gf_pp[1]_i_7 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[61]),
        .I5(key_in[29]),
        .O(\AES_CORE_DATAPATH/g_in [5]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \out_gf_pp[1]_i_7__0 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[37]),
        .I5(key_in[5]),
        .O(\AES_CORE_DATAPATH/g_in [13]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \out_gf_pp[1]_i_7__1 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[53]),
        .I5(key_in[21]),
        .O(\AES_CORE_DATAPATH/g_in [29]));
  LUT6 #(
    .INIT(64'hAAABFFFF55540000)) 
    \out_gf_pp[1]_i_7__2 
       (.I0(enc_dec),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(\FSM_sequential_state_reg[3]_2 ),
        .I4(key_in[45]),
        .I5(key_in[13]),
        .O(\AES_CORE_DATAPATH/g_in [21]));
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT5 #(
    .INIT(32'h33233033)) 
    \rd_count[0]_i_1 
       (.I0(\rd_count_reg[3]_0 ),
        .I1(\rd_count_reg[3]_1 [0]),
        .I2(Q[3]),
        .I3(Q[0]),
        .I4(Q[1]),
        .O(\rd_count[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000F8F8FF000000)) 
    \rd_count[1]_i_1 
       (.I0(Q[1]),
        .I1(\rd_count[1]_i_2_n_0 ),
        .I2(\rd_count[3]_i_4_n_0 ),
        .I3(\rd_count[2]_i_2_n_0 ),
        .I4(\rd_count_reg[3]_1 [0]),
        .I5(\rd_count_reg[3]_1 [1]),
        .O(\rd_count[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \rd_count[1]_i_2 
       (.I0(\rd_count_reg[3]_1 [2]),
        .I1(\rd_count_reg[3]_1 [3]),
        .O(\rd_count[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFF0000000000F4F4)) 
    \rd_count[2]_i_1 
       (.I0(\rd_count_reg[3]_1 [3]),
        .I1(Q[1]),
        .I2(\rd_count[3]_i_4_n_0 ),
        .I3(\rd_count[2]_i_2_n_0 ),
        .I4(\rd_count[2]_i_3_n_0 ),
        .I5(\rd_count_reg[3]_1 [2]),
        .O(\rd_count[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT4 #(
    .INIT(16'hFFDF)) 
    \rd_count[2]_i_2 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(Q[3]),
        .O(\rd_count[2]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rd_count[2]_i_3 
       (.I0(\rd_count_reg[3]_1 [0]),
        .I1(\rd_count_reg[3]_1 [1]),
        .O(\rd_count[2]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00703030)) 
    \rd_count[3]_i_1 
       (.I0(\rd_count_reg[3]_0 ),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(Q[0]),
        .I4(Q[1]),
        .O(\rd_count[3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAEAEAAAAFFAEAAAA)) 
    \rd_count[3]_i_2 
       (.I0(\rd_count[3]_i_3_n_0 ),
        .I1(\rd_count[3]_i_4_n_0 ),
        .I2(\rd_count_reg[3]_1 [2]),
        .I3(\rd_count[3]_i_5_n_0 ),
        .I4(\rd_count_reg[3]_1 [3]),
        .I5(\rd_count_reg[3]_1 [0]),
        .O(\rd_count[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0E00E0E00000E0E0)) 
    \rd_count[3]_i_3 
       (.I0(\rd_count[3]_i_6_n_0 ),
        .I1(\FSM_sequential_state_reg[3]_2 ),
        .I2(\rd_count_reg[3]_1 [3]),
        .I3(\rd_count_reg[3]_1 [2]),
        .I4(\rd_count_reg[3]_1 [1]),
        .I5(\rd_count_reg[3]_1 [0]),
        .O(\rd_count[3]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT4 #(
    .INIT(16'hF7DF)) 
    \rd_count[3]_i_4 
       (.I0(Q[2]),
        .I1(Q[3]),
        .I2(Q[0]),
        .I3(Q[1]),
        .O(\rd_count[3]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT5 #(
    .INIT(32'hAAA2FFFF)) 
    \rd_count[3]_i_5 
       (.I0(\rd_count_reg[3]_1 [2]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(Q[3]),
        .I4(Q[2]),
        .O(\rd_count[3]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \rd_count[3]_i_6 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(\rd_count[3]_i_6_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \rd_count_reg[0] 
       (.C(clk_i),
        .CE(\rd_count[3]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\rd_count[0]_i_1_n_0 ),
        .Q(\rd_count_reg[3]_1 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \rd_count_reg[1] 
       (.C(clk_i),
        .CE(\rd_count[3]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\rd_count[1]_i_1_n_0 ),
        .Q(\rd_count_reg[3]_1 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \rd_count_reg[2] 
       (.C(clk_i),
        .CE(\rd_count[3]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\rd_count[2]_i_1_n_0 ),
        .Q(\rd_count_reg[3]_1 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \rd_count_reg[3] 
       (.C(clk_i),
        .CE(\rd_count[3]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\rd_count[3]_i_2_n_0 ),
        .Q(\rd_count_reg[3]_1 [3]));
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT5 #(
    .INIT(32'h000010E0)) 
    \rk_sel_pp1[0]_i_1 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(Q[3]),
        .I3(Q[2]),
        .I4(\rd_count_reg[3]_0 ),
        .O(\FSM_sequential_state_reg[1]_0 [0]));
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT5 #(
    .INIT(32'h10E00000)) 
    \rk_sel_pp1[1]_i_1 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(Q[3]),
        .I3(Q[2]),
        .I4(\rd_count_reg[3]_0 ),
        .O(\FSM_sequential_state_reg[1]_0 [1]));
endmodule

(* ORIG_REF_NAME = "data_swap" *) 
module switch_elements_data_swap
   (bus_swap,
    enable_i,
    \IV_BKP_REGISTERS[3].bkp[3][31]_i_2 );
  output [31:0]bus_swap;
  input [31:0]enable_i;
  input [1:0]\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 ;

  wire [1:0]\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 ;
  wire [31:0]bus_swap;
  wire [31:0]enable_i;

  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][0]_i_4 
       (.I0(enable_i[16]),
        .I1(enable_i[0]),
        .I2(enable_i[31]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[24]),
        .O(bus_swap[0]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][10]_i_7 
       (.I0(enable_i[26]),
        .I1(enable_i[10]),
        .I2(enable_i[21]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[18]),
        .O(bus_swap[10]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][11]_i_7 
       (.I0(enable_i[27]),
        .I1(enable_i[11]),
        .I2(enable_i[20]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[19]),
        .O(bus_swap[11]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][12]_i_7 
       (.I0(enable_i[28]),
        .I1(enable_i[12]),
        .I2(enable_i[19]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[20]),
        .O(bus_swap[12]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][13]_i_7 
       (.I0(enable_i[29]),
        .I1(enable_i[13]),
        .I2(enable_i[18]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[21]),
        .O(bus_swap[13]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][14]_i_7 
       (.I0(enable_i[30]),
        .I1(enable_i[14]),
        .I2(enable_i[17]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[22]),
        .O(bus_swap[14]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][15]_i_10 
       (.I0(enable_i[31]),
        .I1(enable_i[15]),
        .I2(enable_i[16]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[23]),
        .O(bus_swap[15]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][16]_i_5 
       (.I0(enable_i[0]),
        .I1(enable_i[16]),
        .I2(enable_i[15]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[8]),
        .O(bus_swap[16]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][17]_i_5 
       (.I0(enable_i[1]),
        .I1(enable_i[17]),
        .I2(enable_i[14]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[9]),
        .O(bus_swap[17]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][18]_i_5 
       (.I0(enable_i[2]),
        .I1(enable_i[18]),
        .I2(enable_i[13]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[10]),
        .O(bus_swap[18]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][19]_i_5 
       (.I0(enable_i[3]),
        .I1(enable_i[19]),
        .I2(enable_i[12]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[11]),
        .O(bus_swap[19]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][1]_i_4 
       (.I0(enable_i[17]),
        .I1(enable_i[1]),
        .I2(enable_i[30]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[25]),
        .O(bus_swap[1]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][20]_i_5 
       (.I0(enable_i[4]),
        .I1(enable_i[20]),
        .I2(enable_i[11]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[12]),
        .O(bus_swap[20]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][21]_i_5 
       (.I0(enable_i[5]),
        .I1(enable_i[21]),
        .I2(enable_i[10]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[13]),
        .O(bus_swap[21]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][22]_i_5 
       (.I0(enable_i[6]),
        .I1(enable_i[22]),
        .I2(enable_i[9]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[14]),
        .O(bus_swap[22]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][23]_i_5 
       (.I0(enable_i[7]),
        .I1(enable_i[23]),
        .I2(enable_i[8]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[15]),
        .O(bus_swap[23]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][24]_i_4 
       (.I0(enable_i[8]),
        .I1(enable_i[24]),
        .I2(enable_i[7]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[0]),
        .O(bus_swap[24]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][25]_i_4 
       (.I0(enable_i[9]),
        .I1(enable_i[25]),
        .I2(enable_i[6]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[1]),
        .O(bus_swap[25]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][26]_i_4 
       (.I0(enable_i[10]),
        .I1(enable_i[26]),
        .I2(enable_i[5]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[2]),
        .O(bus_swap[26]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][27]_i_4 
       (.I0(enable_i[11]),
        .I1(enable_i[27]),
        .I2(enable_i[4]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[3]),
        .O(bus_swap[27]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][28]_i_4 
       (.I0(enable_i[12]),
        .I1(enable_i[28]),
        .I2(enable_i[3]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[4]),
        .O(bus_swap[28]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][29]_i_4 
       (.I0(enable_i[13]),
        .I1(enable_i[29]),
        .I2(enable_i[2]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[5]),
        .O(bus_swap[29]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][2]_i_4 
       (.I0(enable_i[18]),
        .I1(enable_i[2]),
        .I2(enable_i[29]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[26]),
        .O(bus_swap[2]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][30]_i_4 
       (.I0(enable_i[14]),
        .I1(enable_i[30]),
        .I2(enable_i[1]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[6]),
        .O(bus_swap[30]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][31]_i_5 
       (.I0(enable_i[15]),
        .I1(enable_i[31]),
        .I2(enable_i[0]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[7]),
        .O(bus_swap[31]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][3]_i_4 
       (.I0(enable_i[19]),
        .I1(enable_i[3]),
        .I2(enable_i[28]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[27]),
        .O(bus_swap[3]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][4]_i_4 
       (.I0(enable_i[20]),
        .I1(enable_i[4]),
        .I2(enable_i[27]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[28]),
        .O(bus_swap[4]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][5]_i_4 
       (.I0(enable_i[21]),
        .I1(enable_i[5]),
        .I2(enable_i[26]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[29]),
        .O(bus_swap[5]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][6]_i_4 
       (.I0(enable_i[22]),
        .I1(enable_i[6]),
        .I2(enable_i[25]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[30]),
        .O(bus_swap[6]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][7]_i_4 
       (.I0(enable_i[23]),
        .I1(enable_i[7]),
        .I2(enable_i[24]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[31]),
        .O(bus_swap[7]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][8]_i_7 
       (.I0(enable_i[24]),
        .I1(enable_i[8]),
        .I2(enable_i[23]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[16]),
        .O(bus_swap[8]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \IV_BKP_REGISTERS[3].bkp[3][9]_i_7 
       (.I0(enable_i[25]),
        .I1(enable_i[9]),
        .I2(enable_i[22]),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 [0]),
        .I5(enable_i[17]),
        .O(bus_swap[9]));
endmodule

(* ORIG_REF_NAME = "data_swap" *) 
module switch_elements_data_swap_0
   (col_out,
    \aes_cr_reg[2] ,
    \aes_cr_reg[2]_0 ,
    sbox_input,
    \info_o[1] );
  output [0:0]col_out;
  output [2:0]\aes_cr_reg[2] ;
  output [26:0]\aes_cr_reg[2]_0 ;
  input [31:0]sbox_input;
  input [1:0]\info_o[1] ;

  wire [2:0]\aes_cr_reg[2] ;
  wire [26:0]\aes_cr_reg[2]_0 ;
  wire [0:0]col_out;
  wire [1:0]\info_o[1] ;
  wire [31:0]sbox_input;

  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[0]_INST_0_i_6 
       (.I0(sbox_input[16]),
        .I1(sbox_input[0]),
        .I2(sbox_input[31]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[24]),
        .O(col_out));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[10]_INST_0_i_2 
       (.I0(sbox_input[26]),
        .I1(sbox_input[10]),
        .I2(sbox_input[21]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[18]),
        .O(\aes_cr_reg[2]_0 [5]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[11]_INST_0_i_2 
       (.I0(sbox_input[27]),
        .I1(sbox_input[11]),
        .I2(sbox_input[20]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[19]),
        .O(\aes_cr_reg[2]_0 [6]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[12]_INST_0_i_2 
       (.I0(sbox_input[28]),
        .I1(sbox_input[12]),
        .I2(sbox_input[19]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[20]),
        .O(\aes_cr_reg[2]_0 [7]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[13]_INST_0_i_1 
       (.I0(sbox_input[29]),
        .I1(sbox_input[13]),
        .I2(sbox_input[18]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[21]),
        .O(\aes_cr_reg[2]_0 [8]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[14]_INST_0_i_1 
       (.I0(sbox_input[30]),
        .I1(sbox_input[14]),
        .I2(sbox_input[17]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[22]),
        .O(\aes_cr_reg[2]_0 [9]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[15]_INST_0_i_1 
       (.I0(sbox_input[31]),
        .I1(sbox_input[15]),
        .I2(sbox_input[16]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[23]),
        .O(\aes_cr_reg[2]_0 [10]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[16]_INST_0_i_1 
       (.I0(sbox_input[0]),
        .I1(sbox_input[16]),
        .I2(sbox_input[15]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[8]),
        .O(\aes_cr_reg[2]_0 [11]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[17]_INST_0_i_1 
       (.I0(sbox_input[1]),
        .I1(sbox_input[17]),
        .I2(sbox_input[14]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[9]),
        .O(\aes_cr_reg[2]_0 [12]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[18]_INST_0_i_1 
       (.I0(sbox_input[2]),
        .I1(sbox_input[18]),
        .I2(sbox_input[13]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[10]),
        .O(\aes_cr_reg[2]_0 [13]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[19]_INST_0_i_1 
       (.I0(sbox_input[3]),
        .I1(sbox_input[19]),
        .I2(sbox_input[12]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[11]),
        .O(\aes_cr_reg[2]_0 [14]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[1]_INST_0_i_1 
       (.I0(sbox_input[17]),
        .I1(sbox_input[1]),
        .I2(sbox_input[30]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[25]),
        .O(\aes_cr_reg[2] [0]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[20]_INST_0_i_1 
       (.I0(sbox_input[4]),
        .I1(sbox_input[20]),
        .I2(sbox_input[11]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[12]),
        .O(\aes_cr_reg[2]_0 [15]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[21]_INST_0_i_1 
       (.I0(sbox_input[5]),
        .I1(sbox_input[21]),
        .I2(sbox_input[10]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[13]),
        .O(\aes_cr_reg[2]_0 [16]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[22]_INST_0_i_1 
       (.I0(sbox_input[6]),
        .I1(sbox_input[22]),
        .I2(sbox_input[9]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[14]),
        .O(\aes_cr_reg[2]_0 [17]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[23]_INST_0_i_1 
       (.I0(sbox_input[7]),
        .I1(sbox_input[23]),
        .I2(sbox_input[8]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[15]),
        .O(\aes_cr_reg[2]_0 [18]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[24]_INST_0_i_1 
       (.I0(sbox_input[8]),
        .I1(sbox_input[24]),
        .I2(sbox_input[7]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[0]),
        .O(\aes_cr_reg[2]_0 [19]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[25]_INST_0_i_1 
       (.I0(sbox_input[9]),
        .I1(sbox_input[25]),
        .I2(sbox_input[6]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[1]),
        .O(\aes_cr_reg[2]_0 [20]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[26]_INST_0_i_1 
       (.I0(sbox_input[10]),
        .I1(sbox_input[26]),
        .I2(sbox_input[5]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[2]),
        .O(\aes_cr_reg[2]_0 [21]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[27]_INST_0_i_1 
       (.I0(sbox_input[11]),
        .I1(sbox_input[27]),
        .I2(sbox_input[4]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[3]),
        .O(\aes_cr_reg[2]_0 [22]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[28]_INST_0_i_1 
       (.I0(sbox_input[12]),
        .I1(sbox_input[28]),
        .I2(sbox_input[3]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[4]),
        .O(\aes_cr_reg[2]_0 [23]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[29]_INST_0_i_1 
       (.I0(sbox_input[13]),
        .I1(sbox_input[29]),
        .I2(sbox_input[2]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[5]),
        .O(\aes_cr_reg[2]_0 [24]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[2]_INST_0_i_3 
       (.I0(sbox_input[18]),
        .I1(sbox_input[2]),
        .I2(sbox_input[29]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[26]),
        .O(\aes_cr_reg[2] [1]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[30]_INST_0_i_1 
       (.I0(sbox_input[14]),
        .I1(sbox_input[30]),
        .I2(sbox_input[1]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[6]),
        .O(\aes_cr_reg[2]_0 [25]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[31]_INST_0_i_2 
       (.I0(sbox_input[15]),
        .I1(sbox_input[31]),
        .I2(sbox_input[0]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[7]),
        .O(\aes_cr_reg[2]_0 [26]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[3]_INST_0_i_3 
       (.I0(sbox_input[19]),
        .I1(sbox_input[3]),
        .I2(sbox_input[28]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[27]),
        .O(\aes_cr_reg[2] [2]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[4]_INST_0_i_2 
       (.I0(sbox_input[20]),
        .I1(sbox_input[4]),
        .I2(sbox_input[27]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[28]),
        .O(\aes_cr_reg[2]_0 [0]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[6]_INST_0_i_2 
       (.I0(sbox_input[22]),
        .I1(sbox_input[6]),
        .I2(sbox_input[25]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[30]),
        .O(\aes_cr_reg[2]_0 [1]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[7]_INST_0_i_1 
       (.I0(sbox_input[23]),
        .I1(sbox_input[7]),
        .I2(sbox_input[24]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[31]),
        .O(\aes_cr_reg[2]_0 [2]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[8]_INST_0_i_1 
       (.I0(sbox_input[24]),
        .I1(sbox_input[8]),
        .I2(sbox_input[23]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[16]),
        .O(\aes_cr_reg[2]_0 [3]));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \info_o[9]_INST_0_i_2 
       (.I0(sbox_input[25]),
        .I1(sbox_input[9]),
        .I2(sbox_input[22]),
        .I3(\info_o[1] [1]),
        .I4(\info_o[1] [0]),
        .I5(sbox_input[17]),
        .O(\aes_cr_reg[2]_0 [4]));
endmodule

(* ORIG_REF_NAME = "datapath" *) 
module switch_elements_datapath
   (key_sel_pp1,
    rk_out_sel_pp2,
    \aes_cr_reg[0] ,
    enable_i_0_sp_1,
    \aes_cr_reg[2] ,
    enable_i_6_sp_1,
    enable_i_3_sp_1,
    \enable_i[6]_0 ,
    enable_i_2_sp_1,
    \round_pp1_reg[0]_0 ,
    \round_pp1_reg[3]_0 ,
    \round_pp1_reg[3]_1 ,
    \round_pp1_reg[0]_1 ,
    \round_pp1_reg[3]_2 ,
    key_out,
    \round_pp1_reg[0]_2 ,
    p_16_in,
    sbox_out_enc,
    isomorphism_inv_return03_out,
    p_93_in,
    isomorphism_inv_return033_out,
    isomorphism_inv_return05_out,
    p_86_in,
    p_16_in_0,
    \KR[1].key_reg[2][10]_0 ,
    isomorphism_inv_return03_out_1,
    p_93_in_2,
    isomorphism_inv_return033_out_3,
    isomorphism_inv_return05_out_4,
    p_86_in_5,
    \KR[1].key_reg[2][11]_0 ,
    \KR[1].key_reg[2][12]_0 ,
    \KR[1].key_reg[2][9]_0 ,
    p_16_in_6,
    isomorphism_inv_return03_out_7,
    p_93_in_8,
    \KR[1].key_reg[2][6]_0 ,
    isomorphism_inv_return033_out_9,
    isomorphism_inv_return05_out_10,
    p_86_in_11,
    \KR[1].key_reg[2][4]_0 ,
    enable_i_16_sp_1,
    bus_swap,
    enable_i_17_sp_1,
    enable_i_18_sp_1,
    enable_i_19_sp_1,
    enable_i_20_sp_1,
    enable_i_21_sp_1,
    enable_i_22_sp_1,
    enable_i_23_sp_1,
    data_in,
    enable_i_24_sp_1,
    \IV_BKP_REGISTERS[3].bkp_reg[3][8]_0 ,
    enable_i_25_sp_1,
    \IV_BKP_REGISTERS[3].bkp_reg[3][9]_0 ,
    enable_i_26_sp_1,
    enable_i_27_sp_1,
    enable_i_28_sp_1,
    enable_i_29_sp_1,
    enable_i_30_sp_1,
    \IV_BKP_REGISTERS[3].bkp_reg[3][14]_0 ,
    enable_i_31_sp_1,
    \IV_BKP_REGISTERS[3].bkp_reg[3][15]_0 ,
    \enable_i[0]_0 ,
    enable_i_1_sp_1,
    \enable_i[2]_0 ,
    \enable_i[3]_0 ,
    enable_i_4_sp_1,
    enable_i_5_sp_1,
    \enable_i[6]_1 ,
    enable_i_7_sp_1,
    enable_i_8_sp_1,
    \IV_BKP_REGISTERS[3].bkp_reg[3][24]_0 ,
    enable_i_9_sp_1,
    \IV_BKP_REGISTERS[3].bkp_reg[3][25]_0 ,
    enable_i_10_sp_1,
    \IV_BKP_REGISTERS[3].bkp_reg[3][26]_0 ,
    enable_i_11_sp_1,
    \IV_BKP_REGISTERS[3].bkp_reg[3][27]_0 ,
    enable_i_12_sp_1,
    enable_i_13_sp_1,
    \IV_BKP_REGISTERS[3].bkp_reg[3][29]_0 ,
    enable_i_14_sp_1,
    \IV_BKP_REGISTERS[3].bkp_reg[3][30]_0 ,
    enable_i_15_sp_1,
    \IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 ,
    key_in,
    g_func,
    add_rk_out,
    \CD[2].col_reg[1][0]_0 ,
    Q,
    \CD[3].col_reg[0][31]_0 ,
    last_round_pp2_reg_0,
    \CD[2].col_reg[1][1]_0 ,
    \CD[2].col_reg[1][6]_0 ,
    \CD[2].col_reg[1][14]_0 ,
    \CD[2].col_reg[1][30]_0 ,
    \CD[2].col_reg[1][5]_0 ,
    \CD[2].col_reg[1][13]_0 ,
    \CD[2].col_reg[1][29]_0 ,
    \CD[2].col_reg[1][9]_0 ,
    \CD[2].col_reg[1][25]_0 ,
    \CD[2].col_reg[1][8]_0 ,
    \CD[2].col_reg[1][24]_0 ,
    \CD[2].col_reg[1][22]_0 ,
    \CD[2].col_reg[1][21]_0 ,
    \CD[2].col_reg[1][17]_0 ,
    \CD[2].col_reg[1][16]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][5]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][31]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][0]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][1]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][2]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][3]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][4]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][5]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][6]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][7]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][10]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][11]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][12]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][13]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][16]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][17]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][18]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][19]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][20]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][21]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][22]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][23]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][28]_0 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][1]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][2]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][3]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][4]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][6]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][7]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][8]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][9]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][10]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][11]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][12]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][13]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][14]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][15]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][16]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][17]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][18]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][19]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][20]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][21]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][22]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][23]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][24]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][25]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][26]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][27]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][28]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][29]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][30]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][31]_1 ,
    \key_out_sel_pp1_reg[1]_0 ,
    \key_out_sel_pp2_reg[1]_0 ,
    \CD[2].col_reg[1][31]_0 ,
    \CD[1].col_reg[2][31]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][5]_1 ,
    \IV_BKP_REGISTERS[2].iv_reg[2][31]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][0]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][1]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][2]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][3]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][4]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][6]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][7]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][8]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][9]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][14]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][15]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][16]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][17]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][18]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][19]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][20]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][21]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][22]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][23]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][24]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][25]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][26]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][27]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][29]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][30]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][31]_2 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][0]_1 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][16]_2 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][24]_2 ,
    O,
    \aes_cr_reg[2]_0 ,
    \key_en_pp1_reg[3]_0 ,
    \KR[2].key_host_reg[1][31]_0 ,
    \col_en_cnt_unit_pp2_reg[3]_0 ,
    \IV_BKP_REGISTERS[1].iv_reg[1][31]_0 ,
    \IV_BKP_REGISTERS[0].iv_reg[0][31]_0 ,
    \col_sel_pp2_reg[1]_0 ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 ,
    key_sel,
    clk_i,
    rst_i,
    last_round,
    rk_out_sel,
    \info_o[0] ,
    \info_o[0]_0 ,
    \info_o[0]_1 ,
    \info_o[0]_2 ,
    enable_i,
    enc_dec_sbox,
    \sbox_pp2_reg[31]_0 ,
    \CD[0].col[3][0]_i_2 ,
    add_rk_sel,
    \IV_BKP_REGISTERS[0].bkp_reg[0][8]_0 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][8]_1 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][9]_0 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][9]_1 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][14]_0 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][14]_1 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][15]_0 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][15]_1 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][24]_0 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][24]_1 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][25]_0 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][25]_1 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][26]_0 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][26]_1 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][27]_0 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][27]_1 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][29]_0 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][29]_1 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][30]_0 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][30]_1 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][31]_2 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][31]_3 ,
    key_en,
    key_sel_mux,
    \CD[0].col[3][0]_i_6_0 ,
    \base_new_pp_reg[4] ,
    \info_o[28]_INST_0_i_7 ,
    \info_o[28]_INST_0_i_7_0 ,
    \CD[0].col[3][7]_i_7_0 ,
    \CD[0].col[3][15]_i_11_0 ,
    \CD[0].col[3][31]_i_12_0 ,
    \CD[0].col[3][1]_i_6_0 ,
    \base_new_pp_reg[4]_0 ,
    \base_new_pp_reg[4]_1 ,
    \base_new_pp_reg[4]_2 ,
    \CD[0].col[3][2]_i_6_0 ,
    \CD[0].col[3][5]_i_6_0 ,
    \CD[0].col[3][13]_i_8_0 ,
    \CD[0].col[3][29]_i_6_0 ,
    \base_new_pp_reg[3] ,
    \CD[0].col[3][4]_i_6_0 ,
    \CD[0].col[3][12]_i_8_0 ,
    \CD[0].col[3][28]_i_6_0 ,
    \base_new_pp_reg[3]_0 ,
    \base_new_pp_reg[3]_1 ,
    \CD[0].col[3][10]_i_8_0 ,
    \CD[0].col[3][26]_i_6_0 ,
    \CD[0].col[3][9]_i_8_0 ,
    \CD[0].col[3][25]_i_6_0 ,
    \CD[0].col[3][8]_i_8_0 ,
    \CD[0].col[3][24]_i_6_0 ,
    \CD[0].col[3][23]_i_7_0 ,
    \base_new_pp_reg[4]_3 ,
    \CD[0].col[3][21]_i_6_0 ,
    \CD[0].col[3][20]_i_6_0 ,
    \base_new_pp_reg[3]_2 ,
    \CD[0].col[3][18]_i_6_0 ,
    \CD[0].col[3][17]_i_6_0 ,
    \CD[0].col[3][16]_i_6_0 ,
    \CD[0].col[3][9]_i_8_1 ,
    \CD[0].col[3][5]_i_7 ,
    \CD[0].col[3][0]_i_2_0 ,
    \CD[0].col[3][31]_i_5 ,
    \IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ,
    \IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ,
    \sbox_pp2_reg[5]_0 ,
    key_sel_rd,
    D,
    bypass_key_en,
    key_derivation_en,
    \CD[0].col[3][7]_i_9_0 ,
    \CD[0].col[3][7]_i_9_1 ,
    iv_mux_out13_out,
    isomorphism_return179_out,
    isomorphism_return114_out,
    isomorphism_return179_out_12,
    isomorphism_return114_out_13,
    isomorphism_return179_out_14,
    isomorphism_return114_out_15,
    isomorphism_return179_out_16,
    isomorphism_return114_out_17,
    \info_o[1] ,
    E,
    \key_en_pp1_reg[3]_1 ,
    \KR[0].key_host_reg[3][0]_0 ,
    \KR[0].key_reg[3][31]_0 ,
    \KR[1].key_host_reg[2][0]_0 ,
    \KR[1].key_reg[2][31]_0 ,
    \KR[2].key_host_reg[1][0]_0 ,
    \KR[2].key_reg[1][31]_0 ,
    \KR[2].key_reg[1][31]_1 ,
    \KR[3].key_host_reg[0][0]_0 ,
    \KR[3].key_reg[0][31]_0 ,
    \col_en_cnt_unit_pp1_reg[0]_0 ,
    \col_en_cnt_unit_pp1_reg[3]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][31]_3 ,
    iv_en,
    \CD[0].col_reg[3][31]_0 ,
    \CD[0].col_reg[3][31]_1 ,
    \CD[1].col_reg[2][31]_1 ,
    \CD[1].col_reg[2][31]_2 ,
    \CD[2].col_reg[1][31]_1 ,
    \CD[2].col_reg[1][31]_2 ,
    \CD[3].col_reg[0][31]_1 ,
    \CD[3].col_reg[0][31]_2 ,
    \col_sel_pp1_reg[1]_0 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 ,
    \rk_sel_pp1_reg[1]_0 ,
    \round_pp1_reg[3]_3 );
  output key_sel_pp1;
  output rk_out_sel_pp2;
  output \aes_cr_reg[0] ;
  output enable_i_0_sp_1;
  output [26:0]\aes_cr_reg[2] ;
  output enable_i_6_sp_1;
  output enable_i_3_sp_1;
  output \enable_i[6]_0 ;
  output enable_i_2_sp_1;
  output \round_pp1_reg[0]_0 ;
  output \round_pp1_reg[3]_0 ;
  output \round_pp1_reg[3]_1 ;
  output \round_pp1_reg[0]_1 ;
  output \round_pp1_reg[3]_2 ;
  output [21:0]key_out;
  output \round_pp1_reg[0]_2 ;
  output p_16_in;
  output [5:0]sbox_out_enc;
  output isomorphism_inv_return03_out;
  output p_93_in;
  output isomorphism_inv_return033_out;
  output isomorphism_inv_return05_out;
  output p_86_in;
  output p_16_in_0;
  output \KR[1].key_reg[2][10]_0 ;
  output isomorphism_inv_return03_out_1;
  output p_93_in_2;
  output isomorphism_inv_return033_out_3;
  output isomorphism_inv_return05_out_4;
  output p_86_in_5;
  output \KR[1].key_reg[2][11]_0 ;
  output \KR[1].key_reg[2][12]_0 ;
  output \KR[1].key_reg[2][9]_0 ;
  output p_16_in_6;
  output isomorphism_inv_return03_out_7;
  output p_93_in_8;
  output \KR[1].key_reg[2][6]_0 ;
  output isomorphism_inv_return033_out_9;
  output isomorphism_inv_return05_out_10;
  output p_86_in_11;
  output \KR[1].key_reg[2][4]_0 ;
  output enable_i_16_sp_1;
  output [31:0]bus_swap;
  output enable_i_17_sp_1;
  output enable_i_18_sp_1;
  output enable_i_19_sp_1;
  output enable_i_20_sp_1;
  output enable_i_21_sp_1;
  output enable_i_22_sp_1;
  output enable_i_23_sp_1;
  output [10:0]data_in;
  output enable_i_24_sp_1;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][8]_0 ;
  output enable_i_25_sp_1;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][9]_0 ;
  output enable_i_26_sp_1;
  output enable_i_27_sp_1;
  output enable_i_28_sp_1;
  output enable_i_29_sp_1;
  output enable_i_30_sp_1;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][14]_0 ;
  output enable_i_31_sp_1;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][15]_0 ;
  output \enable_i[0]_0 ;
  output enable_i_1_sp_1;
  output \enable_i[2]_0 ;
  output \enable_i[3]_0 ;
  output enable_i_4_sp_1;
  output enable_i_5_sp_1;
  output \enable_i[6]_1 ;
  output enable_i_7_sp_1;
  output enable_i_8_sp_1;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][24]_0 ;
  output enable_i_9_sp_1;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][25]_0 ;
  output enable_i_10_sp_1;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][26]_0 ;
  output enable_i_11_sp_1;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][27]_0 ;
  output enable_i_12_sp_1;
  output enable_i_13_sp_1;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][29]_0 ;
  output enable_i_14_sp_1;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][30]_0 ;
  output enable_i_15_sp_1;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 ;
  output [127:0]key_in;
  output [1:0]g_func;
  output [15:0]add_rk_out;
  output \CD[2].col_reg[1][0]_0 ;
  output [31:0]Q;
  output [31:0]\CD[3].col_reg[0][31]_0 ;
  output [15:0]last_round_pp2_reg_0;
  output \CD[2].col_reg[1][1]_0 ;
  output \CD[2].col_reg[1][6]_0 ;
  output \CD[2].col_reg[1][14]_0 ;
  output \CD[2].col_reg[1][30]_0 ;
  output \CD[2].col_reg[1][5]_0 ;
  output \CD[2].col_reg[1][13]_0 ;
  output \CD[2].col_reg[1][29]_0 ;
  output \CD[2].col_reg[1][9]_0 ;
  output \CD[2].col_reg[1][25]_0 ;
  output \CD[2].col_reg[1][8]_0 ;
  output \CD[2].col_reg[1][24]_0 ;
  output \CD[2].col_reg[1][22]_0 ;
  output \CD[2].col_reg[1][21]_0 ;
  output \CD[2].col_reg[1][17]_0 ;
  output \CD[2].col_reg[1][16]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][5]_0 ;
  output [27:0]\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][0]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][1]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][2]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][3]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][4]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][5]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][6]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][7]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][10]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][11]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][12]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][13]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][16]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][17]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][18]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][19]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][20]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][21]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][22]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][23]_0 ;
  output \IV_BKP_REGISTERS[3].bkp_reg[3][28]_0 ;
  output [31:0]\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 ;
  output [31:0]\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][1]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][2]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][3]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][4]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][6]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][7]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][8]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][9]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][10]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][11]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][12]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][13]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][14]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][15]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][16]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][17]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][18]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][19]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][20]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][21]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][22]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][23]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][24]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][25]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][26]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][27]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][28]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][29]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][30]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][31]_1 ;
  output [0:0]\key_out_sel_pp1_reg[1]_0 ;
  output [0:0]\key_out_sel_pp2_reg[1]_0 ;
  output [31:0]\CD[2].col_reg[1][31]_0 ;
  output [31:0]\CD[1].col_reg[2][31]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][5]_1 ;
  output [31:0]\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][0]_0 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][1]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][2]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][3]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][4]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][6]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][7]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][8]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][9]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][14]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][15]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][16]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][17]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][18]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][19]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][20]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][21]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][22]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][23]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][24]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][25]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][26]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][27]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][29]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][30]_1 ;
  output \IV_BKP_REGISTERS[3].iv_reg[3][31]_2 ;
  output [7:0]\IV_BKP_REGISTERS[3].iv_reg[3][0]_1 ;
  output [7:0]\IV_BKP_REGISTERS[3].iv_reg[3][16]_2 ;
  output [7:0]\IV_BKP_REGISTERS[3].iv_reg[3][24]_2 ;
  output [6:0]O;
  output [2:0]\aes_cr_reg[2]_0 ;
  output [3:0]\key_en_pp1_reg[3]_0 ;
  output [31:0]\KR[2].key_host_reg[1][31]_0 ;
  output [3:0]\col_en_cnt_unit_pp2_reg[3]_0 ;
  output [31:0]\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 ;
  output [31:0]\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 ;
  output [1:0]\col_sel_pp2_reg[1]_0 ;
  output [31:0]\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 ;
  output [31:0]\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 ;
  output [31:0]\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 ;
  output [31:0]\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 ;
  input key_sel;
  input clk_i;
  input rst_i;
  input last_round;
  input rk_out_sel;
  input \info_o[0] ;
  input \info_o[0]_0 ;
  input \info_o[0]_1 ;
  input \info_o[0]_2 ;
  input [31:0]enable_i;
  input enc_dec_sbox;
  input \sbox_pp2_reg[31]_0 ;
  input \CD[0].col[3][0]_i_2 ;
  input add_rk_sel;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][8]_0 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][8]_1 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][9]_0 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][9]_1 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][14]_0 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][14]_1 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][15]_0 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][15]_1 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][24]_0 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][24]_1 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][25]_0 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][25]_1 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][26]_0 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][26]_1 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][27]_0 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][27]_1 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][29]_0 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][29]_1 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][30]_0 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][30]_1 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][31]_2 ;
  input \IV_BKP_REGISTERS[1].bkp_reg[1][31]_3 ;
  input [2:0]key_en;
  input key_sel_mux;
  input \CD[0].col[3][0]_i_6_0 ;
  input \base_new_pp_reg[4] ;
  input \info_o[28]_INST_0_i_7 ;
  input \info_o[28]_INST_0_i_7_0 ;
  input \CD[0].col[3][7]_i_7_0 ;
  input \CD[0].col[3][15]_i_11_0 ;
  input \CD[0].col[3][31]_i_12_0 ;
  input \CD[0].col[3][1]_i_6_0 ;
  input \base_new_pp_reg[4]_0 ;
  input \base_new_pp_reg[4]_1 ;
  input \base_new_pp_reg[4]_2 ;
  input \CD[0].col[3][2]_i_6_0 ;
  input \CD[0].col[3][5]_i_6_0 ;
  input \CD[0].col[3][13]_i_8_0 ;
  input \CD[0].col[3][29]_i_6_0 ;
  input \base_new_pp_reg[3] ;
  input \CD[0].col[3][4]_i_6_0 ;
  input \CD[0].col[3][12]_i_8_0 ;
  input \CD[0].col[3][28]_i_6_0 ;
  input \base_new_pp_reg[3]_0 ;
  input \base_new_pp_reg[3]_1 ;
  input \CD[0].col[3][10]_i_8_0 ;
  input \CD[0].col[3][26]_i_6_0 ;
  input \CD[0].col[3][9]_i_8_0 ;
  input \CD[0].col[3][25]_i_6_0 ;
  input \CD[0].col[3][8]_i_8_0 ;
  input \CD[0].col[3][24]_i_6_0 ;
  input \CD[0].col[3][23]_i_7_0 ;
  input \base_new_pp_reg[4]_3 ;
  input \CD[0].col[3][21]_i_6_0 ;
  input \CD[0].col[3][20]_i_6_0 ;
  input \base_new_pp_reg[3]_2 ;
  input \CD[0].col[3][18]_i_6_0 ;
  input \CD[0].col[3][17]_i_6_0 ;
  input \CD[0].col[3][16]_i_6_0 ;
  input [1:0]\CD[0].col[3][9]_i_8_1 ;
  input \CD[0].col[3][5]_i_7 ;
  input \CD[0].col[3][0]_i_2_0 ;
  input \CD[0].col[3][31]_i_5 ;
  input \IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ;
  input \IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ;
  input \sbox_pp2_reg[5]_0 ;
  input [0:0]key_sel_rd;
  input [1:0]D;
  input bypass_key_en;
  input key_derivation_en;
  input \CD[0].col[3][7]_i_9_0 ;
  input \CD[0].col[3][7]_i_9_1 ;
  input iv_mux_out13_out;
  input isomorphism_return179_out;
  input isomorphism_return114_out;
  input isomorphism_return179_out_12;
  input isomorphism_return114_out_13;
  input isomorphism_return179_out_14;
  input isomorphism_return114_out_15;
  input isomorphism_return179_out_16;
  input isomorphism_return114_out_17;
  input [1:0]\info_o[1] ;
  input [0:0]E;
  input [3:0]\key_en_pp1_reg[3]_1 ;
  input [0:0]\KR[0].key_host_reg[3][0]_0 ;
  input [0:0]\KR[0].key_reg[3][31]_0 ;
  input [0:0]\KR[1].key_host_reg[2][0]_0 ;
  input [0:0]\KR[1].key_reg[2][31]_0 ;
  input [0:0]\KR[2].key_host_reg[1][0]_0 ;
  input [0:0]\KR[2].key_reg[1][31]_0 ;
  input [31:0]\KR[2].key_reg[1][31]_1 ;
  input [0:0]\KR[3].key_host_reg[0][0]_0 ;
  input [0:0]\KR[3].key_reg[0][31]_0 ;
  input [0:0]\col_en_cnt_unit_pp1_reg[0]_0 ;
  input [3:0]\col_en_cnt_unit_pp1_reg[3]_0 ;
  input [0:0]\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ;
  input [31:0]\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 ;
  input [2:0]iv_en;
  input [0:0]\CD[0].col_reg[3][31]_0 ;
  input [31:0]\CD[0].col_reg[3][31]_1 ;
  input [0:0]\CD[1].col_reg[2][31]_1 ;
  input [31:0]\CD[1].col_reg[2][31]_2 ;
  input [0:0]\CD[2].col_reg[1][31]_1 ;
  input [31:0]\CD[2].col_reg[1][31]_2 ;
  input [0:0]\CD[3].col_reg[0][31]_1 ;
  input [31:0]\CD[3].col_reg[0][31]_2 ;
  input [1:0]\col_sel_pp1_reg[1]_0 ;
  input [0:0]\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ;
  input [31:0]\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 ;
  input [0:0]\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ;
  input [31:0]\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 ;
  input [0:0]\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ;
  input [31:0]\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 ;
  input [0:0]\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ;
  input [31:0]\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 ;
  input [1:0]\rk_sel_pp1_reg[1]_0 ;
  input [3:0]\round_pp1_reg[3]_3 ;

  wire \CD[0].col[3][0]_i_12_n_0 ;
  wire \CD[0].col[3][0]_i_15_n_0 ;
  wire \CD[0].col[3][0]_i_16_n_0 ;
  wire \CD[0].col[3][0]_i_2 ;
  wire \CD[0].col[3][0]_i_2_0 ;
  wire \CD[0].col[3][0]_i_6_0 ;
  wire \CD[0].col[3][10]_i_11_n_0 ;
  wire \CD[0].col[3][10]_i_14_n_0 ;
  wire \CD[0].col[3][10]_i_8_0 ;
  wire \CD[0].col[3][11]_i_10_n_0 ;
  wire \CD[0].col[3][11]_i_11_n_0 ;
  wire \CD[0].col[3][11]_i_12_n_0 ;
  wire \CD[0].col[3][11]_i_15_n_0 ;
  wire \CD[0].col[3][11]_i_16_n_0 ;
  wire \CD[0].col[3][11]_i_17_n_0 ;
  wire \CD[0].col[3][12]_i_11_n_0 ;
  wire \CD[0].col[3][12]_i_12_n_0 ;
  wire \CD[0].col[3][12]_i_13_n_0 ;
  wire \CD[0].col[3][12]_i_16_n_0 ;
  wire \CD[0].col[3][12]_i_18_n_0 ;
  wire \CD[0].col[3][12]_i_19_n_0 ;
  wire \CD[0].col[3][12]_i_8_0 ;
  wire \CD[0].col[3][13]_i_10_n_0 ;
  wire \CD[0].col[3][13]_i_13_n_0 ;
  wire \CD[0].col[3][13]_i_8_0 ;
  wire \CD[0].col[3][14]_i_10_n_0 ;
  wire \CD[0].col[3][14]_i_13_n_0 ;
  wire \CD[0].col[3][14]_i_16_n_0 ;
  wire \CD[0].col[3][15]_i_11_0 ;
  wire \CD[0].col[3][15]_i_14_n_0 ;
  wire \CD[0].col[3][15]_i_15_n_0 ;
  wire \CD[0].col[3][15]_i_18_n_0 ;
  wire \CD[0].col[3][15]_i_22_n_0 ;
  wire \CD[0].col[3][16]_i_10_n_0 ;
  wire \CD[0].col[3][16]_i_13_n_0 ;
  wire \CD[0].col[3][16]_i_6_0 ;
  wire \CD[0].col[3][17]_i_10_n_0 ;
  wire \CD[0].col[3][17]_i_6_0 ;
  wire \CD[0].col[3][18]_i_10_n_0 ;
  wire \CD[0].col[3][18]_i_6_0 ;
  wire \CD[0].col[3][19]_i_10_n_0 ;
  wire \CD[0].col[3][19]_i_13_n_0 ;
  wire \CD[0].col[3][1]_i_13_n_0 ;
  wire \CD[0].col[3][1]_i_16_n_0 ;
  wire \CD[0].col[3][1]_i_17_n_0 ;
  wire \CD[0].col[3][1]_i_6_0 ;
  wire \CD[0].col[3][20]_i_10_n_0 ;
  wire \CD[0].col[3][20]_i_13_n_0 ;
  wire \CD[0].col[3][20]_i_6_0 ;
  wire \CD[0].col[3][21]_i_10_n_0 ;
  wire \CD[0].col[3][21]_i_13_n_0 ;
  wire \CD[0].col[3][21]_i_6_0 ;
  wire \CD[0].col[3][22]_i_10_n_0 ;
  wire \CD[0].col[3][23]_i_11_n_0 ;
  wire \CD[0].col[3][23]_i_14_n_0 ;
  wire \CD[0].col[3][23]_i_7_0 ;
  wire \CD[0].col[3][24]_i_12_n_0 ;
  wire \CD[0].col[3][24]_i_15_n_0 ;
  wire \CD[0].col[3][24]_i_16_n_0 ;
  wire \CD[0].col[3][24]_i_17_n_0 ;
  wire \CD[0].col[3][24]_i_18_n_0 ;
  wire \CD[0].col[3][24]_i_19_n_0 ;
  wire \CD[0].col[3][24]_i_6_0 ;
  wire \CD[0].col[3][25]_i_12_n_0 ;
  wire \CD[0].col[3][25]_i_15_n_0 ;
  wire \CD[0].col[3][25]_i_6_0 ;
  wire \CD[0].col[3][26]_i_12_n_0 ;
  wire \CD[0].col[3][26]_i_16_n_0 ;
  wire \CD[0].col[3][26]_i_17_n_0 ;
  wire \CD[0].col[3][26]_i_18_n_0 ;
  wire \CD[0].col[3][26]_i_19_n_0 ;
  wire \CD[0].col[3][26]_i_21_n_0 ;
  wire \CD[0].col[3][26]_i_22_n_0 ;
  wire \CD[0].col[3][26]_i_6_0 ;
  wire \CD[0].col[3][27]_i_12_n_0 ;
  wire \CD[0].col[3][27]_i_15_n_0 ;
  wire \CD[0].col[3][27]_i_16_n_0 ;
  wire \CD[0].col[3][27]_i_17_n_0 ;
  wire \CD[0].col[3][27]_i_18_n_0 ;
  wire \CD[0].col[3][27]_i_19_n_0 ;
  wire \CD[0].col[3][27]_i_20_n_0 ;
  wire \CD[0].col[3][27]_i_21_n_0 ;
  wire \CD[0].col[3][28]_i_12_n_0 ;
  wire \CD[0].col[3][28]_i_14_n_0 ;
  wire \CD[0].col[3][28]_i_15_n_0 ;
  wire \CD[0].col[3][28]_i_16_n_0 ;
  wire \CD[0].col[3][28]_i_17_n_0 ;
  wire \CD[0].col[3][28]_i_19_n_0 ;
  wire \CD[0].col[3][28]_i_6_0 ;
  wire \CD[0].col[3][29]_i_12_n_0 ;
  wire \CD[0].col[3][29]_i_15_n_0 ;
  wire \CD[0].col[3][29]_i_16_n_0 ;
  wire \CD[0].col[3][29]_i_17_n_0 ;
  wire \CD[0].col[3][29]_i_18_n_0 ;
  wire \CD[0].col[3][29]_i_19_n_0 ;
  wire \CD[0].col[3][29]_i_20_n_0 ;
  wire \CD[0].col[3][29]_i_6_0 ;
  wire \CD[0].col[3][2]_i_13_n_0 ;
  wire \CD[0].col[3][2]_i_17_n_0 ;
  wire \CD[0].col[3][2]_i_18_n_0 ;
  wire \CD[0].col[3][2]_i_19_n_0 ;
  wire \CD[0].col[3][2]_i_21_n_0 ;
  wire \CD[0].col[3][2]_i_6_0 ;
  wire \CD[0].col[3][30]_i_12_n_0 ;
  wire \CD[0].col[3][30]_i_15_n_0 ;
  wire \CD[0].col[3][30]_i_16_n_0 ;
  wire \CD[0].col[3][30]_i_17_n_0 ;
  wire \CD[0].col[3][30]_i_18_n_0 ;
  wire \CD[0].col[3][30]_i_19_n_0 ;
  wire \CD[0].col[3][31]_i_12_0 ;
  wire \CD[0].col[3][31]_i_25_n_0 ;
  wire \CD[0].col[3][31]_i_29_n_0 ;
  wire \CD[0].col[3][31]_i_31_n_0 ;
  wire \CD[0].col[3][31]_i_32_n_0 ;
  wire \CD[0].col[3][31]_i_33_n_0 ;
  wire \CD[0].col[3][31]_i_34_n_0 ;
  wire \CD[0].col[3][31]_i_35_n_0 ;
  wire \CD[0].col[3][31]_i_37_n_0 ;
  wire \CD[0].col[3][31]_i_39_n_0 ;
  wire \CD[0].col[3][31]_i_5 ;
  wire \CD[0].col[3][3]_i_13_n_0 ;
  wire \CD[0].col[3][3]_i_16_n_0 ;
  wire \CD[0].col[3][3]_i_17_n_0 ;
  wire \CD[0].col[3][3]_i_18_n_0 ;
  wire \CD[0].col[3][3]_i_19_n_0 ;
  wire \CD[0].col[3][4]_i_12_n_0 ;
  wire \CD[0].col[3][4]_i_16_n_0 ;
  wire \CD[0].col[3][4]_i_17_n_0 ;
  wire \CD[0].col[3][4]_i_19_n_0 ;
  wire \CD[0].col[3][4]_i_6_0 ;
  wire \CD[0].col[3][5]_i_13_n_0 ;
  wire \CD[0].col[3][5]_i_16_n_0 ;
  wire \CD[0].col[3][5]_i_17_n_0 ;
  wire \CD[0].col[3][5]_i_18_n_0 ;
  wire \CD[0].col[3][5]_i_19_n_0 ;
  wire \CD[0].col[3][5]_i_20_n_0 ;
  wire \CD[0].col[3][5]_i_21_n_0 ;
  wire \CD[0].col[3][5]_i_6_0 ;
  wire \CD[0].col[3][5]_i_7 ;
  wire \CD[0].col[3][6]_i_12_n_0 ;
  wire \CD[0].col[3][6]_i_15_n_0 ;
  wire \CD[0].col[3][6]_i_16_n_0 ;
  wire \CD[0].col[3][6]_i_17_n_0 ;
  wire \CD[0].col[3][7]_i_13_n_0 ;
  wire \CD[0].col[3][7]_i_17_n_0 ;
  wire \CD[0].col[3][7]_i_18_n_0 ;
  wire \CD[0].col[3][7]_i_19_n_0 ;
  wire \CD[0].col[3][7]_i_7_0 ;
  wire \CD[0].col[3][7]_i_9_0 ;
  wire \CD[0].col[3][7]_i_9_1 ;
  wire \CD[0].col[3][8]_i_10_n_0 ;
  wire \CD[0].col[3][8]_i_11_n_0 ;
  wire \CD[0].col[3][8]_i_14_n_0 ;
  wire \CD[0].col[3][8]_i_17_n_0 ;
  wire \CD[0].col[3][8]_i_8_0 ;
  wire \CD[0].col[3][9]_i_10_n_0 ;
  wire \CD[0].col[3][9]_i_13_n_0 ;
  wire \CD[0].col[3][9]_i_8_0 ;
  wire [1:0]\CD[0].col[3][9]_i_8_1 ;
  wire [0:0]\CD[0].col_reg[3][31]_0 ;
  wire [31:0]\CD[0].col_reg[3][31]_1 ;
  wire \CD[1].col[2][16]_i_5_n_0 ;
  wire \CD[1].col[2][17]_i_5_n_0 ;
  wire \CD[1].col[2][18]_i_6_n_0 ;
  wire \CD[1].col[2][19]_i_5_n_0 ;
  wire \CD[1].col[2][20]_i_6_n_0 ;
  wire \CD[1].col[2][20]_i_7_n_0 ;
  wire \CD[1].col[2][20]_i_8_n_0 ;
  wire \CD[1].col[2][21]_i_5_n_0 ;
  wire \CD[1].col[2][21]_i_6_n_0 ;
  wire \CD[1].col[2][21]_i_7_n_0 ;
  wire \CD[1].col[2][22]_i_5_n_0 ;
  wire \CD[1].col[2][23]_i_6_n_0 ;
  wire [31:0]\CD[1].col_reg[2][31]_0 ;
  wire [0:0]\CD[1].col_reg[2][31]_1 ;
  wire [31:0]\CD[1].col_reg[2][31]_2 ;
  wire \CD[2].col_reg[1][0]_0 ;
  wire \CD[2].col_reg[1][13]_0 ;
  wire \CD[2].col_reg[1][14]_0 ;
  wire \CD[2].col_reg[1][16]_0 ;
  wire \CD[2].col_reg[1][17]_0 ;
  wire \CD[2].col_reg[1][1]_0 ;
  wire \CD[2].col_reg[1][21]_0 ;
  wire \CD[2].col_reg[1][22]_0 ;
  wire \CD[2].col_reg[1][24]_0 ;
  wire \CD[2].col_reg[1][25]_0 ;
  wire \CD[2].col_reg[1][29]_0 ;
  wire \CD[2].col_reg[1][30]_0 ;
  wire [31:0]\CD[2].col_reg[1][31]_0 ;
  wire [0:0]\CD[2].col_reg[1][31]_1 ;
  wire [31:0]\CD[2].col_reg[1][31]_2 ;
  wire \CD[2].col_reg[1][5]_0 ;
  wire \CD[2].col_reg[1][6]_0 ;
  wire \CD[2].col_reg[1][8]_0 ;
  wire \CD[2].col_reg[1][9]_0 ;
  wire [31:0]\CD[3].col_reg[0][31]_0 ;
  wire [0:0]\CD[3].col_reg[0][31]_1 ;
  wire [31:0]\CD[3].col_reg[0][31]_2 ;
  wire [1:0]D;
  wire [0:0]E;
  wire [31:0]\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 ;
  wire [0:0]\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][14]_0 ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][14]_1 ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][15]_0 ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][15]_1 ;
  wire [31:0]\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 ;
  wire [31:0]\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][8]_0 ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][8]_1 ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][9]_0 ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][9]_1 ;
  wire [31:0]\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 ;
  wire [31:0]\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 ;
  wire [0:0]\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][24]_0 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][24]_1 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][25]_0 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][25]_1 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][26]_0 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][26]_1 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][27]_0 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][27]_1 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][29]_0 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][29]_1 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][30]_0 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][30]_1 ;
  wire [31:0]\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][31]_2 ;
  wire \IV_BKP_REGISTERS[1].bkp_reg[1][31]_3 ;
  wire [31:0]\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 ;
  wire [31:0]\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][24]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][25]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][26]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][27]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][29]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][30]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][31]_i_5_n_0 ;
  wire [31:0]\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 ;
  wire [0:0]\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ;
  wire [31:0]\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 ;
  wire [31:0]\IV_BKP_REGISTERS[2].bkp_reg[2]_13 ;
  wire [31:0]\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][14]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][15]_i_7_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][8]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][9]_i_5_n_0 ;
  wire [31:0]\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][0]_0 ;
  wire [0:0]\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][10]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][11]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][12]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][13]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][14]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][15]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][16]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][17]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][18]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][19]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][1]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][20]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][21]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][22]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][23]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][24]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][25]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][26]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][27]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][28]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][29]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][2]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][30]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 ;
  wire [31:0]\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][3]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][4]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][5]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][6]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][7]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][8]_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][9]_0 ;
  wire [31:0]\IV_BKP_REGISTERS[3].bkp_reg[3]_11 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][0]_0 ;
  wire [7:0]\IV_BKP_REGISTERS[3].iv_reg[3][0]_1 ;
  wire [0:0]\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][10]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][11]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][12]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][13]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][14]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][14]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][15]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][15]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][16]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][16]_1 ;
  wire [7:0]\IV_BKP_REGISTERS[3].iv_reg[3][16]_2 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_2 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_3 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_4 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_5 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_6 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_7 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][17]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][17]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][18]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][18]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][19]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][19]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][1]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][1]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][20]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][20]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][21]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][21]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][22]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][22]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][23]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][23]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][24]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][24]_1 ;
  wire [7:0]\IV_BKP_REGISTERS[3].iv_reg[3][24]_2 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_2 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_3 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_4 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_5 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_6 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_7 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][25]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][25]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][26]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][26]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][27]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][27]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][28]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][29]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][29]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][2]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][2]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][30]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][30]_1 ;
  wire [27:0]\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][31]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][31]_2 ;
  wire [31:0]\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_n_2 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_n_3 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_n_4 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_n_5 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_n_6 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_n_7 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][3]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][3]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][4]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][4]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][5]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][5]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][6]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][6]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][7]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][7]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][8]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][8]_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_1 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_2 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_3 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_4 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_5 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_6 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_7 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][9]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][9]_1 ;
  wire [5:1]\IV_BKP_REGISTERS[3].iv_reg[3]_4 ;
  wire [3:2]\KEY_EXPANDER/rc ;
  wire \KR[0].key[3][0]_i_1_n_0 ;
  wire \KR[0].key[3][10]_i_1_n_0 ;
  wire \KR[0].key[3][11]_i_1_n_0 ;
  wire \KR[0].key[3][12]_i_1_n_0 ;
  wire \KR[0].key[3][13]_i_1_n_0 ;
  wire \KR[0].key[3][14]_i_1_n_0 ;
  wire \KR[0].key[3][15]_i_1_n_0 ;
  wire \KR[0].key[3][16]_i_1_n_0 ;
  wire \KR[0].key[3][17]_i_1_n_0 ;
  wire \KR[0].key[3][18]_i_1_n_0 ;
  wire \KR[0].key[3][19]_i_1_n_0 ;
  wire \KR[0].key[3][1]_i_1_n_0 ;
  wire \KR[0].key[3][20]_i_1_n_0 ;
  wire \KR[0].key[3][21]_i_1_n_0 ;
  wire \KR[0].key[3][22]_i_1_n_0 ;
  wire \KR[0].key[3][23]_i_1_n_0 ;
  wire \KR[0].key[3][24]_i_1_n_0 ;
  wire \KR[0].key[3][25]_i_1_n_0 ;
  wire \KR[0].key[3][26]_i_1_n_0 ;
  wire \KR[0].key[3][27]_i_1_n_0 ;
  wire \KR[0].key[3][28]_i_1_n_0 ;
  wire \KR[0].key[3][29]_i_1_n_0 ;
  wire \KR[0].key[3][2]_i_1_n_0 ;
  wire \KR[0].key[3][30]_i_1_n_0 ;
  wire \KR[0].key[3][31]_i_2_n_0 ;
  wire \KR[0].key[3][3]_i_1_n_0 ;
  wire \KR[0].key[3][4]_i_1_n_0 ;
  wire \KR[0].key[3][5]_i_1_n_0 ;
  wire \KR[0].key[3][6]_i_1_n_0 ;
  wire \KR[0].key[3][7]_i_1_n_0 ;
  wire \KR[0].key[3][8]_i_1_n_0 ;
  wire \KR[0].key[3][9]_i_1_n_0 ;
  wire \KR[0].key_host[3][0]_i_1_n_0 ;
  wire \KR[0].key_host[3][10]_i_1_n_0 ;
  wire \KR[0].key_host[3][11]_i_1_n_0 ;
  wire \KR[0].key_host[3][12]_i_1_n_0 ;
  wire \KR[0].key_host[3][13]_i_1_n_0 ;
  wire \KR[0].key_host[3][14]_i_1_n_0 ;
  wire \KR[0].key_host[3][15]_i_1_n_0 ;
  wire \KR[0].key_host[3][16]_i_1_n_0 ;
  wire \KR[0].key_host[3][17]_i_1_n_0 ;
  wire \KR[0].key_host[3][18]_i_1_n_0 ;
  wire \KR[0].key_host[3][19]_i_1_n_0 ;
  wire \KR[0].key_host[3][1]_i_1_n_0 ;
  wire \KR[0].key_host[3][20]_i_1_n_0 ;
  wire \KR[0].key_host[3][21]_i_1_n_0 ;
  wire \KR[0].key_host[3][22]_i_1_n_0 ;
  wire \KR[0].key_host[3][23]_i_1_n_0 ;
  wire \KR[0].key_host[3][24]_i_1_n_0 ;
  wire \KR[0].key_host[3][25]_i_1_n_0 ;
  wire \KR[0].key_host[3][26]_i_1_n_0 ;
  wire \KR[0].key_host[3][27]_i_1_n_0 ;
  wire \KR[0].key_host[3][28]_i_1_n_0 ;
  wire \KR[0].key_host[3][29]_i_1_n_0 ;
  wire \KR[0].key_host[3][2]_i_1_n_0 ;
  wire \KR[0].key_host[3][30]_i_1_n_0 ;
  wire \KR[0].key_host[3][31]_i_2_n_0 ;
  wire \KR[0].key_host[3][3]_i_1_n_0 ;
  wire \KR[0].key_host[3][4]_i_1_n_0 ;
  wire \KR[0].key_host[3][5]_i_1_n_0 ;
  wire \KR[0].key_host[3][6]_i_1_n_0 ;
  wire \KR[0].key_host[3][7]_i_1_n_0 ;
  wire \KR[0].key_host[3][8]_i_1_n_0 ;
  wire \KR[0].key_host[3][9]_i_1_n_0 ;
  wire [0:0]\KR[0].key_host_reg[3][0]_0 ;
  wire [31:0]\KR[0].key_host_reg[3]_0 ;
  wire [0:0]\KR[0].key_reg[3][31]_0 ;
  wire \KR[1].key[2][0]_i_1_n_0 ;
  wire \KR[1].key[2][10]_i_1_n_0 ;
  wire \KR[1].key[2][11]_i_1_n_0 ;
  wire \KR[1].key[2][12]_i_1_n_0 ;
  wire \KR[1].key[2][13]_i_1_n_0 ;
  wire \KR[1].key[2][14]_i_1_n_0 ;
  wire \KR[1].key[2][15]_i_1_n_0 ;
  wire \KR[1].key[2][16]_i_1_n_0 ;
  wire \KR[1].key[2][17]_i_1_n_0 ;
  wire \KR[1].key[2][18]_i_1_n_0 ;
  wire \KR[1].key[2][19]_i_1_n_0 ;
  wire \KR[1].key[2][1]_i_1_n_0 ;
  wire \KR[1].key[2][20]_i_1_n_0 ;
  wire \KR[1].key[2][21]_i_1_n_0 ;
  wire \KR[1].key[2][22]_i_1_n_0 ;
  wire \KR[1].key[2][23]_i_1_n_0 ;
  wire \KR[1].key[2][24]_i_1_n_0 ;
  wire \KR[1].key[2][25]_i_1_n_0 ;
  wire \KR[1].key[2][26]_i_1_n_0 ;
  wire \KR[1].key[2][27]_i_1_n_0 ;
  wire \KR[1].key[2][28]_i_1_n_0 ;
  wire \KR[1].key[2][29]_i_1_n_0 ;
  wire \KR[1].key[2][2]_i_1_n_0 ;
  wire \KR[1].key[2][30]_i_1_n_0 ;
  wire \KR[1].key[2][31]_i_2_n_0 ;
  wire \KR[1].key[2][3]_i_1_n_0 ;
  wire \KR[1].key[2][4]_i_1_n_0 ;
  wire \KR[1].key[2][5]_i_1_n_0 ;
  wire \KR[1].key[2][6]_i_1_n_0 ;
  wire \KR[1].key[2][7]_i_1_n_0 ;
  wire \KR[1].key[2][8]_i_1_n_0 ;
  wire \KR[1].key[2][9]_i_1_n_0 ;
  wire \KR[1].key_host[2][0]_i_1_n_0 ;
  wire \KR[1].key_host[2][10]_i_1_n_0 ;
  wire \KR[1].key_host[2][11]_i_1_n_0 ;
  wire \KR[1].key_host[2][12]_i_1_n_0 ;
  wire \KR[1].key_host[2][13]_i_1_n_0 ;
  wire \KR[1].key_host[2][14]_i_1_n_0 ;
  wire \KR[1].key_host[2][15]_i_1_n_0 ;
  wire \KR[1].key_host[2][16]_i_1_n_0 ;
  wire \KR[1].key_host[2][17]_i_1_n_0 ;
  wire \KR[1].key_host[2][18]_i_1_n_0 ;
  wire \KR[1].key_host[2][19]_i_1_n_0 ;
  wire \KR[1].key_host[2][1]_i_1_n_0 ;
  wire \KR[1].key_host[2][20]_i_1_n_0 ;
  wire \KR[1].key_host[2][21]_i_1_n_0 ;
  wire \KR[1].key_host[2][22]_i_1_n_0 ;
  wire \KR[1].key_host[2][23]_i_1_n_0 ;
  wire \KR[1].key_host[2][24]_i_1_n_0 ;
  wire \KR[1].key_host[2][25]_i_1_n_0 ;
  wire \KR[1].key_host[2][26]_i_1_n_0 ;
  wire \KR[1].key_host[2][27]_i_1_n_0 ;
  wire \KR[1].key_host[2][28]_i_1_n_0 ;
  wire \KR[1].key_host[2][29]_i_1_n_0 ;
  wire \KR[1].key_host[2][2]_i_1_n_0 ;
  wire \KR[1].key_host[2][30]_i_1_n_0 ;
  wire \KR[1].key_host[2][31]_i_2_n_0 ;
  wire \KR[1].key_host[2][3]_i_1_n_0 ;
  wire \KR[1].key_host[2][4]_i_1_n_0 ;
  wire \KR[1].key_host[2][5]_i_1_n_0 ;
  wire \KR[1].key_host[2][6]_i_1_n_0 ;
  wire \KR[1].key_host[2][7]_i_1_n_0 ;
  wire \KR[1].key_host[2][8]_i_1_n_0 ;
  wire \KR[1].key_host[2][9]_i_1_n_0 ;
  wire [0:0]\KR[1].key_host_reg[2][0]_0 ;
  wire [31:0]\KR[1].key_host_reg[2]_1 ;
  wire \KR[1].key_reg[2][10]_0 ;
  wire \KR[1].key_reg[2][11]_0 ;
  wire \KR[1].key_reg[2][12]_0 ;
  wire [0:0]\KR[1].key_reg[2][31]_0 ;
  wire \KR[1].key_reg[2][4]_0 ;
  wire \KR[1].key_reg[2][6]_0 ;
  wire \KR[1].key_reg[2][9]_0 ;
  wire \KR[2].key_host[1][0]_i_1_n_0 ;
  wire \KR[2].key_host[1][10]_i_1_n_0 ;
  wire \KR[2].key_host[1][11]_i_1_n_0 ;
  wire \KR[2].key_host[1][12]_i_1_n_0 ;
  wire \KR[2].key_host[1][13]_i_1_n_0 ;
  wire \KR[2].key_host[1][14]_i_1_n_0 ;
  wire \KR[2].key_host[1][15]_i_1_n_0 ;
  wire \KR[2].key_host[1][16]_i_1_n_0 ;
  wire \KR[2].key_host[1][17]_i_1_n_0 ;
  wire \KR[2].key_host[1][18]_i_1_n_0 ;
  wire \KR[2].key_host[1][19]_i_1_n_0 ;
  wire \KR[2].key_host[1][1]_i_1_n_0 ;
  wire \KR[2].key_host[1][20]_i_1_n_0 ;
  wire \KR[2].key_host[1][21]_i_1_n_0 ;
  wire \KR[2].key_host[1][22]_i_1_n_0 ;
  wire \KR[2].key_host[1][23]_i_1_n_0 ;
  wire \KR[2].key_host[1][24]_i_1_n_0 ;
  wire \KR[2].key_host[1][25]_i_1_n_0 ;
  wire \KR[2].key_host[1][26]_i_1_n_0 ;
  wire \KR[2].key_host[1][27]_i_1_n_0 ;
  wire \KR[2].key_host[1][28]_i_1_n_0 ;
  wire \KR[2].key_host[1][29]_i_1_n_0 ;
  wire \KR[2].key_host[1][2]_i_1_n_0 ;
  wire \KR[2].key_host[1][30]_i_1_n_0 ;
  wire \KR[2].key_host[1][31]_i_2_n_0 ;
  wire \KR[2].key_host[1][3]_i_1_n_0 ;
  wire \KR[2].key_host[1][4]_i_1_n_0 ;
  wire \KR[2].key_host[1][5]_i_1_n_0 ;
  wire \KR[2].key_host[1][6]_i_1_n_0 ;
  wire \KR[2].key_host[1][7]_i_1_n_0 ;
  wire \KR[2].key_host[1][8]_i_1_n_0 ;
  wire \KR[2].key_host[1][9]_i_1_n_0 ;
  wire [0:0]\KR[2].key_host_reg[1][0]_0 ;
  wire [31:0]\KR[2].key_host_reg[1][31]_0 ;
  wire [0:0]\KR[2].key_reg[1][31]_0 ;
  wire [31:0]\KR[2].key_reg[1][31]_1 ;
  wire \KR[3].key_host[0][0]_i_1_n_0 ;
  wire \KR[3].key_host[0][10]_i_1_n_0 ;
  wire \KR[3].key_host[0][11]_i_1_n_0 ;
  wire \KR[3].key_host[0][12]_i_1_n_0 ;
  wire \KR[3].key_host[0][13]_i_1_n_0 ;
  wire \KR[3].key_host[0][14]_i_1_n_0 ;
  wire \KR[3].key_host[0][15]_i_1_n_0 ;
  wire \KR[3].key_host[0][16]_i_1_n_0 ;
  wire \KR[3].key_host[0][17]_i_1_n_0 ;
  wire \KR[3].key_host[0][18]_i_1_n_0 ;
  wire \KR[3].key_host[0][19]_i_1_n_0 ;
  wire \KR[3].key_host[0][1]_i_1_n_0 ;
  wire \KR[3].key_host[0][20]_i_1_n_0 ;
  wire \KR[3].key_host[0][21]_i_1_n_0 ;
  wire \KR[3].key_host[0][22]_i_1_n_0 ;
  wire \KR[3].key_host[0][23]_i_1_n_0 ;
  wire \KR[3].key_host[0][24]_i_1_n_0 ;
  wire \KR[3].key_host[0][25]_i_1_n_0 ;
  wire \KR[3].key_host[0][26]_i_1_n_0 ;
  wire \KR[3].key_host[0][27]_i_1_n_0 ;
  wire \KR[3].key_host[0][28]_i_1_n_0 ;
  wire \KR[3].key_host[0][29]_i_1_n_0 ;
  wire \KR[3].key_host[0][2]_i_1_n_0 ;
  wire \KR[3].key_host[0][30]_i_1_n_0 ;
  wire \KR[3].key_host[0][31]_i_2_n_0 ;
  wire \KR[3].key_host[0][3]_i_1_n_0 ;
  wire \KR[3].key_host[0][4]_i_1_n_0 ;
  wire \KR[3].key_host[0][5]_i_1_n_0 ;
  wire \KR[3].key_host[0][6]_i_1_n_0 ;
  wire \KR[3].key_host[0][7]_i_1_n_0 ;
  wire \KR[3].key_host[0][8]_i_1_n_0 ;
  wire \KR[3].key_host[0][9]_i_1_n_0 ;
  wire [0:0]\KR[3].key_host_reg[0][0]_0 ;
  wire [31:0]\KR[3].key_host_reg[0]_3 ;
  wire [0:0]\KR[3].key_reg[0][31]_0 ;
  wire [6:0]O;
  wire [31:0]Q;
  wire SBOX_n_10;
  wire SBOX_n_11;
  wire SBOX_n_12;
  wire SBOX_n_13;
  wire SBOX_n_130;
  wire SBOX_n_131;
  wire SBOX_n_132;
  wire SBOX_n_137;
  wire SBOX_n_14;
  wire SBOX_n_141;
  wire SBOX_n_142;
  wire SBOX_n_143;
  wire SBOX_n_144;
  wire SBOX_n_145;
  wire SBOX_n_146;
  wire SBOX_n_147;
  wire SBOX_n_148;
  wire SBOX_n_15;
  wire SBOX_n_153;
  wire SBOX_n_156;
  wire SBOX_n_157;
  wire SBOX_n_158;
  wire SBOX_n_16;
  wire SBOX_n_17;
  wire SBOX_n_18;
  wire SBOX_n_19;
  wire SBOX_n_20;
  wire SBOX_n_21;
  wire SBOX_n_22;
  wire SBOX_n_23;
  wire SBOX_n_24;
  wire SBOX_n_25;
  wire SBOX_n_26;
  wire SBOX_n_27;
  wire SBOX_n_28;
  wire SBOX_n_29;
  wire SBOX_n_30;
  wire SBOX_n_31;
  wire SBOX_n_32;
  wire SBOX_n_33;
  wire SBOX_n_34;
  wire SBOX_n_35;
  wire SBOX_n_36;
  wire SBOX_n_37;
  wire SBOX_n_6;
  wire SBOX_n_63;
  wire SBOX_n_64;
  wire SBOX_n_65;
  wire SBOX_n_66;
  wire SBOX_n_67;
  wire SBOX_n_68;
  wire SBOX_n_69;
  wire SBOX_n_7;
  wire SBOX_n_70;
  wire SBOX_n_71;
  wire SBOX_n_72;
  wire SBOX_n_73;
  wire SBOX_n_74;
  wire SBOX_n_75;
  wire SBOX_n_76;
  wire SBOX_n_77;
  wire SBOX_n_78;
  wire SBOX_n_79;
  wire SBOX_n_8;
  wire SBOX_n_80;
  wire SBOX_n_81;
  wire SBOX_n_82;
  wire SBOX_n_83;
  wire SBOX_n_84;
  wire SBOX_n_85;
  wire SBOX_n_86;
  wire SBOX_n_87;
  wire SBOX_n_88;
  wire SBOX_n_89;
  wire SBOX_n_9;
  wire SBOX_n_90;
  wire SBOX_n_91;
  wire SBOX_n_92;
  wire SBOX_n_93;
  wire SBOX_n_94;
  wire [31:0]add_rd_key_in;
  wire [15:0]add_rk_out;
  wire add_rk_sel;
  wire \aes_cr_reg[0] ;
  wire [26:0]\aes_cr_reg[2] ;
  wire [2:0]\aes_cr_reg[2]_0 ;
  wire \base_new_pp_reg[3] ;
  wire \base_new_pp_reg[3]_0 ;
  wire \base_new_pp_reg[3]_1 ;
  wire \base_new_pp_reg[3]_2 ;
  wire \base_new_pp_reg[4] ;
  wire \base_new_pp_reg[4]_0 ;
  wire \base_new_pp_reg[4]_1 ;
  wire \base_new_pp_reg[4]_2 ;
  wire \base_new_pp_reg[4]_3 ;
  wire [31:0]bus_swap;
  wire bypass_key_en;
  wire clk_i;
  wire [3:0]col_en_cnt_unit_pp1;
  wire [0:0]\col_en_cnt_unit_pp1_reg[0]_0 ;
  wire [3:0]\col_en_cnt_unit_pp1_reg[3]_0 ;
  wire [3:0]\col_en_cnt_unit_pp2_reg[3]_0 ;
  wire [0:0]col_out;
  wire [1:0]col_sel_pp1;
  wire [1:0]\col_sel_pp1_reg[1]_0 ;
  wire [1:0]\col_sel_pp2_reg[1]_0 ;
  wire [10:0]data_in;
  wire [31:0]enable_i;
  wire \enable_i[0]_0 ;
  wire \enable_i[2]_0 ;
  wire \enable_i[3]_0 ;
  wire \enable_i[6]_0 ;
  wire \enable_i[6]_1 ;
  wire enable_i_0_sn_1;
  wire enable_i_10_sn_1;
  wire enable_i_11_sn_1;
  wire enable_i_12_sn_1;
  wire enable_i_13_sn_1;
  wire enable_i_14_sn_1;
  wire enable_i_15_sn_1;
  wire enable_i_16_sn_1;
  wire enable_i_17_sn_1;
  wire enable_i_18_sn_1;
  wire enable_i_19_sn_1;
  wire enable_i_1_sn_1;
  wire enable_i_20_sn_1;
  wire enable_i_21_sn_1;
  wire enable_i_22_sn_1;
  wire enable_i_23_sn_1;
  wire enable_i_24_sn_1;
  wire enable_i_25_sn_1;
  wire enable_i_26_sn_1;
  wire enable_i_27_sn_1;
  wire enable_i_28_sn_1;
  wire enable_i_29_sn_1;
  wire enable_i_2_sn_1;
  wire enable_i_30_sn_1;
  wire enable_i_31_sn_1;
  wire enable_i_3_sn_1;
  wire enable_i_4_sn_1;
  wire enable_i_5_sn_1;
  wire enable_i_6_sn_1;
  wire enable_i_7_sn_1;
  wire enable_i_8_sn_1;
  wire enable_i_9_sn_1;
  wire enc_dec_sbox;
  wire [1:0]g_func;
  wire \info_o[0] ;
  wire \info_o[0]_0 ;
  wire \info_o[0]_1 ;
  wire \info_o[0]_2 ;
  wire [1:0]\info_o[1] ;
  wire \info_o[28]_INST_0_i_7 ;
  wire \info_o[28]_INST_0_i_7_0 ;
  wire \info_o[31]_INST_0_i_13_n_0 ;
  wire isomorphism_inv_return033_out;
  wire isomorphism_inv_return033_out_3;
  wire isomorphism_inv_return033_out_9;
  wire isomorphism_inv_return03_out;
  wire isomorphism_inv_return03_out_1;
  wire isomorphism_inv_return03_out_7;
  wire isomorphism_inv_return05_out;
  wire isomorphism_inv_return05_out_10;
  wire isomorphism_inv_return05_out_4;
  wire isomorphism_return114_out;
  wire isomorphism_return114_out_13;
  wire isomorphism_return114_out_15;
  wire isomorphism_return114_out_17;
  wire isomorphism_return179_out;
  wire isomorphism_return179_out_12;
  wire isomorphism_return179_out_14;
  wire isomorphism_return179_out_16;
  wire [2:0]iv_en;
  wire iv_mux_out13_out;
  wire key_derivation_en;
  wire [2:0]key_en;
  wire [3:0]\key_en_pp1_reg[3]_0 ;
  wire [3:0]\key_en_pp1_reg[3]_1 ;
  wire [127:0]key_in;
  wire [21:0]key_out;
  wire [0:0]key_out_sel_pp1;
  wire [0:0]\key_out_sel_pp1_reg[1]_0 ;
  wire [0:0]key_out_sel_pp2;
  wire [0:0]\key_out_sel_pp2_reg[1]_0 ;
  wire key_sel;
  wire key_sel_mux;
  wire key_sel_pp1;
  wire [0:0]key_sel_rd;
  wire last_round;
  wire last_round_pp1;
  wire last_round_pp2;
  wire [15:0]last_round_pp2_reg_0;
  wire [31:0]mix_out_dec;
  wire p_16_in;
  wire p_16_in_0;
  wire p_16_in_6;
  wire p_86_in;
  wire p_86_in_11;
  wire p_86_in_5;
  wire p_93_in;
  wire p_93_in_2;
  wire p_93_in_8;
  wire rk_out_sel;
  wire rk_out_sel_pp1;
  wire rk_out_sel_pp2;
  wire [1:0]rk_sel_pp1;
  wire [1:0]\rk_sel_pp1_reg[1]_0 ;
  wire [1:0]rk_sel_pp2;
  wire [3:0]round_pp1;
  wire \round_pp1_reg[0]_0 ;
  wire \round_pp1_reg[0]_1 ;
  wire \round_pp1_reg[0]_2 ;
  wire \round_pp1_reg[3]_0 ;
  wire \round_pp1_reg[3]_1 ;
  wire \round_pp1_reg[3]_2 ;
  wire [3:0]\round_pp1_reg[3]_3 ;
  wire rst_i;
  wire [31:0]sbox_input;
  wire [5:0]sbox_out_enc;
  wire [31:0]sbox_pp2;
  wire \sbox_pp2[1]_i_3_n_0 ;
  wire \sbox_pp2[2]_i_3_n_0 ;
  wire \sbox_pp2[3]_i_2_n_0 ;
  wire \sbox_pp2[5]_i_3_n_0 ;
  wire \sbox_pp2_reg[31]_0 ;
  wire \sbox_pp2_reg[5]_0 ;
  wire [7:6]\NLW_IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_CO_UNCONNECTED ;
  wire [7:7]\NLW_IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_O_UNCONNECTED ;

  assign enable_i_0_sp_1 = enable_i_0_sn_1;
  assign enable_i_10_sp_1 = enable_i_10_sn_1;
  assign enable_i_11_sp_1 = enable_i_11_sn_1;
  assign enable_i_12_sp_1 = enable_i_12_sn_1;
  assign enable_i_13_sp_1 = enable_i_13_sn_1;
  assign enable_i_14_sp_1 = enable_i_14_sn_1;
  assign enable_i_15_sp_1 = enable_i_15_sn_1;
  assign enable_i_16_sp_1 = enable_i_16_sn_1;
  assign enable_i_17_sp_1 = enable_i_17_sn_1;
  assign enable_i_18_sp_1 = enable_i_18_sn_1;
  assign enable_i_19_sp_1 = enable_i_19_sn_1;
  assign enable_i_1_sp_1 = enable_i_1_sn_1;
  assign enable_i_20_sp_1 = enable_i_20_sn_1;
  assign enable_i_21_sp_1 = enable_i_21_sn_1;
  assign enable_i_22_sp_1 = enable_i_22_sn_1;
  assign enable_i_23_sp_1 = enable_i_23_sn_1;
  assign enable_i_24_sp_1 = enable_i_24_sn_1;
  assign enable_i_25_sp_1 = enable_i_25_sn_1;
  assign enable_i_26_sp_1 = enable_i_26_sn_1;
  assign enable_i_27_sp_1 = enable_i_27_sn_1;
  assign enable_i_28_sp_1 = enable_i_28_sn_1;
  assign enable_i_29_sp_1 = enable_i_29_sn_1;
  assign enable_i_2_sp_1 = enable_i_2_sn_1;
  assign enable_i_30_sp_1 = enable_i_30_sn_1;
  assign enable_i_31_sp_1 = enable_i_31_sn_1;
  assign enable_i_3_sp_1 = enable_i_3_sn_1;
  assign enable_i_4_sp_1 = enable_i_4_sn_1;
  assign enable_i_5_sp_1 = enable_i_5_sn_1;
  assign enable_i_6_sp_1 = enable_i_6_sn_1;
  assign enable_i_7_sp_1 = enable_i_7_sn_1;
  assign enable_i_8_sp_1 = enable_i_8_sn_1;
  assign enable_i_9_sp_1 = enable_i_9_sn_1;
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][0]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [0]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [0]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][0]_0 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][0]_i_12 
       (.I0(sbox_pp2[0]),
        .I1(\CD[0].col[3][0]_i_16_n_0 ),
        .I2(\CD[0].col[3][24]_i_17_n_0 ),
        .I3(\CD[0].col[3][12]_i_13_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][0]_i_15 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[7]),
        .I2(sbox_pp2[31]),
        .I3(sbox_pp2[24]),
        .I4(sbox_pp2[16]),
        .I5(sbox_pp2[8]),
        .O(\CD[0].col[3][0]_i_15_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CD[0].col[3][0]_i_16 
       (.I0(sbox_pp2[24]),
        .I1(sbox_pp2[16]),
        .I2(sbox_pp2[8]),
        .I3(sbox_pp2[22]),
        .I4(sbox_pp2[6]),
        .O(\CD[0].col[3][0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][0]_i_3 
       (.I0(key_out[0]),
        .I1(add_rd_key_in[0]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[0]),
        .I5(sbox_pp2[0]),
        .O(add_rk_out[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][0]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [0]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [0]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][0]_i_6 
       (.I0(bus_swap[0]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][0]_i_12_n_0 ),
        .I3(add_rd_key_in[0]),
        .I4(key_out[0]),
        .I5(add_rk_sel),
        .O(enable_i_16_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][0]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][0]_0 ),
        .I2(\CD[0].col[3][0]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[0]),
        .I5(\CD[0].col[3][0]_i_15_n_0 ),
        .O(add_rd_key_in[0]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][0]_i_9 
       (.I0(\CD[0].col[3][30]_i_17_n_0 ),
        .I1(sbox_pp2[8]),
        .I2(\CD[0].col[3][8]_i_11_n_0 ),
        .I3(\CD[0].col[3][24]_i_17_n_0 ),
        .I4(sbox_pp2[7]),
        .I5(sbox_pp2[31]),
        .O(mix_out_dec[0]));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][10]_i_11 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[26]),
        .I2(sbox_pp2[2]),
        .I3(sbox_pp2[9]),
        .I4(sbox_pp2[18]),
        .I5(sbox_pp2[1]),
        .O(\CD[0].col[3][10]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][10]_i_13 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [6]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][10]_0 ));
  LUT6 #(
    .INIT(64'h0000AAA00000CCC0)) 
    \CD[0].col[3][10]_i_14 
       (.I0(sbox_pp2[10]),
        .I1(mix_out_dec[10]),
        .I2(\CD[0].col[3][9]_i_8_1 [0]),
        .I3(\CD[0].col[3][9]_i_8_1 [1]),
        .I4(rk_out_sel_pp2),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][10]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][10]_i_2 
       (.I0(\KR[1].key_reg[2][10]_0 ),
        .I1(add_rd_key_in[10]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[10]),
        .I5(sbox_pp2[10]),
        .O(last_round_pp2_reg_0[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][10]_i_4 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_147),
        .I2(\CD[0].col[3][10]_i_8_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[10]),
        .I5(\CD[0].col[3][10]_i_11_n_0 ),
        .O(add_rd_key_in[10]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][10]_i_5 
       (.I0(sbox_pp2[18]),
        .I1(sbox_pp2[24]),
        .I2(\CD[0].col[3][29]_i_17_n_0 ),
        .I3(sbox_pp2[9]),
        .I4(sbox_pp2[1]),
        .I5(sbox_pp2[8]),
        .O(mix_out_dec[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][10]_i_7 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [10]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [10]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][10]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][10]_i_8 
       (.I0(bus_swap[10]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][10]_i_14_n_0 ),
        .I3(add_rd_key_in[10]),
        .I4(\KR[1].key_reg[2][10]_0 ),
        .I5(add_rk_sel),
        .O(enable_i_26_sn_1));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][11]_i_10 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(\CD[0].col[3][11]_i_16_n_0 ),
        .I2(sbox_pp2[10]),
        .I3(\CD[0].col[3][27]_i_20_n_0 ),
        .I4(sbox_pp2[2]),
        .I5(sbox_pp2[3]),
        .O(\CD[0].col[3][11]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CD[0].col[3][11]_i_11 
       (.I0(sbox_pp2[27]),
        .I1(sbox_pp2[19]),
        .I2(sbox_pp2[10]),
        .O(\CD[0].col[3][11]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][11]_i_12 
       (.I0(sbox_pp2[31]),
        .I1(sbox_pp2[23]),
        .O(\CD[0].col[3][11]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair270" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][11]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [7]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][11]_0 ));
  LUT5 #(
    .INIT(32'h00AA003C)) 
    \CD[0].col[3][11]_i_15 
       (.I0(sbox_pp2[11]),
        .I1(\CD[0].col[3][27]_i_16_n_0 ),
        .I2(\CD[0].col[3][11]_i_17_n_0 ),
        .I3(add_rk_sel),
        .I4(last_round_pp2),
        .O(\CD[0].col[3][11]_i_15_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair272" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][11]_i_16 
       (.I0(sbox_pp2[19]),
        .I1(sbox_pp2[27]),
        .O(\CD[0].col[3][11]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][11]_i_17 
       (.I0(\CD[0].col[3][11]_i_12_n_0 ),
        .I1(\CD[0].col[3][27]_i_19_n_0 ),
        .I2(sbox_pp2[3]),
        .I3(sbox_pp2[2]),
        .I4(\CD[0].col[3][11]_i_16_n_0 ),
        .I5(sbox_pp2[10]),
        .O(\CD[0].col[3][11]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][11]_i_2 
       (.I0(\KR[1].key_reg[2][11]_0 ),
        .I1(add_rd_key_in[11]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[11]),
        .I5(sbox_pp2[11]),
        .O(last_round_pp2_reg_0[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][11]_i_4 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_145),
        .I2(\base_new_pp_reg[3]_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[11]),
        .I5(\CD[0].col[3][11]_i_10_n_0 ),
        .O(add_rd_key_in[11]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][11]_i_5 
       (.I0(\CD[0].col[3][27]_i_16_n_0 ),
        .I1(\CD[0].col[3][11]_i_11_n_0 ),
        .I2(sbox_pp2[2]),
        .I3(sbox_pp2[3]),
        .I4(\CD[0].col[3][27]_i_19_n_0 ),
        .I5(\CD[0].col[3][11]_i_12_n_0 ),
        .O(mix_out_dec[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][11]_i_7 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [11]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [11]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][11]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][11]_i_8 
       (.I0(bus_swap[11]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][11]_i_15_n_0 ),
        .I3(add_rd_key_in[11]),
        .I4(\KR[1].key_reg[2][11]_0 ),
        .I5(add_rk_sel),
        .O(enable_i_27_sn_1));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][12]_i_11 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(\CD[0].col[3][27]_i_20_n_0 ),
        .I2(sbox_pp2[11]),
        .I3(sbox_pp2[3]),
        .I4(\CD[0].col[3][29]_i_18_n_0 ),
        .I5(sbox_pp2[4]),
        .O(\CD[0].col[3][12]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CD[0].col[3][12]_i_12 
       (.I0(sbox_pp2[4]),
        .I1(sbox_pp2[9]),
        .I2(sbox_pp2[25]),
        .I3(sbox_pp2[26]),
        .I4(sbox_pp2[10]),
        .O(\CD[0].col[3][12]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair275" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][12]_i_13 
       (.I0(sbox_pp2[7]),
        .I1(sbox_pp2[31]),
        .O(\CD[0].col[3][12]_i_13_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair271" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][12]_i_15 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [8]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][12]_0 ));
  LUT5 #(
    .INIT(32'h00AA003C)) 
    \CD[0].col[3][12]_i_16 
       (.I0(sbox_pp2[12]),
        .I1(\CD[0].col[3][28]_i_15_n_0 ),
        .I2(\CD[0].col[3][12]_i_18_n_0 ),
        .I3(add_rk_sel),
        .I4(last_round_pp2),
        .O(\CD[0].col[3][12]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][12]_i_18 
       (.I0(\CD[0].col[3][29]_i_18_n_0 ),
        .I1(\CD[0].col[3][12]_i_19_n_0 ),
        .I2(sbox_pp2[10]),
        .I3(sbox_pp2[26]),
        .I4(\CD[0].col[3][1]_i_17_n_0 ),
        .I5(sbox_pp2[4]),
        .O(\CD[0].col[3][12]_i_18_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CD[0].col[3][12]_i_19 
       (.I0(sbox_pp2[11]),
        .I1(sbox_pp2[3]),
        .I2(sbox_pp2[31]),
        .I3(sbox_pp2[7]),
        .O(\CD[0].col[3][12]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][12]_i_2 
       (.I0(\KR[1].key_reg[2][12]_0 ),
        .I1(add_rd_key_in[12]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[12]),
        .I5(sbox_pp2[12]),
        .O(last_round_pp2_reg_0[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][12]_i_4 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_143),
        .I2(\CD[0].col[3][12]_i_8_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[12]),
        .I5(\CD[0].col[3][12]_i_11_n_0 ),
        .O(add_rd_key_in[12]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][12]_i_5 
       (.I0(\CD[0].col[3][28]_i_15_n_0 ),
        .I1(\CD[0].col[3][12]_i_12_n_0 ),
        .I2(\CD[0].col[3][12]_i_13_n_0 ),
        .I3(sbox_pp2[3]),
        .I4(sbox_pp2[11]),
        .I5(\CD[0].col[3][29]_i_18_n_0 ),
        .O(mix_out_dec[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][12]_i_7 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [12]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [12]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][12]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][12]_i_8 
       (.I0(bus_swap[12]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][12]_i_16_n_0 ),
        .I3(add_rd_key_in[12]),
        .I4(\KR[1].key_reg[2][12]_0 ),
        .I5(add_rk_sel),
        .O(enable_i_28_sn_1));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][13]_i_10 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[4]),
        .I2(sbox_pp2[12]),
        .I3(sbox_pp2[29]),
        .I4(sbox_pp2[21]),
        .I5(sbox_pp2[5]),
        .O(\CD[0].col[3][13]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair271" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][13]_i_12 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [9]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][13]_0 ));
  LUT6 #(
    .INIT(64'h0000AAA00000CCC0)) 
    \CD[0].col[3][13]_i_13 
       (.I0(sbox_pp2[13]),
        .I1(mix_out_dec[13]),
        .I2(\CD[0].col[3][9]_i_8_1 [0]),
        .I3(\CD[0].col[3][9]_i_8_1 [1]),
        .I4(rk_out_sel_pp2),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][13]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][13]_i_2 
       (.I0(key_out[3]),
        .I1(add_rd_key_in[13]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[13]),
        .I5(sbox_pp2[13]),
        .O(last_round_pp2_reg_0[5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][13]_i_4 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][13]_0 ),
        .I2(\CD[0].col[3][13]_i_8_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[13]),
        .I5(\CD[0].col[3][13]_i_10_n_0 ),
        .O(add_rd_key_in[13]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][13]_i_5 
       (.I0(\CD[0].col[3][30]_i_16_n_0 ),
        .I1(sbox_pp2[5]),
        .I2(\CD[0].col[3][29]_i_17_n_0 ),
        .I3(\CD[0].col[3][29]_i_16_n_0 ),
        .I4(\CD[0].col[3][28]_i_16_n_0 ),
        .I5(sbox_pp2[11]),
        .O(mix_out_dec[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][13]_i_7 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [13]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [13]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][13]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][13]_i_8 
       (.I0(bus_swap[13]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][13]_i_13_n_0 ),
        .I3(add_rd_key_in[13]),
        .I4(key_out[3]),
        .I5(add_rk_sel),
        .O(enable_i_29_sn_1));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][14]_i_10 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[5]),
        .I2(sbox_pp2[13]),
        .I3(sbox_pp2[6]),
        .I4(sbox_pp2[22]),
        .I5(sbox_pp2[30]),
        .O(\CD[0].col[3][14]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][14]_i_12 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [10]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [14]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][14]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][14]_i_13 
       (.I0(sbox_pp2[14]),
        .I1(\CD[0].col[3][30]_i_17_n_0 ),
        .I2(\CD[0].col[3][30]_i_18_n_0 ),
        .I3(\CD[0].col[3][14]_i_16_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][14]_i_13_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][14]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [10]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][14]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CD[0].col[3][14]_i_16 
       (.I0(sbox_pp2[30]),
        .I1(sbox_pp2[5]),
        .I2(sbox_pp2[13]),
        .I3(sbox_pp2[28]),
        .I4(sbox_pp2[12]),
        .O(\CD[0].col[3][14]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][14]_i_2 
       (.I0(key_out[4]),
        .I1(add_rd_key_in[14]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[14]),
        .I5(sbox_pp2[14]),
        .O(last_round_pp2_reg_0[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][14]_i_4 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][14]_0 ),
        .I2(\base_new_pp_reg[4]_1 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[14]),
        .I5(\CD[0].col[3][14]_i_10_n_0 ),
        .O(add_rd_key_in[14]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][14]_i_5 
       (.I0(\CD[0].col[3][30]_i_17_n_0 ),
        .I1(\CD[0].col[3][30]_i_18_n_0 ),
        .I2(sbox_pp2[12]),
        .I3(sbox_pp2[28]),
        .I4(\CD[0].col[3][29]_i_19_n_0 ),
        .I5(sbox_pp2[30]),
        .O(mix_out_dec[14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][14]_i_7 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [14]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [14]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][14]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][14]_i_8 
       (.I0(bus_swap[14]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][14]_i_13_n_0 ),
        .I3(add_rd_key_in[14]),
        .I4(key_out[4]),
        .I5(add_rk_sel),
        .O(enable_i_30_sn_1));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][15]_i_10 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [15]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [15]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][15]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][15]_i_11 
       (.I0(bus_swap[15]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][15]_i_18_n_0 ),
        .I3(add_rd_key_in[15]),
        .I4(key_out[5]),
        .I5(add_rk_sel),
        .O(enable_i_31_sn_1));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][15]_i_14 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[23]),
        .I2(sbox_pp2[7]),
        .I3(sbox_pp2[31]),
        .I4(sbox_pp2[6]),
        .I5(sbox_pp2[14]),
        .O(\CD[0].col[3][15]_i_14_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CD[0].col[3][15]_i_15 
       (.I0(sbox_pp2[31]),
        .I1(sbox_pp2[7]),
        .I2(sbox_pp2[14]),
        .O(\CD[0].col[3][15]_i_15_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][15]_i_17 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [11]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [15]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][15]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][15]_i_18 
       (.I0(sbox_pp2[15]),
        .I1(\CD[0].col[3][28]_i_16_n_0 ),
        .I2(\CD[0].col[3][29]_i_18_n_0 ),
        .I3(\CD[0].col[3][15]_i_22_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][15]_i_18_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][15]_i_19 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [11]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][15]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][15]_i_22 
       (.I0(sbox_pp2[14]),
        .I1(\CD[0].col[3][12]_i_13_n_0 ),
        .I2(sbox_pp2[13]),
        .I3(sbox_pp2[29]),
        .I4(sbox_pp2[23]),
        .I5(sbox_pp2[6]),
        .O(\CD[0].col[3][15]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][15]_i_4 
       (.I0(key_out[5]),
        .I1(add_rd_key_in[15]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[15]),
        .I5(sbox_pp2[15]),
        .O(last_round_pp2_reg_0[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][15]_i_7 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_131),
        .I2(\CD[0].col[3][15]_i_11_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[15]),
        .I5(\CD[0].col[3][15]_i_14_n_0 ),
        .O(add_rd_key_in[15]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][15]_i_8 
       (.I0(\CD[0].col[3][31]_i_33_n_0 ),
        .I1(sbox_pp2[6]),
        .I2(sbox_pp2[23]),
        .I3(sbox_pp2[29]),
        .I4(sbox_pp2[13]),
        .I5(\CD[0].col[3][15]_i_15_n_0 ),
        .O(mix_out_dec[15]));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][16]_i_10 
       (.I0(sbox_pp2[16]),
        .I1(\CD[0].col[3][16]_i_13_n_0 ),
        .I2(\CD[0].col[3][24]_i_17_n_0 ),
        .I3(\CD[0].col[3][31]_i_35_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][16]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][16]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [12]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][16]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CD[0].col[3][16]_i_13 
       (.I0(sbox_pp2[8]),
        .I1(sbox_pp2[0]),
        .I2(sbox_pp2[24]),
        .I3(sbox_pp2[22]),
        .I4(sbox_pp2[6]),
        .O(\CD[0].col[3][16]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][16]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [16]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [16]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][16]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][16]_i_6 
       (.I0(bus_swap[16]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][16]_i_10_n_0 ),
        .I3(add_rd_key_in[16]),
        .I4(key_out[6]),
        .I5(add_rk_sel),
        .O(\enable_i[0]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][16]_i_9 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [12]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [16]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][16]_1 ));
  LUT6 #(
    .INIT(64'h0000AAA00000CCC0)) 
    \CD[0].col[3][17]_i_10 
       (.I0(sbox_pp2[17]),
        .I1(mix_out_dec[17]),
        .I2(\CD[0].col[3][9]_i_8_1 [0]),
        .I3(\CD[0].col[3][9]_i_8_1 [1]),
        .I4(rk_out_sel_pp2),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][17]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][17]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [13]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][17]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][17]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [17]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [17]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][17]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][17]_i_6 
       (.I0(bus_swap[17]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][17]_i_10_n_0 ),
        .I3(add_rd_key_in[17]),
        .I4(key_out[7]),
        .I5(add_rk_sel),
        .O(enable_i_1_sn_1));
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][17]_i_9 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [13]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [17]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][17]_1 ));
  LUT6 #(
    .INIT(64'h0000AAA00000CCC0)) 
    \CD[0].col[3][18]_i_10 
       (.I0(sbox_pp2[18]),
        .I1(mix_out_dec[18]),
        .I2(\CD[0].col[3][9]_i_8_1 [0]),
        .I3(\CD[0].col[3][9]_i_8_1 [1]),
        .I4(rk_out_sel_pp2),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][18]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][18]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [14]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][18]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][18]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [18]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [18]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][18]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][18]_i_6 
       (.I0(bus_swap[18]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][18]_i_10_n_0 ),
        .I3(add_rd_key_in[18]),
        .I4(key_out[8]),
        .I5(add_rk_sel),
        .O(\enable_i[2]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][18]_i_9 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [14]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [18]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][18]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][19]_i_10 
       (.I0(sbox_pp2[19]),
        .I1(\CD[0].col[3][19]_i_13_n_0 ),
        .I2(\CD[0].col[3][27]_i_19_n_0 ),
        .I3(\CD[0].col[3][29]_i_16_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][19]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][19]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [15]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][19]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CD[0].col[3][19]_i_13 
       (.I0(\CD[0].col[3][28]_i_15_n_0 ),
        .I1(sbox_pp2[7]),
        .I2(sbox_pp2[31]),
        .I3(sbox_pp2[3]),
        .I4(sbox_pp2[11]),
        .O(\CD[0].col[3][19]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][19]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [19]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [19]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][19]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][19]_i_6 
       (.I0(bus_swap[19]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][19]_i_10_n_0 ),
        .I3(add_rd_key_in[19]),
        .I4(key_out[9]),
        .I5(add_rk_sel),
        .O(\enable_i[3]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][19]_i_9 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [15]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [19]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][19]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][1]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3]_4 [1]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [1]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][1]_1 ));
  LUT6 #(
    .INIT(64'h0000AAA00000CCC0)) 
    \CD[0].col[3][1]_i_13 
       (.I0(sbox_pp2[1]),
        .I1(mix_out_dec[1]),
        .I2(\CD[0].col[3][9]_i_8_1 [0]),
        .I3(\CD[0].col[3][9]_i_8_1 [1]),
        .I4(rk_out_sel_pp2),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][1]_i_13_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][1]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3]_4 [1]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][1]_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][1]_i_16 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[17]),
        .I2(sbox_pp2[0]),
        .I3(\CD[0].col[3][1]_i_17_n_0 ),
        .I4(\CD[0].col[3][12]_i_13_n_0 ),
        .I5(sbox_pp2[24]),
        .O(\CD[0].col[3][1]_i_16_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][1]_i_17 
       (.I0(sbox_pp2[9]),
        .I1(sbox_pp2[25]),
        .O(\CD[0].col[3][1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][1]_i_3 
       (.I0(\sbox_pp2[1]_i_3_n_0 ),
        .I1(add_rd_key_in[1]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[1]),
        .I5(sbox_pp2[1]),
        .O(add_rk_out[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][1]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [1]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [1]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][1]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][1]_i_6 
       (.I0(bus_swap[1]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][1]_i_13_n_0 ),
        .I3(add_rd_key_in[1]),
        .I4(\sbox_pp2[1]_i_3_n_0 ),
        .I5(add_rk_sel),
        .O(enable_i_17_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][1]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][1]_0 ),
        .I2(\CD[0].col[3][1]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[1]),
        .I5(\CD[0].col[3][1]_i_16_n_0 ),
        .O(add_rd_key_in[1]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][1]_i_9 
       (.I0(sbox_pp2[24]),
        .I1(sbox_pp2[31]),
        .I2(sbox_pp2[23]),
        .I3(\CD[0].col[3][27]_i_16_n_0 ),
        .I4(sbox_pp2[0]),
        .I5(sbox_pp2[17]),
        .O(mix_out_dec[1]));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][20]_i_10 
       (.I0(sbox_pp2[20]),
        .I1(sbox_pp2[11]),
        .I2(\CD[0].col[3][28]_i_16_n_0 ),
        .I3(\CD[0].col[3][20]_i_13_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][20]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][20]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [16]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][20]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][20]_i_13 
       (.I0(\CD[1].col[2][20]_i_8_n_0 ),
        .I1(\CD[0].col[3][27]_i_17_n_0 ),
        .I2(sbox_pp2[28]),
        .I3(sbox_pp2[2]),
        .I4(\CD[0].col[3][4]_i_19_n_0 ),
        .I5(\CD[0].col[3][27]_i_20_n_0 ),
        .O(\CD[0].col[3][20]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][20]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [20]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [20]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][20]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][20]_i_6 
       (.I0(bus_swap[20]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][20]_i_10_n_0 ),
        .I3(add_rd_key_in[20]),
        .I4(key_out[10]),
        .I5(add_rk_sel),
        .O(enable_i_4_sn_1));
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][20]_i_9 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [16]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [20]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][20]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][21]_i_10 
       (.I0(sbox_pp2[21]),
        .I1(\CD[1].col[2][21]_i_6_n_0 ),
        .I2(\CD[0].col[3][5]_i_18_n_0 ),
        .I3(\CD[0].col[3][21]_i_13_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][21]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][21]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [17]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][21]_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][21]_i_13 
       (.I0(sbox_pp2[10]),
        .I1(sbox_pp2[18]),
        .I2(sbox_pp2[3]),
        .I3(sbox_pp2[12]),
        .I4(sbox_pp2[19]),
        .I5(\CD[0].col[3][29]_i_19_n_0 ),
        .O(\CD[0].col[3][21]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][21]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [21]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [21]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][21]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][21]_i_6 
       (.I0(bus_swap[21]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][21]_i_10_n_0 ),
        .I3(add_rd_key_in[21]),
        .I4(key_out[11]),
        .I5(add_rk_sel),
        .O(enable_i_5_sn_1));
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][21]_i_9 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [17]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [21]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][21]_1 ));
  LUT6 #(
    .INIT(64'h0000AAA00000CCC0)) 
    \CD[0].col[3][22]_i_10 
       (.I0(sbox_pp2[22]),
        .I1(mix_out_dec[22]),
        .I2(\CD[0].col[3][9]_i_8_1 [0]),
        .I3(\CD[0].col[3][9]_i_8_1 [1]),
        .I4(rk_out_sel_pp2),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][22]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][22]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [18]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][22]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][22]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [22]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [22]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][22]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][22]_i_6 
       (.I0(bus_swap[22]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][22]_i_10_n_0 ),
        .I3(add_rd_key_in[22]),
        .I4(key_out[12]),
        .I5(add_rk_sel),
        .O(\enable_i[6]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][22]_i_9 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [18]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [22]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][22]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][23]_i_10 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [19]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [23]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][23]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][23]_i_11 
       (.I0(sbox_pp2[23]),
        .I1(\CD[0].col[3][31]_i_33_n_0 ),
        .I2(\CD[0].col[3][6]_i_16_n_0 ),
        .I3(\CD[0].col[3][23]_i_14_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][23]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][23]_i_12 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [19]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][23]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CD[0].col[3][23]_i_14 
       (.I0(sbox_pp2[14]),
        .I1(sbox_pp2[7]),
        .I2(sbox_pp2[31]),
        .I3(sbox_pp2[21]),
        .I4(sbox_pp2[15]),
        .O(\CD[0].col[3][23]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][23]_i_6 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [23]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [23]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][23]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][23]_i_7 
       (.I0(bus_swap[23]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][23]_i_11_n_0 ),
        .I3(add_rd_key_in[23]),
        .I4(key_out[13]),
        .I5(add_rk_sel),
        .O(enable_i_7_sn_1));
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][24]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [20]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [24]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][24]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][24]_i_12 
       (.I0(sbox_pp2[24]),
        .I1(\CD[0].col[3][24]_i_19_n_0 ),
        .I2(\CD[0].col[3][24]_i_17_n_0 ),
        .I3(\CD[0].col[3][24]_i_18_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][24]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][24]_i_13 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [20]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][24]_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][24]_i_15 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[0]),
        .I2(sbox_pp2[8]),
        .I3(sbox_pp2[23]),
        .I4(sbox_pp2[31]),
        .I5(sbox_pp2[16]),
        .O(\CD[0].col[3][24]_i_15_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][24]_i_16 
       (.I0(sbox_pp2[30]),
        .I1(sbox_pp2[14]),
        .O(\CD[0].col[3][24]_i_16_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CD[0].col[3][24]_i_17 
       (.I0(sbox_pp2[29]),
        .I1(sbox_pp2[21]),
        .I2(sbox_pp2[13]),
        .I3(sbox_pp2[5]),
        .O(\CD[0].col[3][24]_i_17_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][24]_i_18 
       (.I0(sbox_pp2[0]),
        .I1(sbox_pp2[8]),
        .O(\CD[0].col[3][24]_i_18_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CD[0].col[3][24]_i_19 
       (.I0(sbox_pp2[23]),
        .I1(sbox_pp2[31]),
        .I2(sbox_pp2[16]),
        .I3(sbox_pp2[30]),
        .I4(sbox_pp2[14]),
        .O(\CD[0].col[3][24]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][24]_i_3 
       (.I0(key_out[14]),
        .I1(add_rd_key_in[24]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[24]),
        .I5(sbox_pp2[24]),
        .O(last_round_pp2_reg_0[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][24]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [24]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [24]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][24]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][24]_i_6 
       (.I0(bus_swap[24]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][24]_i_12_n_0 ),
        .I3(add_rd_key_in[24]),
        .I4(key_out[14]),
        .I5(add_rk_sel),
        .O(enable_i_8_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][24]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][24]_0 ),
        .I2(\CD[0].col[3][24]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[24]),
        .I5(\CD[0].col[3][24]_i_15_n_0 ),
        .O(add_rd_key_in[24]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][24]_i_9 
       (.I0(\CD[0].col[3][24]_i_16_n_0 ),
        .I1(sbox_pp2[16]),
        .I2(sbox_pp2[31]),
        .I3(sbox_pp2[23]),
        .I4(\CD[0].col[3][24]_i_17_n_0 ),
        .I5(\CD[0].col[3][24]_i_18_n_0 ),
        .O(mix_out_dec[24]));
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][25]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [21]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [25]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][25]_1 ));
  LUT6 #(
    .INIT(64'h0000AAA00000CCC0)) 
    \CD[0].col[3][25]_i_12 
       (.I0(sbox_pp2[25]),
        .I1(mix_out_dec[25]),
        .I2(\CD[0].col[3][9]_i_8_1 [0]),
        .I3(\CD[0].col[3][9]_i_8_1 [1]),
        .I4(rk_out_sel_pp2),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][25]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][25]_i_13 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [21]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][25]_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][25]_i_15 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(\CD[0].col[3][11]_i_12_n_0 ),
        .I2(\CD[0].col[3][8]_i_11_n_0 ),
        .I3(sbox_pp2[17]),
        .I4(sbox_pp2[1]),
        .I5(sbox_pp2[9]),
        .O(\CD[0].col[3][25]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][25]_i_3 
       (.I0(key_out[15]),
        .I1(add_rd_key_in[25]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[25]),
        .I5(sbox_pp2[25]),
        .O(last_round_pp2_reg_0[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][25]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [25]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [25]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][25]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][25]_i_6 
       (.I0(bus_swap[25]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][25]_i_12_n_0 ),
        .I3(add_rd_key_in[25]),
        .I4(key_out[15]),
        .I5(add_rk_sel),
        .O(enable_i_9_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][25]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][25]_0 ),
        .I2(\CD[0].col[3][25]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[25]),
        .I5(\CD[0].col[3][25]_i_15_n_0 ),
        .O(add_rd_key_in[25]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][25]_i_9 
       (.I0(sbox_pp2[9]),
        .I1(sbox_pp2[15]),
        .I2(sbox_pp2[23]),
        .I3(sbox_pp2[16]),
        .I4(sbox_pp2[24]),
        .I5(\CD[0].col[3][28]_i_15_n_0 ),
        .O(mix_out_dec[25]));
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][26]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [22]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [26]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][26]_1 ));
  LUT5 #(
    .INIT(32'h00AA003C)) 
    \CD[0].col[3][26]_i_12 
       (.I0(sbox_pp2[26]),
        .I1(\CD[0].col[3][26]_i_17_n_0 ),
        .I2(\CD[0].col[3][26]_i_19_n_0 ),
        .I3(add_rk_sel),
        .I4(last_round_pp2),
        .O(\CD[0].col[3][26]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][26]_i_13 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [22]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][26]_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][26]_i_16 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[18]),
        .I2(sbox_pp2[10]),
        .I3(sbox_pp2[25]),
        .I4(sbox_pp2[2]),
        .I5(sbox_pp2[17]),
        .O(\CD[0].col[3][26]_i_16_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair269" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CD[0].col[3][26]_i_17 
       (.I0(sbox_pp2[18]),
        .I1(sbox_pp2[10]),
        .I2(sbox_pp2[25]),
        .O(\CD[0].col[3][26]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][26]_i_18 
       (.I0(sbox_pp2[23]),
        .I1(sbox_pp2[7]),
        .I2(sbox_pp2[30]),
        .I3(sbox_pp2[14]),
        .I4(sbox_pp2[22]),
        .I5(sbox_pp2[6]),
        .O(\CD[0].col[3][26]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][26]_i_19 
       (.I0(\CD[0].col[3][26]_i_21_n_0 ),
        .I1(\CD[0].col[3][26]_i_22_n_0 ),
        .I2(sbox_pp2[2]),
        .I3(sbox_pp2[24]),
        .I4(sbox_pp2[8]),
        .I5(sbox_pp2[17]),
        .O(\CD[0].col[3][26]_i_19_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CD[0].col[3][26]_i_21 
       (.I0(sbox_pp2[6]),
        .I1(sbox_pp2[22]),
        .I2(sbox_pp2[14]),
        .I3(sbox_pp2[30]),
        .O(\CD[0].col[3][26]_i_21_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair275" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][26]_i_22 
       (.I0(sbox_pp2[7]),
        .I1(sbox_pp2[23]),
        .O(\CD[0].col[3][26]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][26]_i_3 
       (.I0(key_out[16]),
        .I1(add_rd_key_in[26]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[26]),
        .I5(sbox_pp2[26]),
        .O(last_round_pp2_reg_0[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][26]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [26]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [26]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][26]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][26]_i_6 
       (.I0(bus_swap[26]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][26]_i_12_n_0 ),
        .I3(add_rd_key_in[26]),
        .I4(key_out[16]),
        .I5(add_rk_sel),
        .O(enable_i_10_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][26]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_148),
        .I2(\CD[0].col[3][26]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[26]),
        .I5(\CD[0].col[3][26]_i_16_n_0 ),
        .O(add_rd_key_in[26]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][26]_i_9 
       (.I0(\CD[0].col[3][26]_i_17_n_0 ),
        .I1(sbox_pp2[17]),
        .I2(sbox_pp2[8]),
        .I3(sbox_pp2[24]),
        .I4(sbox_pp2[2]),
        .I5(\CD[0].col[3][26]_i_18_n_0 ),
        .O(mix_out_dec[26]));
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][27]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [23]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [27]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][27]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][27]_i_12 
       (.I0(sbox_pp2[27]),
        .I1(\CD[0].col[3][27]_i_16_n_0 ),
        .I2(\CD[0].col[3][27]_i_17_n_0 ),
        .I3(\CD[0].col[3][27]_i_21_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][27]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][27]_i_13 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [23]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][27]_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][27]_i_15 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[19]),
        .I2(sbox_pp2[18]),
        .I3(\CD[0].col[3][11]_i_12_n_0 ),
        .I4(\CD[0].col[3][27]_i_18_n_0 ),
        .I5(sbox_pp2[26]),
        .O(\CD[0].col[3][27]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][27]_i_16 
       (.I0(\CD[0].col[3][24]_i_16_n_0 ),
        .I1(sbox_pp2[9]),
        .I2(sbox_pp2[25]),
        .I3(\CD[0].col[3][29]_i_19_n_0 ),
        .I4(sbox_pp2[21]),
        .I5(sbox_pp2[29]),
        .O(\CD[0].col[3][27]_i_16_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair272" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][27]_i_17 
       (.I0(sbox_pp2[18]),
        .I1(sbox_pp2[19]),
        .O(\CD[0].col[3][27]_i_17_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair273" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][27]_i_18 
       (.I0(sbox_pp2[3]),
        .I1(sbox_pp2[11]),
        .O(\CD[0].col[3][27]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \CD[0].col[3][27]_i_19 
       (.I0(sbox_pp2[24]),
        .I1(sbox_pp2[16]),
        .I2(sbox_pp2[8]),
        .I3(sbox_pp2[0]),
        .O(\CD[0].col[3][27]_i_19_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][27]_i_20 
       (.I0(sbox_pp2[7]),
        .I1(sbox_pp2[15]),
        .O(\CD[0].col[3][27]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][27]_i_21 
       (.I0(\CD[0].col[3][27]_i_20_n_0 ),
        .I1(\CD[0].col[3][8]_i_11_n_0 ),
        .I2(\CD[0].col[3][24]_i_18_n_0 ),
        .I3(sbox_pp2[26]),
        .I4(sbox_pp2[3]),
        .I5(sbox_pp2[11]),
        .O(\CD[0].col[3][27]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][27]_i_3 
       (.I0(key_out[17]),
        .I1(add_rd_key_in[27]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[27]),
        .I5(sbox_pp2[27]),
        .O(last_round_pp2_reg_0[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][27]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [27]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [27]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][27]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][27]_i_6 
       (.I0(bus_swap[27]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][27]_i_12_n_0 ),
        .I3(add_rd_key_in[27]),
        .I4(key_out[17]),
        .I5(add_rk_sel),
        .O(enable_i_11_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][27]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_146),
        .I2(\base_new_pp_reg[3]_1 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[27]),
        .I5(\CD[0].col[3][27]_i_15_n_0 ),
        .O(add_rd_key_in[27]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][27]_i_9 
       (.I0(\CD[0].col[3][27]_i_16_n_0 ),
        .I1(\CD[0].col[3][27]_i_17_n_0 ),
        .I2(\CD[0].col[3][27]_i_18_n_0 ),
        .I3(sbox_pp2[26]),
        .I4(\CD[0].col[3][27]_i_19_n_0 ),
        .I5(\CD[0].col[3][27]_i_20_n_0 ),
        .O(mix_out_dec[27]));
  (* SOFT_HLUTNM = "soft_lutpair270" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][28]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [24]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][28]_0 ));
  LUT5 #(
    .INIT(32'h00AA003C)) 
    \CD[0].col[3][28]_i_12 
       (.I0(sbox_pp2[28]),
        .I1(\CD[0].col[3][28]_i_15_n_0 ),
        .I2(\CD[0].col[3][28]_i_19_n_0 ),
        .I3(add_rk_sel),
        .I4(last_round_pp2),
        .O(\CD[0].col[3][28]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][28]_i_14 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(\CD[0].col[3][11]_i_12_n_0 ),
        .I2(sbox_pp2[27]),
        .I3(sbox_pp2[19]),
        .I4(\CD[0].col[3][28]_i_16_n_0 ),
        .I5(sbox_pp2[20]),
        .O(\CD[0].col[3][28]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][28]_i_15 
       (.I0(sbox_pp2[29]),
        .I1(sbox_pp2[21]),
        .I2(\CD[0].col[3][29]_i_19_n_0 ),
        .I3(sbox_pp2[1]),
        .I4(sbox_pp2[17]),
        .I5(\CD[0].col[3][30]_i_17_n_0 ),
        .O(\CD[0].col[3][28]_i_15_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair274" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][28]_i_16 
       (.I0(sbox_pp2[4]),
        .I1(sbox_pp2[12]),
        .O(\CD[0].col[3][28]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][28]_i_17 
       (.I0(sbox_pp2[15]),
        .I1(sbox_pp2[23]),
        .I2(sbox_pp2[19]),
        .I3(sbox_pp2[27]),
        .I4(sbox_pp2[25]),
        .I5(sbox_pp2[9]),
        .O(\CD[0].col[3][28]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][28]_i_19 
       (.I0(\CD[0].col[3][1]_i_17_n_0 ),
        .I1(\CD[0].col[3][3]_i_17_n_0 ),
        .I2(sbox_pp2[20]),
        .I3(sbox_pp2[26]),
        .I4(\CD[0].col[3][28]_i_16_n_0 ),
        .I5(sbox_pp2[10]),
        .O(\CD[0].col[3][28]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][28]_i_3 
       (.I0(key_out[18]),
        .I1(add_rd_key_in[28]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[28]),
        .I5(sbox_pp2[28]),
        .O(last_round_pp2_reg_0[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][28]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [28]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [28]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][28]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][28]_i_6 
       (.I0(bus_swap[28]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][28]_i_12_n_0 ),
        .I3(add_rd_key_in[28]),
        .I4(key_out[18]),
        .I5(add_rk_sel),
        .O(enable_i_12_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][28]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_144),
        .I2(\CD[0].col[3][28]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[28]),
        .I5(\CD[0].col[3][28]_i_14_n_0 ),
        .O(add_rd_key_in[28]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][28]_i_9 
       (.I0(\CD[0].col[3][28]_i_15_n_0 ),
        .I1(sbox_pp2[10]),
        .I2(\CD[0].col[3][28]_i_16_n_0 ),
        .I3(sbox_pp2[26]),
        .I4(sbox_pp2[20]),
        .I5(\CD[0].col[3][28]_i_17_n_0 ),
        .O(mix_out_dec[28]));
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][29]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [25]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [29]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][29]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][29]_i_12 
       (.I0(sbox_pp2[29]),
        .I1(\CD[0].col[3][29]_i_16_n_0 ),
        .I2(\CD[0].col[3][29]_i_17_n_0 ),
        .I3(\CD[0].col[3][29]_i_20_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][29]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][29]_i_13 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [25]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][29]_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][29]_i_15 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[20]),
        .I2(sbox_pp2[28]),
        .I3(sbox_pp2[13]),
        .I4(sbox_pp2[5]),
        .I5(sbox_pp2[21]),
        .O(\CD[0].col[3][29]_i_15_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair269" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CD[0].col[3][29]_i_16 
       (.I0(sbox_pp2[18]),
        .I1(sbox_pp2[10]),
        .I2(sbox_pp2[27]),
        .O(\CD[0].col[3][29]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][29]_i_17 
       (.I0(sbox_pp2[23]),
        .I1(sbox_pp2[7]),
        .I2(sbox_pp2[2]),
        .I3(sbox_pp2[26]),
        .I4(\CD[0].col[3][30]_i_17_n_0 ),
        .I5(\CD[0].col[3][24]_i_16_n_0 ),
        .O(\CD[0].col[3][29]_i_17_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][29]_i_18 
       (.I0(sbox_pp2[20]),
        .I1(sbox_pp2[28]),
        .O(\CD[0].col[3][29]_i_18_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][29]_i_19 
       (.I0(sbox_pp2[5]),
        .I1(sbox_pp2[13]),
        .O(\CD[0].col[3][29]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][29]_i_20 
       (.I0(sbox_pp2[5]),
        .I1(sbox_pp2[13]),
        .I2(sbox_pp2[20]),
        .I3(sbox_pp2[28]),
        .I4(sbox_pp2[11]),
        .I5(sbox_pp2[21]),
        .O(\CD[0].col[3][29]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][29]_i_3 
       (.I0(key_out[19]),
        .I1(add_rd_key_in[29]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[29]),
        .I5(sbox_pp2[29]),
        .O(last_round_pp2_reg_0[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][29]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [29]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [29]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][29]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][29]_i_6 
       (.I0(bus_swap[29]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][29]_i_12_n_0 ),
        .I3(add_rd_key_in[29]),
        .I4(key_out[19]),
        .I5(add_rk_sel),
        .O(enable_i_13_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][29]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][29]_0 ),
        .I2(\CD[0].col[3][29]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[29]),
        .I5(\CD[0].col[3][29]_i_15_n_0 ),
        .O(add_rd_key_in[29]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][29]_i_9 
       (.I0(\CD[0].col[3][29]_i_16_n_0 ),
        .I1(\CD[0].col[3][29]_i_17_n_0 ),
        .I2(sbox_pp2[21]),
        .I3(sbox_pp2[11]),
        .I4(\CD[0].col[3][29]_i_18_n_0 ),
        .I5(\CD[0].col[3][29]_i_19_n_0 ),
        .O(mix_out_dec[29]));
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][2]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3]_4 [2]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [2]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][2]_1 ));
  LUT5 #(
    .INIT(32'h00AA003C)) 
    \CD[0].col[3][2]_i_13 
       (.I0(sbox_pp2[2]),
        .I1(\CD[0].col[3][26]_i_17_n_0 ),
        .I2(\CD[0].col[3][2]_i_19_n_0 ),
        .I3(add_rk_sel),
        .I4(last_round_pp2),
        .O(\CD[0].col[3][2]_i_13_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][2]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3]_4 [2]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][2]_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][2]_i_17 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[18]),
        .I2(sbox_pp2[10]),
        .I3(sbox_pp2[25]),
        .I4(sbox_pp2[1]),
        .I5(sbox_pp2[26]),
        .O(\CD[0].col[3][2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][2]_i_18 
       (.I0(sbox_pp2[15]),
        .I1(sbox_pp2[31]),
        .I2(sbox_pp2[30]),
        .I3(sbox_pp2[14]),
        .I4(sbox_pp2[22]),
        .I5(sbox_pp2[6]),
        .O(\CD[0].col[3][2]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][2]_i_19 
       (.I0(\CD[0].col[3][26]_i_21_n_0 ),
        .I1(\CD[0].col[3][2]_i_21_n_0 ),
        .I2(sbox_pp2[16]),
        .I3(sbox_pp2[26]),
        .I4(sbox_pp2[0]),
        .I5(sbox_pp2[1]),
        .O(\CD[0].col[3][2]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][2]_i_21 
       (.I0(sbox_pp2[31]),
        .I1(sbox_pp2[15]),
        .O(\CD[0].col[3][2]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][2]_i_3 
       (.I0(\sbox_pp2[2]_i_3_n_0 ),
        .I1(add_rd_key_in[2]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[2]),
        .I5(sbox_pp2[2]),
        .O(add_rk_out[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][2]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [2]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [2]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][2]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][2]_i_6 
       (.I0(bus_swap[2]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][2]_i_13_n_0 ),
        .I3(add_rd_key_in[2]),
        .I4(\sbox_pp2[2]_i_3_n_0 ),
        .I5(add_rk_sel),
        .O(enable_i_18_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][2]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_137),
        .I2(\CD[0].col[3][2]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[2]),
        .I5(\CD[0].col[3][2]_i_17_n_0 ),
        .O(add_rd_key_in[2]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][2]_i_9 
       (.I0(\CD[0].col[3][26]_i_17_n_0 ),
        .I1(sbox_pp2[1]),
        .I2(sbox_pp2[0]),
        .I3(sbox_pp2[26]),
        .I4(sbox_pp2[16]),
        .I5(\CD[0].col[3][2]_i_18_n_0 ),
        .O(mix_out_dec[2]));
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][30]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [26]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [30]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][30]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][30]_i_12 
       (.I0(sbox_pp2[30]),
        .I1(\CD[0].col[3][30]_i_19_n_0 ),
        .I2(\CD[0].col[3][30]_i_17_n_0 ),
        .I3(\CD[0].col[3][30]_i_18_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][30]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][30]_i_13 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [26]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][30]_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][30]_i_15 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[22]),
        .I2(sbox_pp2[6]),
        .I3(sbox_pp2[29]),
        .I4(sbox_pp2[21]),
        .I5(sbox_pp2[14]),
        .O(\CD[0].col[3][30]_i_15_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][30]_i_16 
       (.I0(sbox_pp2[21]),
        .I1(sbox_pp2[29]),
        .O(\CD[0].col[3][30]_i_16_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][30]_i_17 
       (.I0(sbox_pp2[22]),
        .I1(sbox_pp2[6]),
        .O(\CD[0].col[3][30]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][30]_i_18 
       (.I0(\CD[0].col[3][12]_i_13_n_0 ),
        .I1(sbox_pp2[3]),
        .I2(sbox_pp2[11]),
        .I3(\CD[0].col[3][31]_i_35_n_0 ),
        .I4(sbox_pp2[19]),
        .I5(sbox_pp2[27]),
        .O(\CD[0].col[3][30]_i_18_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CD[0].col[3][30]_i_19 
       (.I0(sbox_pp2[28]),
        .I1(sbox_pp2[21]),
        .I2(sbox_pp2[29]),
        .I3(sbox_pp2[12]),
        .I4(sbox_pp2[14]),
        .O(\CD[0].col[3][30]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][30]_i_3 
       (.I0(key_out[20]),
        .I1(add_rd_key_in[30]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[30]),
        .I5(sbox_pp2[30]),
        .O(last_round_pp2_reg_0[14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][30]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [30]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [30]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][30]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][30]_i_6 
       (.I0(bus_swap[30]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][30]_i_12_n_0 ),
        .I3(add_rd_key_in[30]),
        .I4(key_out[20]),
        .I5(add_rk_sel),
        .O(enable_i_14_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][30]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][30]_0 ),
        .I2(\base_new_pp_reg[4]_2 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[30]),
        .I5(\CD[0].col[3][30]_i_15_n_0 ),
        .O(add_rd_key_in[30]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][30]_i_9 
       (.I0(sbox_pp2[14]),
        .I1(sbox_pp2[12]),
        .I2(\CD[0].col[3][30]_i_16_n_0 ),
        .I3(sbox_pp2[28]),
        .I4(\CD[0].col[3][30]_i_17_n_0 ),
        .I5(\CD[0].col[3][30]_i_18_n_0 ),
        .O(mix_out_dec[30]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][31]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [31]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [31]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][31]_i_12 
       (.I0(bus_swap[31]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][31]_i_25_n_0 ),
        .I3(add_rd_key_in[31]),
        .I4(key_out[21]),
        .I5(add_rk_sel),
        .O(enable_i_15_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][31]_i_14 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_132),
        .I2(\CD[0].col[3][31]_i_12_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[31]),
        .I5(\CD[0].col[3][31]_i_32_n_0 ),
        .O(add_rd_key_in[31]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][31]_i_16 
       (.I0(\CD[0].col[3][31]_i_33_n_0 ),
        .I1(sbox_pp2[22]),
        .I2(sbox_pp2[30]),
        .I3(\CD[0].col[3][31]_i_34_n_0 ),
        .I4(\CD[0].col[3][31]_i_35_n_0 ),
        .I5(sbox_pp2[7]),
        .O(mix_out_dec[31]));
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][31]_i_20 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [27]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [31]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][31]_2 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][31]_i_25 
       (.I0(sbox_pp2[31]),
        .I1(\CD[0].col[3][28]_i_16_n_0 ),
        .I2(\CD[0].col[3][29]_i_18_n_0 ),
        .I3(\CD[0].col[3][31]_i_37_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][31]_i_25_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][31]_i_26 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [27]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][31]_1 ));
  LUT4 #(
    .INIT(16'h111F)) 
    \CD[0].col[3][31]_i_29 
       (.I0(rk_sel_pp2[0]),
        .I1(rk_sel_pp2[1]),
        .I2(\CD[0].col[3][9]_i_8_1 [1]),
        .I3(\CD[0].col[3][9]_i_8_1 [0]),
        .O(\CD[0].col[3][31]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h2220)) 
    \CD[0].col[3][31]_i_31 
       (.I0(rk_sel_pp2[0]),
        .I1(rk_sel_pp2[1]),
        .I2(\CD[0].col[3][9]_i_8_1 [1]),
        .I3(\CD[0].col[3][9]_i_8_1 [0]),
        .O(\CD[0].col[3][31]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][31]_i_32 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[30]),
        .I2(sbox_pp2[15]),
        .I3(sbox_pp2[23]),
        .I4(sbox_pp2[7]),
        .I5(sbox_pp2[22]),
        .O(\CD[0].col[3][31]_i_32_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CD[0].col[3][31]_i_33 
       (.I0(sbox_pp2[28]),
        .I1(sbox_pp2[20]),
        .I2(sbox_pp2[12]),
        .I3(sbox_pp2[4]),
        .O(\CD[0].col[3][31]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][31]_i_34 
       (.I0(sbox_pp2[13]),
        .I1(sbox_pp2[29]),
        .O(\CD[0].col[3][31]_i_34_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][31]_i_35 
       (.I0(sbox_pp2[15]),
        .I1(sbox_pp2[23]),
        .O(\CD[0].col[3][31]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][31]_i_37 
       (.I0(sbox_pp2[7]),
        .I1(\CD[0].col[3][31]_i_35_n_0 ),
        .I2(sbox_pp2[13]),
        .I3(sbox_pp2[29]),
        .I4(sbox_pp2[30]),
        .I5(sbox_pp2[22]),
        .O(\CD[0].col[3][31]_i_37_n_0 ));
  LUT4 #(
    .INIT(16'h2220)) 
    \CD[0].col[3][31]_i_39 
       (.I0(rk_sel_pp2[1]),
        .I1(rk_sel_pp2[0]),
        .I2(\CD[0].col[3][9]_i_8_1 [1]),
        .I3(\CD[0].col[3][9]_i_8_1 [0]),
        .O(\CD[0].col[3][31]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][31]_i_6 
       (.I0(key_out[21]),
        .I1(add_rd_key_in[31]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[31]),
        .I5(sbox_pp2[31]),
        .O(last_round_pp2_reg_0[15]));
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][3]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3]_4 [3]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [3]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][3]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][3]_i_13 
       (.I0(sbox_pp2[3]),
        .I1(\CD[0].col[3][3]_i_18_n_0 ),
        .I2(\CD[0].col[3][3]_i_17_n_0 ),
        .I3(\CD[0].col[3][28]_i_15_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][3]_i_13_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][3]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3]_4 [3]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][3]_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][3]_i_16 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(\CD[0].col[3][3]_i_19_n_0 ),
        .I2(sbox_pp2[27]),
        .I3(sbox_pp2[19]),
        .I4(\CD[0].col[3][12]_i_13_n_0 ),
        .I5(sbox_pp2[11]),
        .O(\CD[0].col[3][3]_i_16_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CD[0].col[3][3]_i_17 
       (.I0(sbox_pp2[27]),
        .I1(sbox_pp2[19]),
        .I2(sbox_pp2[23]),
        .I3(sbox_pp2[15]),
        .O(\CD[0].col[3][3]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][3]_i_18 
       (.I0(\CD[0].col[3][24]_i_18_n_0 ),
        .I1(sbox_pp2[16]),
        .I2(sbox_pp2[24]),
        .I3(sbox_pp2[11]),
        .I4(sbox_pp2[2]),
        .I5(sbox_pp2[26]),
        .O(\CD[0].col[3][3]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][3]_i_19 
       (.I0(sbox_pp2[2]),
        .I1(sbox_pp2[26]),
        .O(\CD[0].col[3][3]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][3]_i_3 
       (.I0(\sbox_pp2[3]_i_2_n_0 ),
        .I1(add_rd_key_in[3]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[3]),
        .I5(sbox_pp2[3]),
        .O(add_rk_out[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][3]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [3]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [3]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][3]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][3]_i_6 
       (.I0(bus_swap[3]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][3]_i_13_n_0 ),
        .I3(add_rd_key_in[3]),
        .I4(\sbox_pp2[3]_i_2_n_0 ),
        .I5(add_rk_sel),
        .O(enable_i_19_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][3]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_141),
        .I2(\base_new_pp_reg[3] ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[3]),
        .I5(\CD[0].col[3][3]_i_16_n_0 ),
        .O(add_rd_key_in[3]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][3]_i_9 
       (.I0(sbox_pp2[26]),
        .I1(sbox_pp2[2]),
        .I2(sbox_pp2[11]),
        .I3(\CD[0].col[3][27]_i_19_n_0 ),
        .I4(\CD[0].col[3][3]_i_17_n_0 ),
        .I5(\CD[0].col[3][28]_i_15_n_0 ),
        .O(mix_out_dec[3]));
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][4]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [1]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [4]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][4]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][4]_i_12 
       (.I0(sbox_pp2[4]),
        .I1(\CD[1].col[2][21]_i_7_n_0 ),
        .I2(\CD[1].col[2][20]_i_8_n_0 ),
        .I3(\CD[0].col[3][4]_i_17_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][4]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][4]_i_13 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [1]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][4]_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][4]_i_16 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[12]),
        .I2(sbox_pp2[3]),
        .I3(\CD[0].col[3][29]_i_18_n_0 ),
        .I4(\CD[0].col[3][12]_i_13_n_0 ),
        .I5(sbox_pp2[27]),
        .O(\CD[0].col[3][4]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][4]_i_17 
       (.I0(\CD[0].col[3][11]_i_12_n_0 ),
        .I1(\CD[0].col[3][4]_i_19_n_0 ),
        .I2(sbox_pp2[27]),
        .I3(sbox_pp2[2]),
        .I4(\CD[0].col[3][29]_i_18_n_0 ),
        .I5(sbox_pp2[18]),
        .O(\CD[0].col[3][4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][4]_i_19 
       (.I0(sbox_pp2[17]),
        .I1(sbox_pp2[1]),
        .I2(sbox_pp2[5]),
        .I3(sbox_pp2[13]),
        .I4(sbox_pp2[21]),
        .I5(sbox_pp2[29]),
        .O(\CD[0].col[3][4]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][4]_i_3 
       (.I0(\KR[1].key_reg[2][4]_0 ),
        .I1(add_rd_key_in[4]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[4]),
        .I5(sbox_pp2[4]),
        .O(add_rk_out[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][4]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [4]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [4]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][4]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][4]_i_6 
       (.I0(bus_swap[4]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][4]_i_12_n_0 ),
        .I3(add_rd_key_in[4]),
        .I4(\KR[1].key_reg[2][4]_0 ),
        .I5(add_rk_sel),
        .O(enable_i_20_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][4]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_142),
        .I2(\CD[0].col[3][4]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[4]),
        .I5(\CD[0].col[3][4]_i_16_n_0 ),
        .O(add_rd_key_in[4]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][4]_i_9 
       (.I0(sbox_pp2[3]),
        .I1(sbox_pp2[12]),
        .I2(sbox_pp2[25]),
        .I3(sbox_pp2[9]),
        .I4(\CD[0].col[3][24]_i_16_n_0 ),
        .I5(\CD[0].col[3][4]_i_17_n_0 ),
        .O(mix_out_dec[4]));
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][5]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3]_4 [5]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [5]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][5]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][5]_i_13 
       (.I0(sbox_pp2[5]),
        .I1(\CD[0].col[3][5]_i_17_n_0 ),
        .I2(\CD[0].col[3][5]_i_18_n_0 ),
        .I3(\CD[0].col[3][5]_i_21_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][5]_i_13_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][5]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3]_4 [5]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][5]_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][5]_i_16 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[4]),
        .I2(sbox_pp2[13]),
        .I3(sbox_pp2[29]),
        .I4(sbox_pp2[21]),
        .I5(sbox_pp2[28]),
        .O(\CD[0].col[3][5]_i_16_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \CD[0].col[3][5]_i_17 
       (.I0(sbox_pp2[29]),
        .I1(sbox_pp2[21]),
        .I2(sbox_pp2[28]),
        .O(\CD[0].col[3][5]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][5]_i_18 
       (.I0(sbox_pp2[15]),
        .I1(sbox_pp2[31]),
        .I2(sbox_pp2[2]),
        .I3(sbox_pp2[26]),
        .I4(\CD[0].col[3][30]_i_17_n_0 ),
        .I5(\CD[0].col[3][24]_i_16_n_0 ),
        .O(\CD[0].col[3][5]_i_18_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair274" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][5]_i_19 
       (.I0(sbox_pp2[4]),
        .I1(sbox_pp2[13]),
        .O(\CD[0].col[3][5]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][5]_i_20 
       (.I0(sbox_pp2[10]),
        .I1(sbox_pp2[18]),
        .O(\CD[0].col[3][5]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][5]_i_21 
       (.I0(sbox_pp2[10]),
        .I1(sbox_pp2[18]),
        .I2(sbox_pp2[4]),
        .I3(sbox_pp2[13]),
        .I4(sbox_pp2[19]),
        .I5(sbox_pp2[3]),
        .O(\CD[0].col[3][5]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][5]_i_3 
       (.I0(\sbox_pp2[5]_i_3_n_0 ),
        .I1(add_rd_key_in[5]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[5]),
        .I5(sbox_pp2[5]),
        .O(add_rk_out[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][5]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [5]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [5]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][5]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][5]_i_6 
       (.I0(bus_swap[5]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][5]_i_13_n_0 ),
        .I3(add_rd_key_in[5]),
        .I4(\sbox_pp2[5]_i_3_n_0 ),
        .I5(add_rk_sel),
        .O(enable_i_21_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][5]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][5]_0 ),
        .I2(\CD[0].col[3][5]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[5]),
        .I5(\CD[0].col[3][5]_i_16_n_0 ),
        .O(add_rd_key_in[5]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][5]_i_9 
       (.I0(\CD[0].col[3][5]_i_17_n_0 ),
        .I1(\CD[0].col[3][5]_i_18_n_0 ),
        .I2(sbox_pp2[3]),
        .I3(sbox_pp2[19]),
        .I4(\CD[0].col[3][5]_i_19_n_0 ),
        .I5(\CD[0].col[3][5]_i_20_n_0 ),
        .O(mix_out_dec[5]));
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][6]_i_11 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [2]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [6]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][6]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][6]_i_12 
       (.I0(sbox_pp2[6]),
        .I1(\CD[0].col[3][6]_i_17_n_0 ),
        .I2(\CD[0].col[3][30]_i_18_n_0 ),
        .I3(\CD[0].col[3][6]_i_16_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][6]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][6]_i_13 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [2]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][6]_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][6]_i_15 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[22]),
        .I2(sbox_pp2[5]),
        .I3(sbox_pp2[14]),
        .I4(sbox_pp2[30]),
        .I5(sbox_pp2[29]),
        .O(\CD[0].col[3][6]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][6]_i_16 
       (.I0(sbox_pp2[22]),
        .I1(sbox_pp2[5]),
        .O(\CD[0].col[3][6]_i_16_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CD[0].col[3][6]_i_17 
       (.I0(sbox_pp2[29]),
        .I1(sbox_pp2[20]),
        .I2(sbox_pp2[4]),
        .I3(sbox_pp2[30]),
        .I4(sbox_pp2[14]),
        .O(\CD[0].col[3][6]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][6]_i_3 
       (.I0(\KR[1].key_reg[2][6]_0 ),
        .I1(add_rd_key_in[6]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[6]),
        .I5(sbox_pp2[6]),
        .O(add_rk_out[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][6]_i_5 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [6]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [6]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][6]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][6]_i_6 
       (.I0(bus_swap[6]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][6]_i_12_n_0 ),
        .I3(add_rd_key_in[6]),
        .I4(\KR[1].key_reg[2][6]_0 ),
        .I5(add_rk_sel),
        .O(enable_i_22_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][6]_i_8 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][6]_0 ),
        .I2(\base_new_pp_reg[4]_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[6]),
        .I5(\CD[0].col[3][6]_i_15_n_0 ),
        .O(add_rd_key_in[6]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][6]_i_9 
       (.I0(\CD[0].col[3][24]_i_16_n_0 ),
        .I1(sbox_pp2[4]),
        .I2(sbox_pp2[20]),
        .I3(sbox_pp2[29]),
        .I4(\CD[0].col[3][30]_i_18_n_0 ),
        .I5(\CD[0].col[3][6]_i_16_n_0 ),
        .O(mix_out_dec[6]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][7]_i_10 
       (.I0(\CD[0].col[3][31]_i_33_n_0 ),
        .I1(\CD[0].col[3][7]_i_18_n_0 ),
        .I2(sbox_pp2[31]),
        .I3(sbox_pp2[5]),
        .I4(\CD[0].col[3][31]_i_35_n_0 ),
        .I5(sbox_pp2[30]),
        .O(mix_out_dec[7]));
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][7]_i_12 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [3]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [7]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][7]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][7]_i_13 
       (.I0(sbox_pp2[7]),
        .I1(\CD[0].col[3][31]_i_33_n_0 ),
        .I2(\CD[0].col[3][7]_i_18_n_0 ),
        .I3(\CD[0].col[3][7]_i_19_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][7]_i_13_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][7]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [3]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][7]_0 ));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][7]_i_17 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[30]),
        .I2(sbox_pp2[15]),
        .I3(sbox_pp2[23]),
        .I4(sbox_pp2[31]),
        .I5(sbox_pp2[6]),
        .O(\CD[0].col[3][7]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][7]_i_18 
       (.I0(sbox_pp2[6]),
        .I1(sbox_pp2[21]),
        .O(\CD[0].col[3][7]_i_18_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CD[0].col[3][7]_i_19 
       (.I0(sbox_pp2[30]),
        .I1(sbox_pp2[15]),
        .I2(sbox_pp2[23]),
        .I3(sbox_pp2[5]),
        .I4(sbox_pp2[31]),
        .O(\CD[0].col[3][7]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][7]_i_3 
       (.I0(key_out[1]),
        .I1(add_rd_key_in[7]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[7]),
        .I5(sbox_pp2[7]),
        .O(add_rk_out[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][7]_i_6 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [7]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [7]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][7]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][7]_i_7 
       (.I0(bus_swap[7]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][7]_i_13_n_0 ),
        .I3(add_rd_key_in[7]),
        .I4(key_out[1]),
        .I5(add_rk_sel),
        .O(enable_i_23_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][7]_i_9 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_130),
        .I2(\CD[0].col[3][7]_i_7_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[7]),
        .I5(\CD[0].col[3][7]_i_17_n_0 ),
        .O(add_rd_key_in[7]));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][8]_i_10 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[7]),
        .I2(sbox_pp2[15]),
        .I3(sbox_pp2[24]),
        .I4(sbox_pp2[16]),
        .I5(sbox_pp2[0]),
        .O(\CD[0].col[3][8]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[0].col[3][8]_i_11 
       (.I0(sbox_pp2[16]),
        .I1(sbox_pp2[24]),
        .O(\CD[0].col[3][8]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][8]_i_13 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [4]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [8]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][8]_1 ));
  LUT6 #(
    .INIT(64'h0000AAAA0000C33C)) 
    \CD[0].col[3][8]_i_14 
       (.I0(sbox_pp2[8]),
        .I1(\CD[0].col[3][8]_i_17_n_0 ),
        .I2(\CD[0].col[3][24]_i_17_n_0 ),
        .I3(\CD[0].col[3][8]_i_11_n_0 ),
        .I4(add_rk_sel),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][8]_i_14_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][8]_i_15 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [4]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][8]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \CD[0].col[3][8]_i_17 
       (.I0(sbox_pp2[15]),
        .I1(sbox_pp2[7]),
        .I2(sbox_pp2[0]),
        .I3(sbox_pp2[30]),
        .I4(sbox_pp2[14]),
        .O(\CD[0].col[3][8]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][8]_i_2 
       (.I0(key_out[2]),
        .I1(add_rd_key_in[8]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[8]),
        .I5(sbox_pp2[8]),
        .O(last_round_pp2_reg_0[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][8]_i_4 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][8]_0 ),
        .I2(\CD[0].col[3][8]_i_8_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[8]),
        .I5(\CD[0].col[3][8]_i_10_n_0 ),
        .O(add_rd_key_in[8]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][8]_i_5 
       (.I0(\CD[0].col[3][24]_i_16_n_0 ),
        .I1(sbox_pp2[0]),
        .I2(sbox_pp2[7]),
        .I3(sbox_pp2[15]),
        .I4(\CD[0].col[3][24]_i_17_n_0 ),
        .I5(\CD[0].col[3][8]_i_11_n_0 ),
        .O(mix_out_dec[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][8]_i_7 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [8]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [8]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][8]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][8]_i_8 
       (.I0(bus_swap[8]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][8]_i_14_n_0 ),
        .I3(add_rd_key_in[8]),
        .I4(key_out[2]),
        .I5(add_rk_sel),
        .O(enable_i_24_sn_1));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[0].col[3][9]_i_10 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(\CD[0].col[3][27]_i_20_n_0 ),
        .I2(sbox_pp2[17]),
        .I3(sbox_pp2[1]),
        .I4(\CD[0].col[3][24]_i_18_n_0 ),
        .I5(sbox_pp2[25]),
        .O(\CD[0].col[3][9]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT4 #(
    .INIT(16'hAAC0)) 
    \CD[0].col[3][9]_i_12 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [5]),
        .I1(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [9]),
        .I2(iv_mux_out13_out),
        .I3(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][9]_1 ));
  LUT6 #(
    .INIT(64'h0000AAA00000CCC0)) 
    \CD[0].col[3][9]_i_13 
       (.I0(sbox_pp2[9]),
        .I1(mix_out_dec[9]),
        .I2(\CD[0].col[3][9]_i_8_1 [0]),
        .I3(\CD[0].col[3][9]_i_8_1 [1]),
        .I4(rk_out_sel_pp2),
        .I5(last_round_pp2),
        .O(\CD[0].col[3][9]_i_13_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \CD[0].col[3][9]_i_14 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [5]),
        .I1(\CD[0].col[3][5]_i_7 ),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][9]_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[0].col[3][9]_i_2 
       (.I0(\KR[1].key_reg[2][9]_0 ),
        .I1(add_rd_key_in[9]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[9]),
        .I5(sbox_pp2[9]),
        .O(last_round_pp2_reg_0[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[0].col[3][9]_i_4 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][9]_0 ),
        .I2(\CD[0].col[3][9]_i_8_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[9]),
        .I5(\CD[0].col[3][9]_i_10_n_0 ),
        .O(add_rd_key_in[9]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[0].col[3][9]_i_5 
       (.I0(sbox_pp2[25]),
        .I1(sbox_pp2[7]),
        .I2(sbox_pp2[31]),
        .I3(sbox_pp2[0]),
        .I4(sbox_pp2[8]),
        .I5(\CD[0].col[3][28]_i_15_n_0 ),
        .O(mix_out_dec[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \CD[0].col[3][9]_i_7 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [9]),
        .I1(\CD[0].col[3][0]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [9]),
        .I3(\CD[0].col[3][31]_i_5 ),
        .O(\IV_BKP_REGISTERS[3].bkp_reg[3][9]_0 ));
  LUT6 #(
    .INIT(64'h4744444747474747)) 
    \CD[0].col[3][9]_i_8 
       (.I0(bus_swap[9]),
        .I1(\CD[0].col[3][0]_i_2 ),
        .I2(\CD[0].col[3][9]_i_13_n_0 ),
        .I3(add_rd_key_in[9]),
        .I4(\KR[1].key_reg[2][9]_0 ),
        .I5(add_rk_sel),
        .O(enable_i_25_sn_1));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][0] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [0]),
        .Q(Q[0]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][10] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [10]),
        .Q(Q[10]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][11] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [11]),
        .Q(Q[11]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][12] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [12]),
        .Q(Q[12]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][13] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [13]),
        .Q(Q[13]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][14] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [14]),
        .Q(Q[14]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][15] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [15]),
        .Q(Q[15]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][16] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [16]),
        .Q(Q[16]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][17] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [17]),
        .Q(Q[17]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][18] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [18]),
        .Q(Q[18]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][19] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [19]),
        .Q(Q[19]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][1] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [1]),
        .Q(Q[1]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][20] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [20]),
        .Q(Q[20]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][21] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [21]),
        .Q(Q[21]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][22] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [22]),
        .Q(Q[22]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][23] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [23]),
        .Q(Q[23]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][24] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [24]),
        .Q(Q[24]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][25] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [25]),
        .Q(Q[25]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][26] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [26]),
        .Q(Q[26]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][27] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [27]),
        .Q(Q[27]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][28] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [28]),
        .Q(Q[28]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][29] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [29]),
        .Q(Q[29]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][2] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [2]),
        .Q(Q[2]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][30] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [30]),
        .Q(Q[30]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][31] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [31]),
        .Q(Q[31]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][3] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [3]),
        .Q(Q[3]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][4] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [4]),
        .Q(Q[4]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][5] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [5]),
        .Q(Q[5]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][6] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [6]),
        .Q(Q[6]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][7] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [7]),
        .Q(Q[7]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][8] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [8]),
        .Q(Q[8]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[0].col_reg[3][9] 
       (.C(clk_i),
        .CE(\CD[0].col_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [9]),
        .Q(Q[9]));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[1].col[2][16]_i_2 
       (.I0(key_out[6]),
        .I1(add_rd_key_in[16]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[16]),
        .I5(sbox_pp2[16]),
        .O(add_rk_out[8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[1].col[2][16]_i_3 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][16]_0 ),
        .I2(\CD[0].col[3][16]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[16]),
        .I5(\CD[1].col[2][16]_i_5_n_0 ),
        .O(add_rd_key_in[16]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[1].col[2][16]_i_4 
       (.I0(\CD[0].col[3][30]_i_17_n_0 ),
        .I1(sbox_pp2[24]),
        .I2(sbox_pp2[0]),
        .I3(sbox_pp2[8]),
        .I4(\CD[0].col[3][24]_i_17_n_0 ),
        .I5(\CD[0].col[3][31]_i_35_n_0 ),
        .O(mix_out_dec[16]));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[1].col[2][16]_i_5 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[15]),
        .I2(sbox_pp2[23]),
        .I3(sbox_pp2[8]),
        .I4(sbox_pp2[0]),
        .I5(sbox_pp2[24]),
        .O(\CD[1].col[2][16]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[1].col[2][17]_i_2 
       (.I0(key_out[7]),
        .I1(add_rd_key_in[17]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[17]),
        .I5(sbox_pp2[17]),
        .O(add_rk_out[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[1].col[2][17]_i_3 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][17]_0 ),
        .I2(\CD[0].col[3][17]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[17]),
        .I5(\CD[1].col[2][17]_i_5_n_0 ),
        .O(add_rd_key_in[17]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[1].col[2][17]_i_4 
       (.I0(sbox_pp2[16]),
        .I1(sbox_pp2[7]),
        .I2(sbox_pp2[15]),
        .I3(\CD[0].col[3][27]_i_16_n_0 ),
        .I4(sbox_pp2[1]),
        .I5(sbox_pp2[8]),
        .O(mix_out_dec[17]));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[1].col[2][17]_i_5 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[8]),
        .I2(sbox_pp2[1]),
        .I3(\CD[0].col[3][1]_i_17_n_0 ),
        .I4(\CD[0].col[3][31]_i_35_n_0 ),
        .I5(sbox_pp2[16]),
        .O(\CD[1].col[2][17]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[1].col[2][18]_i_2 
       (.I0(key_out[8]),
        .I1(add_rd_key_in[18]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[18]),
        .I5(sbox_pp2[18]),
        .O(add_rk_out[10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[1].col[2][18]_i_3 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_158),
        .I2(\CD[0].col[3][18]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[18]),
        .I5(\CD[1].col[2][18]_i_6_n_0 ),
        .O(add_rd_key_in[18]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[1].col[2][18]_i_4 
       (.I0(sbox_pp2[9]),
        .I1(sbox_pp2[16]),
        .I2(\CD[0].col[3][5]_i_18_n_0 ),
        .I3(sbox_pp2[10]),
        .I4(sbox_pp2[0]),
        .I5(sbox_pp2[17]),
        .O(mix_out_dec[18]));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[1].col[2][18]_i_6 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[26]),
        .I2(sbox_pp2[2]),
        .I3(sbox_pp2[10]),
        .I4(sbox_pp2[9]),
        .I5(sbox_pp2[17]),
        .O(\CD[1].col[2][18]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[1].col[2][19]_i_2 
       (.I0(key_out[9]),
        .I1(add_rd_key_in[19]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[19]),
        .I5(sbox_pp2[19]),
        .O(add_rk_out[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[1].col[2][19]_i_3 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_157),
        .I2(\base_new_pp_reg[3]_2 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[19]),
        .I5(\CD[1].col[2][19]_i_5_n_0 ),
        .O(add_rd_key_in[19]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[1].col[2][19]_i_4 
       (.I0(sbox_pp2[11]),
        .I1(sbox_pp2[3]),
        .I2(\CD[0].col[3][12]_i_13_n_0 ),
        .I3(\CD[0].col[3][28]_i_15_n_0 ),
        .I4(\CD[0].col[3][27]_i_19_n_0 ),
        .I5(\CD[0].col[3][29]_i_16_n_0 ),
        .O(mix_out_dec[19]));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[1].col[2][19]_i_5 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(\CD[0].col[3][29]_i_16_n_0 ),
        .I2(sbox_pp2[23]),
        .I3(sbox_pp2[15]),
        .I4(sbox_pp2[11]),
        .I5(sbox_pp2[3]),
        .O(\CD[1].col[2][19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[1].col[2][20]_i_2 
       (.I0(key_out[10]),
        .I1(add_rd_key_in[20]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[20]),
        .I5(sbox_pp2[20]),
        .O(add_rk_out[12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[1].col[2][20]_i_3 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_156),
        .I2(\CD[0].col[3][20]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[20]),
        .I5(\CD[1].col[2][20]_i_6_n_0 ),
        .O(add_rd_key_in[20]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[1].col[2][20]_i_4 
       (.I0(sbox_pp2[11]),
        .I1(\CD[0].col[3][28]_i_16_n_0 ),
        .I2(\CD[1].col[2][20]_i_7_n_0 ),
        .I3(sbox_pp2[19]),
        .I4(sbox_pp2[18]),
        .I5(\CD[1].col[2][20]_i_8_n_0 ),
        .O(mix_out_dec[20]));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[1].col[2][20]_i_6 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[11]),
        .I2(\CD[0].col[3][28]_i_16_n_0 ),
        .I3(\CD[0].col[3][31]_i_35_n_0 ),
        .I4(sbox_pp2[28]),
        .I5(sbox_pp2[19]),
        .O(\CD[1].col[2][20]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[1].col[2][20]_i_7 
       (.I0(\CD[0].col[3][27]_i_20_n_0 ),
        .I1(sbox_pp2[17]),
        .I2(sbox_pp2[1]),
        .I3(\CD[0].col[3][24]_i_17_n_0 ),
        .I4(sbox_pp2[2]),
        .I5(sbox_pp2[28]),
        .O(\CD[1].col[2][20]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \CD[1].col[2][20]_i_8 
       (.I0(sbox_pp2[25]),
        .I1(sbox_pp2[9]),
        .I2(sbox_pp2[14]),
        .I3(sbox_pp2[30]),
        .O(\CD[1].col[2][20]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[1].col[2][21]_i_2 
       (.I0(key_out[11]),
        .I1(add_rd_key_in[21]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[21]),
        .I5(sbox_pp2[21]),
        .O(add_rk_out[13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[1].col[2][21]_i_3 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][21]_0 ),
        .I2(\CD[0].col[3][21]_i_6_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[21]),
        .I5(\CD[1].col[2][21]_i_5_n_0 ),
        .O(add_rd_key_in[21]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[1].col[2][21]_i_4 
       (.I0(\CD[1].col[2][21]_i_6_n_0 ),
        .I1(\CD[0].col[3][5]_i_18_n_0 ),
        .I2(\CD[0].col[3][29]_i_19_n_0 ),
        .I3(sbox_pp2[19]),
        .I4(\CD[1].col[2][21]_i_7_n_0 ),
        .I5(\CD[0].col[3][5]_i_20_n_0 ),
        .O(mix_out_dec[21]));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[1].col[2][21]_i_5 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[20]),
        .I2(sbox_pp2[29]),
        .I3(sbox_pp2[13]),
        .I4(sbox_pp2[5]),
        .I5(sbox_pp2[12]),
        .O(\CD[1].col[2][21]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[1].col[2][21]_i_6 
       (.I0(sbox_pp2[20]),
        .I1(sbox_pp2[29]),
        .O(\CD[1].col[2][21]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair273" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \CD[1].col[2][21]_i_7 
       (.I0(sbox_pp2[3]),
        .I1(sbox_pp2[12]),
        .O(\CD[1].col[2][21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[1].col[2][22]_i_2 
       (.I0(key_out[12]),
        .I1(add_rd_key_in[22]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[22]),
        .I5(sbox_pp2[22]),
        .O(add_rk_out[14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[1].col[2][22]_i_3 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(\CD[2].col_reg[1][22]_0 ),
        .I2(\base_new_pp_reg[4]_3 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[22]),
        .I5(\CD[1].col[2][22]_i_5_n_0 ),
        .O(add_rd_key_in[22]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[1].col[2][22]_i_4 
       (.I0(\CD[0].col[3][24]_i_16_n_0 ),
        .I1(sbox_pp2[20]),
        .I2(\CD[0].col[3][7]_i_18_n_0 ),
        .I3(\CD[0].col[3][30]_i_18_n_0 ),
        .I4(sbox_pp2[4]),
        .I5(sbox_pp2[13]),
        .O(mix_out_dec[22]));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[1].col[2][22]_i_5 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[6]),
        .I2(sbox_pp2[21]),
        .I3(sbox_pp2[14]),
        .I4(sbox_pp2[30]),
        .I5(sbox_pp2[13]),
        .O(\CD[1].col[2][22]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h66FF66F0660F6600)) 
    \CD[1].col[2][23]_i_2 
       (.I0(key_out[13]),
        .I1(add_rd_key_in[23]),
        .I2(last_round_pp2),
        .I3(add_rk_sel),
        .I4(mix_out_dec[23]),
        .I5(sbox_pp2[23]),
        .O(add_rk_out[15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8A8A8)) 
    \CD[1].col[2][23]_i_3 
       (.I0(\CD[0].col[3][31]_i_29_n_0 ),
        .I1(SBOX_n_153),
        .I2(\CD[0].col[3][23]_i_7_0 ),
        .I3(\CD[0].col[3][31]_i_31_n_0 ),
        .I4(sbox_pp2[23]),
        .I5(\CD[1].col[2][23]_i_6_n_0 ),
        .O(add_rd_key_in[23]));
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \CD[1].col[2][23]_i_4 
       (.I0(\CD[0].col[3][31]_i_33_n_0 ),
        .I1(\CD[0].col[3][6]_i_16_n_0 ),
        .I2(sbox_pp2[15]),
        .I3(sbox_pp2[21]),
        .I4(\CD[0].col[3][12]_i_13_n_0 ),
        .I5(sbox_pp2[14]),
        .O(mix_out_dec[23]));
  LUT6 #(
    .INIT(64'h8228288228828228)) 
    \CD[1].col[2][23]_i_6 
       (.I0(\CD[0].col[3][31]_i_39_n_0 ),
        .I1(sbox_pp2[15]),
        .I2(sbox_pp2[7]),
        .I3(sbox_pp2[31]),
        .I4(sbox_pp2[22]),
        .I5(sbox_pp2[14]),
        .O(\CD[1].col[2][23]_i_6_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][0] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [0]),
        .Q(\CD[1].col_reg[2][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][10] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [10]),
        .Q(\CD[1].col_reg[2][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][11] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [11]),
        .Q(\CD[1].col_reg[2][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][12] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [12]),
        .Q(\CD[1].col_reg[2][31]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][13] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [13]),
        .Q(\CD[1].col_reg[2][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][14] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [14]),
        .Q(\CD[1].col_reg[2][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][15] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [15]),
        .Q(\CD[1].col_reg[2][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][16] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [16]),
        .Q(\CD[1].col_reg[2][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][17] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [17]),
        .Q(\CD[1].col_reg[2][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][18] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [18]),
        .Q(\CD[1].col_reg[2][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][19] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [19]),
        .Q(\CD[1].col_reg[2][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][1] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [1]),
        .Q(\CD[1].col_reg[2][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][20] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [20]),
        .Q(\CD[1].col_reg[2][31]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][21] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [21]),
        .Q(\CD[1].col_reg[2][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][22] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [22]),
        .Q(\CD[1].col_reg[2][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][23] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [23]),
        .Q(\CD[1].col_reg[2][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][24] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [24]),
        .Q(\CD[1].col_reg[2][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][25] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [25]),
        .Q(\CD[1].col_reg[2][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][26] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [26]),
        .Q(\CD[1].col_reg[2][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][27] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [27]),
        .Q(\CD[1].col_reg[2][31]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][28] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [28]),
        .Q(\CD[1].col_reg[2][31]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][29] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [29]),
        .Q(\CD[1].col_reg[2][31]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][2] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [2]),
        .Q(\CD[1].col_reg[2][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][30] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [30]),
        .Q(\CD[1].col_reg[2][31]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][31] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [31]),
        .Q(\CD[1].col_reg[2][31]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][3] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [3]),
        .Q(\CD[1].col_reg[2][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][4] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [4]),
        .Q(\CD[1].col_reg[2][31]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][5] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [5]),
        .Q(\CD[1].col_reg[2][31]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][6] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [6]),
        .Q(\CD[1].col_reg[2][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][7] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [7]),
        .Q(\CD[1].col_reg[2][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][8] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [8]),
        .Q(\CD[1].col_reg[2][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[1].col_reg[2][9] 
       (.C(clk_i),
        .CE(\CD[1].col_reg[2][31]_1 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [9]),
        .Q(\CD[1].col_reg[2][31]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][0] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [0]),
        .Q(\CD[2].col_reg[1][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][10] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [10]),
        .Q(\CD[2].col_reg[1][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][11] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [11]),
        .Q(\CD[2].col_reg[1][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][12] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [12]),
        .Q(\CD[2].col_reg[1][31]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][13] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [13]),
        .Q(\CD[2].col_reg[1][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][14] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [14]),
        .Q(\CD[2].col_reg[1][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][15] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [15]),
        .Q(\CD[2].col_reg[1][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][16] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [16]),
        .Q(\CD[2].col_reg[1][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][17] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [17]),
        .Q(\CD[2].col_reg[1][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][18] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [18]),
        .Q(\CD[2].col_reg[1][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][19] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [19]),
        .Q(\CD[2].col_reg[1][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][1] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [1]),
        .Q(\CD[2].col_reg[1][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][20] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [20]),
        .Q(\CD[2].col_reg[1][31]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][21] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [21]),
        .Q(\CD[2].col_reg[1][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][22] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [22]),
        .Q(\CD[2].col_reg[1][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][23] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [23]),
        .Q(\CD[2].col_reg[1][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][24] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [24]),
        .Q(\CD[2].col_reg[1][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][25] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [25]),
        .Q(\CD[2].col_reg[1][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][26] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [26]),
        .Q(\CD[2].col_reg[1][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][27] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [27]),
        .Q(\CD[2].col_reg[1][31]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][28] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [28]),
        .Q(\CD[2].col_reg[1][31]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][29] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [29]),
        .Q(\CD[2].col_reg[1][31]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][2] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [2]),
        .Q(\CD[2].col_reg[1][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][30] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [30]),
        .Q(\CD[2].col_reg[1][31]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][31] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [31]),
        .Q(\CD[2].col_reg[1][31]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][3] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [3]),
        .Q(\CD[2].col_reg[1][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][4] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [4]),
        .Q(\CD[2].col_reg[1][31]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][5] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [5]),
        .Q(\CD[2].col_reg[1][31]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][6] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [6]),
        .Q(\CD[2].col_reg[1][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][7] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [7]),
        .Q(\CD[2].col_reg[1][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][8] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [8]),
        .Q(\CD[2].col_reg[1][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[2].col_reg[1][9] 
       (.C(clk_i),
        .CE(\CD[2].col_reg[1][31]_1 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [9]),
        .Q(\CD[2].col_reg[1][31]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][0] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [0]),
        .Q(\CD[3].col_reg[0][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][10] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [10]),
        .Q(\CD[3].col_reg[0][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][11] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [11]),
        .Q(\CD[3].col_reg[0][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][12] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [12]),
        .Q(\CD[3].col_reg[0][31]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][13] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [13]),
        .Q(\CD[3].col_reg[0][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][14] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [14]),
        .Q(\CD[3].col_reg[0][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][15] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [15]),
        .Q(\CD[3].col_reg[0][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][16] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [16]),
        .Q(\CD[3].col_reg[0][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][17] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [17]),
        .Q(\CD[3].col_reg[0][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][18] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [18]),
        .Q(\CD[3].col_reg[0][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][19] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [19]),
        .Q(\CD[3].col_reg[0][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][1] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [1]),
        .Q(\CD[3].col_reg[0][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][20] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [20]),
        .Q(\CD[3].col_reg[0][31]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][21] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [21]),
        .Q(\CD[3].col_reg[0][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][22] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [22]),
        .Q(\CD[3].col_reg[0][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][23] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [23]),
        .Q(\CD[3].col_reg[0][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][24] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [24]),
        .Q(\CD[3].col_reg[0][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][25] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [25]),
        .Q(\CD[3].col_reg[0][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][26] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [26]),
        .Q(\CD[3].col_reg[0][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][27] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [27]),
        .Q(\CD[3].col_reg[0][31]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][28] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [28]),
        .Q(\CD[3].col_reg[0][31]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][29] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [29]),
        .Q(\CD[3].col_reg[0][31]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][2] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [2]),
        .Q(\CD[3].col_reg[0][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][30] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [30]),
        .Q(\CD[3].col_reg[0][31]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][31] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [31]),
        .Q(\CD[3].col_reg[0][31]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][3] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [3]),
        .Q(\CD[3].col_reg[0][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][4] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [4]),
        .Q(\CD[3].col_reg[0][31]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][5] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [5]),
        .Q(\CD[3].col_reg[0][31]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][6] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [6]),
        .Q(\CD[3].col_reg[0][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][7] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [7]),
        .Q(\CD[3].col_reg[0][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][8] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [8]),
        .Q(\CD[3].col_reg[0][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \CD[3].col_reg[0][9] 
       (.C(clk_i),
        .CE(\CD[3].col_reg[0][31]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [9]),
        .Q(\CD[3].col_reg[0][31]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][0] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [0]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][10] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [10]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][11] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [11]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][12] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [12]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][13] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [13]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][14] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [14]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][15] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [15]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][16] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [16]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][17] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [17]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][18] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [18]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][19] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [19]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][1] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [1]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][20] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [20]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][21] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [21]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][22] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [22]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][23] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [23]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][24] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [24]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][25] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [25]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][26] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [26]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][27] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [27]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][28] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [28]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][29] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [29]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][2] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [2]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][30] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [30]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][31] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [31]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][3] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [3]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][4] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [4]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][5] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [5]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][6] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [6]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][7] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [7]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][8] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [8]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][9] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\CD[0].col_reg[3][31]_1 [9]),
        .Q(\IV_BKP_REGISTERS[0].bkp_1_reg[0][31]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][0] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [0]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][10] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [10]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][11] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [11]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][12] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [12]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][13] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [13]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][14] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [14]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][15] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [15]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][16] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [16]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][17] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [17]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][18] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [18]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][19] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [19]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][1] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [1]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][20] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [20]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][21] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [21]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][22] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [22]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][23] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [23]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][24] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [24]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][25] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [25]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][26] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [26]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][27] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [27]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][28] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [28]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][29] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [29]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][2] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [2]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][30] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [30]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][31] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [31]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][3] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [3]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][4] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [4]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][5] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [5]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][6] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [6]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][7] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [7]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][8] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [8]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].bkp_reg[0][9] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[0].bkp_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_1 [9]),
        .Q(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][0] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][10] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][11] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][12] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][13] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][14] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][15] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][16] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][17] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][18] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][19] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][1] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][20] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][21] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][22] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][23] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][24] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][25] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][26] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][27] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][28] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][29] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][2] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][30] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][31] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][3] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][4] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][5] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][6] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][7] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][8] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[0].iv_reg[0][9] 
       (.C(clk_i),
        .CE(iv_en[0]),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(\IV_BKP_REGISTERS[0].iv_reg[0][31]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][0] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [0]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][10] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [10]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][11] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [11]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][12] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [12]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][13] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [13]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][14] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [14]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][15] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [15]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][16] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [16]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][17] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [17]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][18] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [18]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][19] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [19]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][1] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [1]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][20] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [20]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][21] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [21]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][22] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [22]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][23] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [23]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][24] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [24]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][25] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [25]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][26] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [26]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][27] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [27]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][28] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [28]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][29] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [29]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][2] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [2]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][30] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [30]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][31] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [31]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][3] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [3]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][4] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [4]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][5] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [5]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][6] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [6]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][7] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [7]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][8] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [8]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][9] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\CD[1].col_reg[2][31]_2 [9]),
        .Q(\IV_BKP_REGISTERS[1].bkp_1_reg[1][31]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][0] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [0]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][10] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [10]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][11] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [11]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][12] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [12]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][13] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [13]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][14] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [14]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][15] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [15]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][16] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [16]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][17] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [17]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][18] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [18]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][19] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [19]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][1] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [1]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][20] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [20]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][21] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [21]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][22] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [22]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][23] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [23]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][24] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [24]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][25] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [25]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][26] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [26]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][27] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [27]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][28] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [28]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][29] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [29]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][2] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [2]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][30] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [30]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][31] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [31]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][3] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [3]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][4] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [4]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][5] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [5]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][6] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [6]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][7] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [7]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][8] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [8]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].bkp_reg[1][9] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[1].bkp_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_4 [9]),
        .Q(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][0] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][10] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][11] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][12] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][13] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][14] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][15] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][16] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][17] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][18] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][19] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][1] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][20] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][21] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][22] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][23] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][24] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][25] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][26] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][27] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][28] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][29] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][2] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][30] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][31] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][3] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][4] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][5] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][6] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][7] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][8] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[1].iv_reg[1][9] 
       (.C(clk_i),
        .CE(iv_en[1]),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(\IV_BKP_REGISTERS[1].iv_reg[1][31]_0 [9]));
  LUT6 #(
    .INIT(64'hEEEEEEEBAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][24]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][24]_0 ),
        .I1(enable_i_8_sn_1),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][24]_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][24]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp_reg[1][24]_1 ),
        .I5(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ),
        .O(data_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][24]_i_5 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [24]),
        .I1(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [24]),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][24]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEBAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][25]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][25]_0 ),
        .I1(enable_i_9_sn_1),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][25]_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][25]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp_reg[1][25]_1 ),
        .I5(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ),
        .O(data_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][25]_i_5 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [25]),
        .I1(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [25]),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][25]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEBAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][26]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][26]_0 ),
        .I1(enable_i_10_sn_1),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][26]_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][26]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp_reg[1][26]_1 ),
        .I5(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ),
        .O(data_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][26]_i_5 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [26]),
        .I1(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [26]),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][26]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEBAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][27]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][27]_0 ),
        .I1(enable_i_11_sn_1),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][27]_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][27]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp_reg[1][27]_1 ),
        .I5(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ),
        .O(data_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][27]_i_5 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [27]),
        .I1(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [27]),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEBAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][29]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][29]_0 ),
        .I1(enable_i_13_sn_1),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][29]_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][29]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp_reg[1][29]_1 ),
        .I5(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ),
        .O(data_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][29]_i_5 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [29]),
        .I1(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [29]),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][29]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEBAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][30]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][30]_0 ),
        .I1(enable_i_14_sn_1),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][30]_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][30]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp_reg[1][30]_1 ),
        .I5(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ),
        .O(data_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][30]_i_5 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [30]),
        .I1(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [30]),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][30]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEBAAAAAAAA)) 
    \IV_BKP_REGISTERS[2].bkp[2][31]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_2 ),
        .I1(enable_i_15_sn_1),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_0 ),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][31]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_3 ),
        .I5(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ),
        .O(data_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][31]_i_5 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [31]),
        .I1(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [31]),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ),
        .O(\IV_BKP_REGISTERS[2].bkp[2][31]_i_5_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][0] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [0]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][10] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [10]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][11] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [11]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][12] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [12]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][13] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [13]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][14] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [14]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][15] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [15]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][16] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [16]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][17] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [17]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][18] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [18]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][19] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [19]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][1] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [1]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][20] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [20]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][21] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [21]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][22] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [22]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][23] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [23]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][24] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [24]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][25] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [25]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][26] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [26]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][27] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [27]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][28] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [28]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][29] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [29]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][2] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [2]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][30] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [30]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][31] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [31]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][3] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [3]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][4] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [4]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][5] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [5]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][6] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [6]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][7] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [7]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][8] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [8]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][9] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\CD[2].col_reg[1][31]_2 [9]),
        .Q(\IV_BKP_REGISTERS[2].bkp_1_reg[2][31]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][0] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [0]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][10] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [10]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][11] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [11]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][12] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [12]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][13] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [13]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][14] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [14]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][15] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [15]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][16] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [16]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][17] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [17]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][18] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [18]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][19] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [19]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][1] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [1]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][20] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [20]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][21] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [21]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][22] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [22]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][23] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [23]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][24] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [24]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][25] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [25]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][26] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [26]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][27] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [27]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][28] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [28]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][29] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [29]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][2] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [2]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][30] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [30]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][31] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [31]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][3] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [3]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][4] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [4]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][5] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [5]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][6] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [6]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][7] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [7]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][8] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [8]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].bkp_reg[2][9] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[2].bkp_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [9]),
        .Q(\IV_BKP_REGISTERS[2].bkp_reg[2]_13 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][0] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[0]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][10] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][11] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][12] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[12]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][13] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[13]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][14] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[14]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][15] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[15]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][16] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[16]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][17] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[17]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][18] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[18]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][19] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[19]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][1] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][20] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[20]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][21] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[21]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][22] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[22]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][23] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[23]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][24] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[24]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][25] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[25]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][26] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[26]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][27] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[27]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][28] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[28]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][29] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[29]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][2] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][30] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[30]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][31] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[31]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][3] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[3]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][4] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][5] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][6] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][7] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[7]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][8] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[2].iv_reg[2][9] 
       (.C(clk_i),
        .CE(iv_en[2]),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(\IV_BKP_REGISTERS[2].iv_reg[2][31]_0 [9]));
  LUT6 #(
    .INIT(64'hEEEEEEEBAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][14]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][14]_0 ),
        .I1(enable_i_30_sn_1),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][14]_0 ),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][14]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][14]_1 ),
        .I5(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ),
        .O(data_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \IV_BKP_REGISTERS[3].bkp[3][14]_i_5 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [14]),
        .I1(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [14]),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][14]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEBAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][15]_i_4 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][15]_0 ),
        .I1(enable_i_31_sn_1),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][15]_0 ),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][15]_i_7_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][15]_1 ),
        .I5(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ),
        .O(data_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \IV_BKP_REGISTERS[3].bkp[3][15]_i_7 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [15]),
        .I1(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [15]),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEBAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][8]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][8]_0 ),
        .I1(enable_i_24_sn_1),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][8]_0 ),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][8]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][8]_1 ),
        .I5(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ),
        .O(data_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \IV_BKP_REGISTERS[3].bkp[3][8]_i_5 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [8]),
        .I1(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [8]),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEBAAAAAAAA)) 
    \IV_BKP_REGISTERS[3].bkp[3][9]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][9]_0 ),
        .I1(enable_i_25_sn_1),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][9]_0 ),
        .I3(\IV_BKP_REGISTERS[3].bkp[3][9]_i_5_n_0 ),
        .I4(\IV_BKP_REGISTERS[0].bkp_reg[0][9]_1 ),
        .I5(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_1 ),
        .O(data_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \IV_BKP_REGISTERS[3].bkp[3][9]_i_5 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31]_0 [9]),
        .I1(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_0 ),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][31]_0 [9]),
        .I3(\IV_BKP_REGISTERS[2].bkp[2][31]_i_2_1 ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][9]_i_5_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][0] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [0]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][10] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [10]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][11] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [11]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][12] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [12]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][13] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [13]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][14] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [14]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][15] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [15]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][16] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [16]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][17] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [17]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][18] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [18]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][19] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [19]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][1] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [1]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][20] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [20]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][21] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [21]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][22] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [22]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][23] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [23]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][24] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [24]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][25] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [25]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][26] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [26]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][27] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [27]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][28] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [28]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][29] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [29]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][2] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [2]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][30] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [30]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][31] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [31]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][3] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [3]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][4] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [4]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][5] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [5]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][6] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [6]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][7] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [7]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][8] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [8]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][9] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\CD[3].col_reg[0][31]_2 [9]),
        .Q(\IV_BKP_REGISTERS[3].bkp_1_reg[3][31]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][0] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [0]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][10] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [10]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][11] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [11]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][12] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [12]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][13] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [13]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][14] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [14]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][15] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [15]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][16] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [16]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][17] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [17]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][18] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [18]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][19] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [19]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][1] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [1]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][20] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [20]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][21] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [21]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][22] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [22]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][23] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [23]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][24] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [24]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][25] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [25]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][26] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [26]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][27] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [27]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][28] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [28]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][29] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [29]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][2] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [2]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][30] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [30]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][31] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [31]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][3] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [3]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][4] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [4]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][5] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [5]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][6] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [6]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][7] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [7]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][8] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [8]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].bkp_reg[3][9] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].bkp_reg[3][0]_1 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].bkp_reg[3][31]_1 [9]),
        .Q(\IV_BKP_REGISTERS[3].bkp_reg[3]_11 [9]));
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT4 #(
    .INIT(16'h0080)) 
    \IV_BKP_REGISTERS[3].iv[3][31]_i_3 
       (.I0(enable_i[6]),
        .I1(enable_i[5]),
        .I2(enable_i[4]),
        .I3(enable_i[0]),
        .O(enable_i_6_sn_1));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][0] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [0]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][10] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [10]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][11] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [11]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][12] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [12]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][13] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [13]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][14] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [14]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][15] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [15]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][16] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [16]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [12]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2 
       (.CI(\IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_0 ),
        .CI_TOP(1'b0),
        .CO({\IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_0 ,\IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_1 ,\IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_2 ,\IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_3 ,\IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_4 ,\IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_5 ,\IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_6 ,\IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][16]_2 ),
        .S(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [12:5]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][17] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [17]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][18] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [18]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][19] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [19]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][1] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [1]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3]_4 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][20] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [20]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][21] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [21]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][22] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [22]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][23] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [23]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][24] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [24]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [20]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2 
       (.CI(\IV_BKP_REGISTERS[3].iv_reg[3][16]_i_2_n_0 ),
        .CI_TOP(1'b0),
        .CO({\IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_0 ,\IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_1 ,\IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_2 ,\IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_3 ,\IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_4 ,\IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_5 ,\IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_6 ,\IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][24]_2 ),
        .S(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [20:13]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][25] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [25]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][26] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [26]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][27] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [27]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][28] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [28]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][29] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [29]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][2] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [2]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3]_4 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][30] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [30]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][31] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [31]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [27]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7 
       (.CI(\IV_BKP_REGISTERS[3].iv_reg[3][24]_i_2_n_0 ),
        .CI_TOP(1'b0),
        .CO({\NLW_IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_CO_UNCONNECTED [7:6],\IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_n_2 ,\IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_n_3 ,\IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_n_4 ,\IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_n_5 ,\IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_n_6 ,\IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O({\NLW_IV_BKP_REGISTERS[3].iv_reg[3][31]_i_7_O_UNCONNECTED [7],O}),
        .S({1'b0,\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [27:21]}));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][3] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [3]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3]_4 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][4] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [4]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][5] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [5]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3]_4 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][6] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [6]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][7] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [7]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][8] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [8]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [4]));
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2 
       (.CI(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [0]),
        .CI_TOP(1'b0),
        .CO({\IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_0 ,\IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_1 ,\IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_2 ,\IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_3 ,\IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_4 ,\IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_5 ,\IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_6 ,\IV_BKP_REGISTERS[3].iv_reg[3][8]_i_2_n_7 }),
        .DI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .O(\IV_BKP_REGISTERS[3].iv_reg[3][0]_1 ),
        .S({\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [4:2],\IV_BKP_REGISTERS[3].iv_reg[3]_4 [5],\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [1],\IV_BKP_REGISTERS[3].iv_reg[3]_4 [3:1]}));
  FDCE #(
    .INIT(1'b0)) 
    \IV_BKP_REGISTERS[3].iv_reg[3][9] 
       (.C(clk_i),
        .CE(\IV_BKP_REGISTERS[3].iv_reg[3][0]_2 ),
        .CLR(rst_i),
        .D(\IV_BKP_REGISTERS[3].iv_reg[3][31]_3 [9]),
        .Q(\IV_BKP_REGISTERS[3].iv_reg[3][31]_0 [5]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][0]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [0]),
        .I2(enable_i[0]),
        .I3(key_sel_mux),
        .I4(key_in[32]),
        .I5(key_in[0]),
        .O(\KR[0].key[3][0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][10]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [10]),
        .I2(enable_i[10]),
        .I3(key_sel_mux),
        .I4(key_in[42]),
        .I5(key_in[10]),
        .O(\KR[0].key[3][10]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][11]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [11]),
        .I2(enable_i[11]),
        .I3(key_sel_mux),
        .I4(key_in[43]),
        .I5(key_in[11]),
        .O(\KR[0].key[3][11]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][12]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [12]),
        .I2(enable_i[12]),
        .I3(key_sel_mux),
        .I4(key_in[44]),
        .I5(key_in[12]),
        .O(\KR[0].key[3][12]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][13]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [13]),
        .I2(enable_i[13]),
        .I3(key_sel_mux),
        .I4(key_in[45]),
        .I5(key_in[13]),
        .O(\KR[0].key[3][13]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][14]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [14]),
        .I2(enable_i[14]),
        .I3(key_sel_mux),
        .I4(key_in[46]),
        .I5(key_in[14]),
        .O(\KR[0].key[3][14]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][15]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [15]),
        .I2(enable_i[15]),
        .I3(key_sel_mux),
        .I4(key_in[47]),
        .I5(key_in[15]),
        .O(\KR[0].key[3][15]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][16]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [16]),
        .I2(enable_i[16]),
        .I3(key_sel_mux),
        .I4(key_in[48]),
        .I5(key_in[16]),
        .O(\KR[0].key[3][16]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][17]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [17]),
        .I2(enable_i[17]),
        .I3(key_sel_mux),
        .I4(key_in[49]),
        .I5(key_in[17]),
        .O(\KR[0].key[3][17]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][18]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [18]),
        .I2(enable_i[18]),
        .I3(key_sel_mux),
        .I4(key_in[50]),
        .I5(key_in[18]),
        .O(\KR[0].key[3][18]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][19]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [19]),
        .I2(enable_i[19]),
        .I3(key_sel_mux),
        .I4(key_in[51]),
        .I5(key_in[19]),
        .O(\KR[0].key[3][19]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][1]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [1]),
        .I2(enable_i[1]),
        .I3(key_sel_mux),
        .I4(key_in[33]),
        .I5(key_in[1]),
        .O(\KR[0].key[3][1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][20]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [20]),
        .I2(enable_i[20]),
        .I3(key_sel_mux),
        .I4(key_in[52]),
        .I5(key_in[20]),
        .O(\KR[0].key[3][20]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][21]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [21]),
        .I2(enable_i[21]),
        .I3(key_sel_mux),
        .I4(key_in[53]),
        .I5(key_in[21]),
        .O(\KR[0].key[3][21]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][22]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [22]),
        .I2(enable_i[22]),
        .I3(key_sel_mux),
        .I4(key_in[54]),
        .I5(key_in[22]),
        .O(\KR[0].key[3][22]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][23]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [23]),
        .I2(enable_i[23]),
        .I3(key_sel_mux),
        .I4(key_in[55]),
        .I5(key_in[23]),
        .O(\KR[0].key[3][23]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][24]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [24]),
        .I2(enable_i[24]),
        .I3(key_sel_mux),
        .I4(key_in[56]),
        .I5(key_in[24]),
        .O(\KR[0].key[3][24]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][25]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [25]),
        .I2(enable_i[25]),
        .I3(key_sel_mux),
        .I4(key_in[57]),
        .I5(key_in[25]),
        .O(\KR[0].key[3][25]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][26]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [26]),
        .I2(enable_i[26]),
        .I3(key_sel_mux),
        .I4(key_in[58]),
        .I5(key_in[26]),
        .O(\KR[0].key[3][26]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][27]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [27]),
        .I2(enable_i[27]),
        .I3(key_sel_mux),
        .I4(key_in[59]),
        .I5(key_in[27]),
        .O(\KR[0].key[3][27]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][28]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [28]),
        .I2(enable_i[28]),
        .I3(key_sel_mux),
        .I4(key_in[60]),
        .I5(key_in[28]),
        .O(\KR[0].key[3][28]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][29]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [29]),
        .I2(enable_i[29]),
        .I3(key_sel_mux),
        .I4(key_in[61]),
        .I5(key_in[29]),
        .O(\KR[0].key[3][29]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][2]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [2]),
        .I2(enable_i[2]),
        .I3(key_sel_mux),
        .I4(key_in[34]),
        .I5(key_in[2]),
        .O(\KR[0].key[3][2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][30]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [30]),
        .I2(enable_i[30]),
        .I3(key_sel_mux),
        .I4(key_in[62]),
        .I5(key_in[30]),
        .O(\KR[0].key[3][30]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][31]_i_2 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [31]),
        .I2(enable_i[31]),
        .I3(key_sel_mux),
        .I4(key_in[63]),
        .I5(key_in[31]),
        .O(\KR[0].key[3][31]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][3]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [3]),
        .I2(enable_i[3]),
        .I3(key_sel_mux),
        .I4(key_in[35]),
        .I5(key_in[3]),
        .O(\KR[0].key[3][3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][4]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [4]),
        .I2(enable_i[4]),
        .I3(key_sel_mux),
        .I4(key_in[36]),
        .I5(key_in[4]),
        .O(\KR[0].key[3][4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][5]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [5]),
        .I2(enable_i[5]),
        .I3(key_sel_mux),
        .I4(key_in[37]),
        .I5(key_in[5]),
        .O(\KR[0].key[3][5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][6]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [6]),
        .I2(enable_i[6]),
        .I3(key_sel_mux),
        .I4(key_in[38]),
        .I5(key_in[6]),
        .O(\KR[0].key[3][6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][7]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [7]),
        .I2(enable_i[7]),
        .I3(key_sel_mux),
        .I4(key_in[39]),
        .I5(key_in[7]),
        .O(\KR[0].key[3][7]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][8]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [8]),
        .I2(enable_i[8]),
        .I3(key_sel_mux),
        .I4(key_in[40]),
        .I5(key_in[8]),
        .O(\KR[0].key[3][8]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[0].key[3][9]_i_1 
       (.I0(key_en[2]),
        .I1(\KR[0].key_host_reg[3]_0 [9]),
        .I2(enable_i[9]),
        .I3(key_sel_mux),
        .I4(key_in[41]),
        .I5(key_in[9]),
        .O(\KR[0].key[3][9]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair236" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][0]_i_1 
       (.I0(key_in[0]),
        .I1(key_derivation_en),
        .I2(enable_i[0]),
        .O(\KR[0].key_host[3][0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][10]_i_1 
       (.I0(key_in[10]),
        .I1(key_derivation_en),
        .I2(enable_i[10]),
        .O(\KR[0].key_host[3][10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][11]_i_1 
       (.I0(key_in[11]),
        .I1(key_derivation_en),
        .I2(enable_i[11]),
        .O(\KR[0].key_host[3][11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][12]_i_1 
       (.I0(key_in[12]),
        .I1(key_derivation_en),
        .I2(enable_i[12]),
        .O(\KR[0].key_host[3][12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][13]_i_1 
       (.I0(key_in[13]),
        .I1(key_derivation_en),
        .I2(enable_i[13]),
        .O(\KR[0].key_host[3][13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][14]_i_1 
       (.I0(key_in[14]),
        .I1(key_derivation_en),
        .I2(enable_i[14]),
        .O(\KR[0].key_host[3][14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][15]_i_1 
       (.I0(key_in[15]),
        .I1(key_derivation_en),
        .I2(enable_i[15]),
        .O(\KR[0].key_host[3][15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair237" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][16]_i_1 
       (.I0(key_in[16]),
        .I1(key_derivation_en),
        .I2(enable_i[16]),
        .O(\KR[0].key_host[3][16]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][17]_i_1 
       (.I0(key_in[17]),
        .I1(key_derivation_en),
        .I2(enable_i[17]),
        .O(\KR[0].key_host[3][17]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][18]_i_1 
       (.I0(key_in[18]),
        .I1(key_derivation_en),
        .I2(enable_i[18]),
        .O(\KR[0].key_host[3][18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair243" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][19]_i_1 
       (.I0(key_in[19]),
        .I1(key_derivation_en),
        .I2(enable_i[19]),
        .O(\KR[0].key_host[3][19]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][1]_i_1 
       (.I0(key_in[1]),
        .I1(key_derivation_en),
        .I2(enable_i[1]),
        .O(\KR[0].key_host[3][1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair245" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][20]_i_1 
       (.I0(key_in[20]),
        .I1(key_derivation_en),
        .I2(enable_i[20]),
        .O(\KR[0].key_host[3][20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair247" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][21]_i_1 
       (.I0(key_in[21]),
        .I1(key_derivation_en),
        .I2(enable_i[21]),
        .O(\KR[0].key_host[3][21]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair267" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][22]_i_1 
       (.I0(key_in[22]),
        .I1(key_derivation_en),
        .I2(enable_i[22]),
        .O(\KR[0].key_host[3][22]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair249" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][23]_i_1 
       (.I0(key_in[23]),
        .I1(key_derivation_en),
        .I2(enable_i[23]),
        .O(\KR[0].key_host[3][23]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair251" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][24]_i_1 
       (.I0(key_in[24]),
        .I1(key_derivation_en),
        .I2(enable_i[24]),
        .O(\KR[0].key_host[3][24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair253" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][25]_i_1 
       (.I0(key_in[25]),
        .I1(key_derivation_en),
        .I2(enable_i[25]),
        .O(\KR[0].key_host[3][25]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair255" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][26]_i_1 
       (.I0(key_in[26]),
        .I1(key_derivation_en),
        .I2(enable_i[26]),
        .O(\KR[0].key_host[3][26]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair257" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][27]_i_1 
       (.I0(key_in[27]),
        .I1(key_derivation_en),
        .I2(enable_i[27]),
        .O(\KR[0].key_host[3][27]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair259" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][28]_i_1 
       (.I0(key_in[28]),
        .I1(key_derivation_en),
        .I2(enable_i[28]),
        .O(\KR[0].key_host[3][28]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair261" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][29]_i_1 
       (.I0(key_in[29]),
        .I1(key_derivation_en),
        .I2(enable_i[29]),
        .O(\KR[0].key_host[3][29]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][2]_i_1 
       (.I0(key_in[2]),
        .I1(key_derivation_en),
        .I2(enable_i[2]),
        .O(\KR[0].key_host[3][2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair263" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][30]_i_1 
       (.I0(key_in[30]),
        .I1(key_derivation_en),
        .I2(enable_i[30]),
        .O(\KR[0].key_host[3][30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair265" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][31]_i_2 
       (.I0(key_in[31]),
        .I1(key_derivation_en),
        .I2(enable_i[31]),
        .O(\KR[0].key_host[3][31]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][3]_i_1 
       (.I0(key_in[3]),
        .I1(key_derivation_en),
        .I2(enable_i[3]),
        .O(\KR[0].key_host[3][3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][4]_i_1 
       (.I0(key_in[4]),
        .I1(key_derivation_en),
        .I2(enable_i[4]),
        .O(\KR[0].key_host[3][4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][5]_i_1 
       (.I0(key_in[5]),
        .I1(key_derivation_en),
        .I2(enable_i[5]),
        .O(\KR[0].key_host[3][5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][6]_i_1 
       (.I0(key_in[6]),
        .I1(key_derivation_en),
        .I2(enable_i[6]),
        .O(\KR[0].key_host[3][6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][7]_i_1 
       (.I0(key_in[7]),
        .I1(key_derivation_en),
        .I2(enable_i[7]),
        .O(\KR[0].key_host[3][7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][8]_i_1 
       (.I0(key_in[8]),
        .I1(key_derivation_en),
        .I2(enable_i[8]),
        .O(\KR[0].key_host[3][8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[0].key_host[3][9]_i_1 
       (.I0(key_in[9]),
        .I1(key_derivation_en),
        .I2(enable_i[9]),
        .O(\KR[0].key_host[3][9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][0] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][0]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][10] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][10]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][11] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][11]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][12] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][12]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][13] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][13]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][14] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][14]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][15] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][15]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][16] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][16]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][17] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][17]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][18] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][18]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][19] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][19]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][1] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][1]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][20] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][20]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][21] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][21]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][22] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][22]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][23] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][23]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][24] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][24]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][25] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][25]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][26] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][26]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][27] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][27]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][28] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][28]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][29] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][29]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][2] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][2]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][30] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][30]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][31] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][31]_i_2_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][3] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][3]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][4] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][4]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][5] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][5]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][6] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][6]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][7] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][7]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][8] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][8]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_host_reg[3][9] 
       (.C(clk_i),
        .CE(\KR[0].key_host_reg[3][0]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key_host[3][9]_i_1_n_0 ),
        .Q(\KR[0].key_host_reg[3]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][0] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][0]_i_1_n_0 ),
        .Q(key_in[0]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][10] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][10]_i_1_n_0 ),
        .Q(key_in[10]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][11] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][11]_i_1_n_0 ),
        .Q(key_in[11]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][12] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][12]_i_1_n_0 ),
        .Q(key_in[12]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][13] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][13]_i_1_n_0 ),
        .Q(key_in[13]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][14] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][14]_i_1_n_0 ),
        .Q(key_in[14]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][15] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][15]_i_1_n_0 ),
        .Q(key_in[15]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][16] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][16]_i_1_n_0 ),
        .Q(key_in[16]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][17] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][17]_i_1_n_0 ),
        .Q(key_in[17]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][18] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][18]_i_1_n_0 ),
        .Q(key_in[18]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][19] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][19]_i_1_n_0 ),
        .Q(key_in[19]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][1] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][1]_i_1_n_0 ),
        .Q(key_in[1]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][20] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][20]_i_1_n_0 ),
        .Q(key_in[20]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][21] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][21]_i_1_n_0 ),
        .Q(key_in[21]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][22] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][22]_i_1_n_0 ),
        .Q(key_in[22]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][23] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][23]_i_1_n_0 ),
        .Q(key_in[23]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][24] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][24]_i_1_n_0 ),
        .Q(key_in[24]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][25] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][25]_i_1_n_0 ),
        .Q(key_in[25]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][26] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][26]_i_1_n_0 ),
        .Q(key_in[26]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][27] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][27]_i_1_n_0 ),
        .Q(key_in[27]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][28] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][28]_i_1_n_0 ),
        .Q(key_in[28]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][29] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][29]_i_1_n_0 ),
        .Q(key_in[29]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][2] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][2]_i_1_n_0 ),
        .Q(key_in[2]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][30] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][30]_i_1_n_0 ),
        .Q(key_in[30]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][31] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][31]_i_2_n_0 ),
        .Q(key_in[31]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][3] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][3]_i_1_n_0 ),
        .Q(key_in[3]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][4] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][4]_i_1_n_0 ),
        .Q(key_in[4]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][5] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][5]_i_1_n_0 ),
        .Q(key_in[5]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][6] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][6]_i_1_n_0 ),
        .Q(key_in[6]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][7] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][7]_i_1_n_0 ),
        .Q(key_in[7]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][8] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][8]_i_1_n_0 ),
        .Q(key_in[8]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[0].key_reg[3][9] 
       (.C(clk_i),
        .CE(\KR[0].key_reg[3][31]_0 ),
        .CLR(rst_i),
        .D(\KR[0].key[3][9]_i_1_n_0 ),
        .Q(key_in[9]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][0]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [0]),
        .I2(enable_i[0]),
        .I3(key_sel_mux),
        .I4(key_in[64]),
        .I5(key_in[32]),
        .O(\KR[1].key[2][0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][10]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [10]),
        .I2(enable_i[10]),
        .I3(key_sel_mux),
        .I4(key_in[74]),
        .I5(key_in[42]),
        .O(\KR[1].key[2][10]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][11]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [11]),
        .I2(enable_i[11]),
        .I3(key_sel_mux),
        .I4(key_in[75]),
        .I5(key_in[43]),
        .O(\KR[1].key[2][11]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][12]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [12]),
        .I2(enable_i[12]),
        .I3(key_sel_mux),
        .I4(key_in[76]),
        .I5(key_in[44]),
        .O(\KR[1].key[2][12]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][13]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [13]),
        .I2(enable_i[13]),
        .I3(key_sel_mux),
        .I4(key_in[77]),
        .I5(key_in[45]),
        .O(\KR[1].key[2][13]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][14]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [14]),
        .I2(enable_i[14]),
        .I3(key_sel_mux),
        .I4(key_in[78]),
        .I5(key_in[46]),
        .O(\KR[1].key[2][14]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][15]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [15]),
        .I2(enable_i[15]),
        .I3(key_sel_mux),
        .I4(key_in[79]),
        .I5(key_in[47]),
        .O(\KR[1].key[2][15]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][16]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [16]),
        .I2(enable_i[16]),
        .I3(key_sel_mux),
        .I4(key_in[80]),
        .I5(key_in[48]),
        .O(\KR[1].key[2][16]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][17]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [17]),
        .I2(enable_i[17]),
        .I3(key_sel_mux),
        .I4(key_in[81]),
        .I5(key_in[49]),
        .O(\KR[1].key[2][17]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][18]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [18]),
        .I2(enable_i[18]),
        .I3(key_sel_mux),
        .I4(key_in[82]),
        .I5(key_in[50]),
        .O(\KR[1].key[2][18]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][19]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [19]),
        .I2(enable_i[19]),
        .I3(key_sel_mux),
        .I4(key_in[83]),
        .I5(key_in[51]),
        .O(\KR[1].key[2][19]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][1]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [1]),
        .I2(enable_i[1]),
        .I3(key_sel_mux),
        .I4(key_in[65]),
        .I5(key_in[33]),
        .O(\KR[1].key[2][1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][20]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [20]),
        .I2(enable_i[20]),
        .I3(key_sel_mux),
        .I4(key_in[84]),
        .I5(key_in[52]),
        .O(\KR[1].key[2][20]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][21]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [21]),
        .I2(enable_i[21]),
        .I3(key_sel_mux),
        .I4(key_in[85]),
        .I5(key_in[53]),
        .O(\KR[1].key[2][21]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][22]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [22]),
        .I2(enable_i[22]),
        .I3(key_sel_mux),
        .I4(key_in[86]),
        .I5(key_in[54]),
        .O(\KR[1].key[2][22]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][23]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [23]),
        .I2(enable_i[23]),
        .I3(key_sel_mux),
        .I4(key_in[87]),
        .I5(key_in[55]),
        .O(\KR[1].key[2][23]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][24]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [24]),
        .I2(enable_i[24]),
        .I3(key_sel_mux),
        .I4(key_in[88]),
        .I5(key_in[56]),
        .O(\KR[1].key[2][24]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][25]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [25]),
        .I2(enable_i[25]),
        .I3(key_sel_mux),
        .I4(key_in[89]),
        .I5(key_in[57]),
        .O(\KR[1].key[2][25]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][26]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [26]),
        .I2(enable_i[26]),
        .I3(key_sel_mux),
        .I4(key_in[90]),
        .I5(key_in[58]),
        .O(\KR[1].key[2][26]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][27]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [27]),
        .I2(enable_i[27]),
        .I3(key_sel_mux),
        .I4(key_in[91]),
        .I5(key_in[59]),
        .O(\KR[1].key[2][27]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][28]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [28]),
        .I2(enable_i[28]),
        .I3(key_sel_mux),
        .I4(key_in[92]),
        .I5(key_in[60]),
        .O(\KR[1].key[2][28]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][29]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [29]),
        .I2(enable_i[29]),
        .I3(key_sel_mux),
        .I4(key_in[93]),
        .I5(key_in[61]),
        .O(\KR[1].key[2][29]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][2]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [2]),
        .I2(enable_i[2]),
        .I3(key_sel_mux),
        .I4(key_in[66]),
        .I5(key_in[34]),
        .O(\KR[1].key[2][2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][30]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [30]),
        .I2(enable_i[30]),
        .I3(key_sel_mux),
        .I4(key_in[94]),
        .I5(key_in[62]),
        .O(\KR[1].key[2][30]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][31]_i_2 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [31]),
        .I2(enable_i[31]),
        .I3(key_sel_mux),
        .I4(key_in[95]),
        .I5(key_in[63]),
        .O(\KR[1].key[2][31]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][3]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [3]),
        .I2(enable_i[3]),
        .I3(key_sel_mux),
        .I4(key_in[67]),
        .I5(key_in[35]),
        .O(\KR[1].key[2][3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][4]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [4]),
        .I2(enable_i[4]),
        .I3(key_sel_mux),
        .I4(key_in[68]),
        .I5(key_in[36]),
        .O(\KR[1].key[2][4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][5]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [5]),
        .I2(enable_i[5]),
        .I3(key_sel_mux),
        .I4(key_in[69]),
        .I5(key_in[37]),
        .O(\KR[1].key[2][5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][6]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [6]),
        .I2(enable_i[6]),
        .I3(key_sel_mux),
        .I4(key_in[70]),
        .I5(key_in[38]),
        .O(\KR[1].key[2][6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][7]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [7]),
        .I2(enable_i[7]),
        .I3(key_sel_mux),
        .I4(key_in[71]),
        .I5(key_in[39]),
        .O(\KR[1].key[2][7]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][8]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [8]),
        .I2(enable_i[8]),
        .I3(key_sel_mux),
        .I4(key_in[72]),
        .I5(key_in[40]),
        .O(\KR[1].key[2][8]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[1].key[2][9]_i_1 
       (.I0(key_en[1]),
        .I1(\KR[1].key_host_reg[2]_1 [9]),
        .I2(enable_i[9]),
        .I3(key_sel_mux),
        .I4(key_in[73]),
        .I5(key_in[41]),
        .O(\KR[1].key[2][9]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair236" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][0]_i_1 
       (.I0(key_in[32]),
        .I1(key_derivation_en),
        .I2(enable_i[0]),
        .O(\KR[1].key_host[2][0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][10]_i_1 
       (.I0(key_in[42]),
        .I1(key_derivation_en),
        .I2(enable_i[10]),
        .O(\KR[1].key_host[2][10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][11]_i_1 
       (.I0(key_in[43]),
        .I1(key_derivation_en),
        .I2(enable_i[11]),
        .O(\KR[1].key_host[2][11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][12]_i_1 
       (.I0(key_in[44]),
        .I1(key_derivation_en),
        .I2(enable_i[12]),
        .O(\KR[1].key_host[2][12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][13]_i_1 
       (.I0(key_in[45]),
        .I1(key_derivation_en),
        .I2(enable_i[13]),
        .O(\KR[1].key_host[2][13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][14]_i_1 
       (.I0(key_in[46]),
        .I1(key_derivation_en),
        .I2(enable_i[14]),
        .O(\KR[1].key_host[2][14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][15]_i_1 
       (.I0(key_in[47]),
        .I1(key_derivation_en),
        .I2(enable_i[15]),
        .O(\KR[1].key_host[2][15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][16]_i_1 
       (.I0(key_in[48]),
        .I1(key_derivation_en),
        .I2(enable_i[16]),
        .O(\KR[1].key_host[2][16]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair240" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][17]_i_1 
       (.I0(key_in[49]),
        .I1(key_derivation_en),
        .I2(enable_i[17]),
        .O(\KR[1].key_host[2][17]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][18]_i_1 
       (.I0(key_in[50]),
        .I1(key_derivation_en),
        .I2(enable_i[18]),
        .O(\KR[1].key_host[2][18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair244" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][19]_i_1 
       (.I0(key_in[51]),
        .I1(key_derivation_en),
        .I2(enable_i[19]),
        .O(\KR[1].key_host[2][19]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][1]_i_1 
       (.I0(key_in[33]),
        .I1(key_derivation_en),
        .I2(enable_i[1]),
        .O(\KR[1].key_host[2][1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair246" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][20]_i_1 
       (.I0(key_in[52]),
        .I1(key_derivation_en),
        .I2(enable_i[20]),
        .O(\KR[1].key_host[2][20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair248" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][21]_i_1 
       (.I0(key_in[53]),
        .I1(key_derivation_en),
        .I2(enable_i[21]),
        .O(\KR[1].key_host[2][21]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair268" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][22]_i_1 
       (.I0(key_in[54]),
        .I1(key_derivation_en),
        .I2(enable_i[22]),
        .O(\KR[1].key_host[2][22]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair250" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][23]_i_1 
       (.I0(key_in[55]),
        .I1(key_derivation_en),
        .I2(enable_i[23]),
        .O(\KR[1].key_host[2][23]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair252" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][24]_i_1 
       (.I0(key_in[56]),
        .I1(key_derivation_en),
        .I2(enable_i[24]),
        .O(\KR[1].key_host[2][24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair254" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][25]_i_1 
       (.I0(key_in[57]),
        .I1(key_derivation_en),
        .I2(enable_i[25]),
        .O(\KR[1].key_host[2][25]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair256" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][26]_i_1 
       (.I0(key_in[58]),
        .I1(key_derivation_en),
        .I2(enable_i[26]),
        .O(\KR[1].key_host[2][26]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair258" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][27]_i_1 
       (.I0(key_in[59]),
        .I1(key_derivation_en),
        .I2(enable_i[27]),
        .O(\KR[1].key_host[2][27]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair260" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][28]_i_1 
       (.I0(key_in[60]),
        .I1(key_derivation_en),
        .I2(enable_i[28]),
        .O(\KR[1].key_host[2][28]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair262" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][29]_i_1 
       (.I0(key_in[61]),
        .I1(key_derivation_en),
        .I2(enable_i[29]),
        .O(\KR[1].key_host[2][29]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][2]_i_1 
       (.I0(key_in[34]),
        .I1(key_derivation_en),
        .I2(enable_i[2]),
        .O(\KR[1].key_host[2][2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair264" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][30]_i_1 
       (.I0(key_in[62]),
        .I1(key_derivation_en),
        .I2(enable_i[30]),
        .O(\KR[1].key_host[2][30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair266" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][31]_i_2 
       (.I0(key_in[63]),
        .I1(key_derivation_en),
        .I2(enable_i[31]),
        .O(\KR[1].key_host[2][31]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hF7)) 
    \KR[1].key_host[2][31]_i_4 
       (.I0(enable_i[6]),
        .I1(enable_i[5]),
        .I2(enable_i[3]),
        .O(\enable_i[6]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][3]_i_1 
       (.I0(key_in[35]),
        .I1(key_derivation_en),
        .I2(enable_i[3]),
        .O(\KR[1].key_host[2][3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][4]_i_1 
       (.I0(key_in[36]),
        .I1(key_derivation_en),
        .I2(enable_i[4]),
        .O(\KR[1].key_host[2][4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][5]_i_1 
       (.I0(key_in[37]),
        .I1(key_derivation_en),
        .I2(enable_i[5]),
        .O(\KR[1].key_host[2][5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][6]_i_1 
       (.I0(key_in[38]),
        .I1(key_derivation_en),
        .I2(enable_i[6]),
        .O(\KR[1].key_host[2][6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][7]_i_1 
       (.I0(key_in[39]),
        .I1(key_derivation_en),
        .I2(enable_i[7]),
        .O(\KR[1].key_host[2][7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][8]_i_1 
       (.I0(key_in[40]),
        .I1(key_derivation_en),
        .I2(enable_i[8]),
        .O(\KR[1].key_host[2][8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[1].key_host[2][9]_i_1 
       (.I0(key_in[41]),
        .I1(key_derivation_en),
        .I2(enable_i[9]),
        .O(\KR[1].key_host[2][9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][0] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][0]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][10] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][10]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][11] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][11]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][12] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][12]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][13] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][13]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][14] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][14]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][15] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][15]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][16] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][16]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][17] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][17]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][18] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][18]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][19] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][19]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][1] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][1]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][20] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][20]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][21] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][21]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][22] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][22]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][23] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][23]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][24] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][24]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][25] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][25]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][26] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][26]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][27] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][27]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][28] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][28]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][29] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][29]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][2] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][2]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][30] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][30]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][31] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][31]_i_2_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][3] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][3]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][4] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][4]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][5] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][5]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][6] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][6]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][7] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][7]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][8] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][8]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_host_reg[2][9] 
       (.C(clk_i),
        .CE(\KR[1].key_host_reg[2][0]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key_host[2][9]_i_1_n_0 ),
        .Q(\KR[1].key_host_reg[2]_1 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][0] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][0]_i_1_n_0 ),
        .Q(key_in[32]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][10] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][10]_i_1_n_0 ),
        .Q(key_in[42]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][11] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][11]_i_1_n_0 ),
        .Q(key_in[43]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][12] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][12]_i_1_n_0 ),
        .Q(key_in[44]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][13] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][13]_i_1_n_0 ),
        .Q(key_in[45]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][14] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][14]_i_1_n_0 ),
        .Q(key_in[46]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][15] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][15]_i_1_n_0 ),
        .Q(key_in[47]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][16] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][16]_i_1_n_0 ),
        .Q(key_in[48]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][17] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][17]_i_1_n_0 ),
        .Q(key_in[49]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][18] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][18]_i_1_n_0 ),
        .Q(key_in[50]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][19] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][19]_i_1_n_0 ),
        .Q(key_in[51]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][1] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][1]_i_1_n_0 ),
        .Q(key_in[33]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][20] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][20]_i_1_n_0 ),
        .Q(key_in[52]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][21] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][21]_i_1_n_0 ),
        .Q(key_in[53]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][22] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][22]_i_1_n_0 ),
        .Q(key_in[54]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][23] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][23]_i_1_n_0 ),
        .Q(key_in[55]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][24] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][24]_i_1_n_0 ),
        .Q(key_in[56]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][25] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][25]_i_1_n_0 ),
        .Q(key_in[57]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][26] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][26]_i_1_n_0 ),
        .Q(key_in[58]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][27] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][27]_i_1_n_0 ),
        .Q(key_in[59]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][28] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][28]_i_1_n_0 ),
        .Q(key_in[60]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][29] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][29]_i_1_n_0 ),
        .Q(key_in[61]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][2] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][2]_i_1_n_0 ),
        .Q(key_in[34]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][30] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][30]_i_1_n_0 ),
        .Q(key_in[62]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][31] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][31]_i_2_n_0 ),
        .Q(key_in[63]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][3] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][3]_i_1_n_0 ),
        .Q(key_in[35]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][4] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][4]_i_1_n_0 ),
        .Q(key_in[36]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][5] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][5]_i_1_n_0 ),
        .Q(key_in[37]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][6] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][6]_i_1_n_0 ),
        .Q(key_in[38]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][7] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][7]_i_1_n_0 ),
        .Q(key_in[39]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][8] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][8]_i_1_n_0 ),
        .Q(key_in[40]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[1].key_reg[2][9] 
       (.C(clk_i),
        .CE(\KR[1].key_reg[2][31]_0 ),
        .CLR(rst_i),
        .D(\KR[1].key[2][9]_i_1_n_0 ),
        .Q(key_in[41]));
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT5 #(
    .INIT(32'h10080021)) 
    \KR[2].key[1][26]_i_4 
       (.I0(enc_dec_sbox),
        .I1(round_pp1[3]),
        .I2(round_pp1[1]),
        .I3(round_pp1[2]),
        .I4(round_pp1[0]),
        .O(\KEY_EXPANDER/rc [2]));
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT5 #(
    .INIT(32'h00211008)) 
    \KR[2].key[1][27]_i_4 
       (.I0(enc_dec_sbox),
        .I1(round_pp1[3]),
        .I2(round_pp1[1]),
        .I3(round_pp1[2]),
        .I4(round_pp1[0]),
        .O(\KEY_EXPANDER/rc [3]));
  (* SOFT_HLUTNM = "soft_lutpair235" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][0]_i_1 
       (.I0(key_in[64]),
        .I1(key_derivation_en),
        .I2(enable_i[0]),
        .O(\KR[2].key_host[1][0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][10]_i_1 
       (.I0(key_in[74]),
        .I1(key_derivation_en),
        .I2(enable_i[10]),
        .O(\KR[2].key_host[1][10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][11]_i_1 
       (.I0(key_in[75]),
        .I1(key_derivation_en),
        .I2(enable_i[11]),
        .O(\KR[2].key_host[1][11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][12]_i_1 
       (.I0(key_in[76]),
        .I1(key_derivation_en),
        .I2(enable_i[12]),
        .O(\KR[2].key_host[1][12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][13]_i_1 
       (.I0(key_in[77]),
        .I1(key_derivation_en),
        .I2(enable_i[13]),
        .O(\KR[2].key_host[1][13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][14]_i_1 
       (.I0(key_in[78]),
        .I1(key_derivation_en),
        .I2(enable_i[14]),
        .O(\KR[2].key_host[1][14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][15]_i_1 
       (.I0(key_in[79]),
        .I1(key_derivation_en),
        .I2(enable_i[15]),
        .O(\KR[2].key_host[1][15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][16]_i_1 
       (.I0(key_in[80]),
        .I1(key_derivation_en),
        .I2(enable_i[16]),
        .O(\KR[2].key_host[1][16]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair240" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][17]_i_1 
       (.I0(key_in[81]),
        .I1(key_derivation_en),
        .I2(enable_i[17]),
        .O(\KR[2].key_host[1][17]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][18]_i_1 
       (.I0(key_in[82]),
        .I1(key_derivation_en),
        .I2(enable_i[18]),
        .O(\KR[2].key_host[1][18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair244" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][19]_i_1 
       (.I0(key_in[83]),
        .I1(key_derivation_en),
        .I2(enable_i[19]),
        .O(\KR[2].key_host[1][19]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][1]_i_1 
       (.I0(key_in[65]),
        .I1(key_derivation_en),
        .I2(enable_i[1]),
        .O(\KR[2].key_host[1][1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair246" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][20]_i_1 
       (.I0(key_in[84]),
        .I1(key_derivation_en),
        .I2(enable_i[20]),
        .O(\KR[2].key_host[1][20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair248" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][21]_i_1 
       (.I0(key_in[85]),
        .I1(key_derivation_en),
        .I2(enable_i[21]),
        .O(\KR[2].key_host[1][21]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair268" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][22]_i_1 
       (.I0(key_in[86]),
        .I1(key_derivation_en),
        .I2(enable_i[22]),
        .O(\KR[2].key_host[1][22]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair250" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][23]_i_1 
       (.I0(key_in[87]),
        .I1(key_derivation_en),
        .I2(enable_i[23]),
        .O(\KR[2].key_host[1][23]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair252" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][24]_i_1 
       (.I0(key_in[88]),
        .I1(key_derivation_en),
        .I2(enable_i[24]),
        .O(\KR[2].key_host[1][24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair254" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][25]_i_1 
       (.I0(key_in[89]),
        .I1(key_derivation_en),
        .I2(enable_i[25]),
        .O(\KR[2].key_host[1][25]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair256" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][26]_i_1 
       (.I0(key_in[90]),
        .I1(key_derivation_en),
        .I2(enable_i[26]),
        .O(\KR[2].key_host[1][26]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair258" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][27]_i_1 
       (.I0(key_in[91]),
        .I1(key_derivation_en),
        .I2(enable_i[27]),
        .O(\KR[2].key_host[1][27]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair260" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][28]_i_1 
       (.I0(key_in[92]),
        .I1(key_derivation_en),
        .I2(enable_i[28]),
        .O(\KR[2].key_host[1][28]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair262" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][29]_i_1 
       (.I0(key_in[93]),
        .I1(key_derivation_en),
        .I2(enable_i[29]),
        .O(\KR[2].key_host[1][29]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][2]_i_1 
       (.I0(key_in[66]),
        .I1(key_derivation_en),
        .I2(enable_i[2]),
        .O(\KR[2].key_host[1][2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair264" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][30]_i_1 
       (.I0(key_in[94]),
        .I1(key_derivation_en),
        .I2(enable_i[30]),
        .O(\KR[2].key_host[1][30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair266" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][31]_i_2 
       (.I0(key_in[95]),
        .I1(key_derivation_en),
        .I2(enable_i[31]),
        .O(\KR[2].key_host[1][31]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][3]_i_1 
       (.I0(key_in[67]),
        .I1(key_derivation_en),
        .I2(enable_i[3]),
        .O(\KR[2].key_host[1][3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][4]_i_1 
       (.I0(key_in[68]),
        .I1(key_derivation_en),
        .I2(enable_i[4]),
        .O(\KR[2].key_host[1][4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][5]_i_1 
       (.I0(key_in[69]),
        .I1(key_derivation_en),
        .I2(enable_i[5]),
        .O(\KR[2].key_host[1][5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][6]_i_1 
       (.I0(key_in[70]),
        .I1(key_derivation_en),
        .I2(enable_i[6]),
        .O(\KR[2].key_host[1][6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][7]_i_1 
       (.I0(key_in[71]),
        .I1(key_derivation_en),
        .I2(enable_i[7]),
        .O(\KR[2].key_host[1][7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][8]_i_1 
       (.I0(key_in[72]),
        .I1(key_derivation_en),
        .I2(enable_i[8]),
        .O(\KR[2].key_host[1][8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[2].key_host[1][9]_i_1 
       (.I0(key_in[73]),
        .I1(key_derivation_en),
        .I2(enable_i[9]),
        .O(\KR[2].key_host[1][9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][0] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][0]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][10] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][10]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][11] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][11]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][12] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][12]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][13] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][13]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][14] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][14]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][15] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][15]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][16] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][16]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][17] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][17]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][18] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][18]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][19] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][19]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][1] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][1]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][20] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][20]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][21] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][21]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][22] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][22]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][23] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][23]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][24] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][24]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][25] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][25]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][26] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][26]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][27] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][27]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][28] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][28]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][29] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][29]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][2] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][2]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][30] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][30]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][31] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][31]_i_2_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][3] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][3]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][4] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][4]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][5] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][5]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][6] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][6]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][7] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][7]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][8] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][8]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_host_reg[1][9] 
       (.C(clk_i),
        .CE(\KR[2].key_host_reg[1][0]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_host[1][9]_i_1_n_0 ),
        .Q(\KR[2].key_host_reg[1][31]_0 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][0] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [0]),
        .Q(key_in[64]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][10] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [10]),
        .Q(key_in[74]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][11] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [11]),
        .Q(key_in[75]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][12] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [12]),
        .Q(key_in[76]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][13] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [13]),
        .Q(key_in[77]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][14] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [14]),
        .Q(key_in[78]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][15] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [15]),
        .Q(key_in[79]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][16] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [16]),
        .Q(key_in[80]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][17] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [17]),
        .Q(key_in[81]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][18] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [18]),
        .Q(key_in[82]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][19] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [19]),
        .Q(key_in[83]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][1] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [1]),
        .Q(key_in[65]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][20] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [20]),
        .Q(key_in[84]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][21] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [21]),
        .Q(key_in[85]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][22] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [22]),
        .Q(key_in[86]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][23] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [23]),
        .Q(key_in[87]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][24] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [24]),
        .Q(key_in[88]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][25] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [25]),
        .Q(key_in[89]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][26] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [26]),
        .Q(key_in[90]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][27] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [27]),
        .Q(key_in[91]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][28] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [28]),
        .Q(key_in[92]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][29] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [29]),
        .Q(key_in[93]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][2] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [2]),
        .Q(key_in[66]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][30] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [30]),
        .Q(key_in[94]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][31] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [31]),
        .Q(key_in[95]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][3] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [3]),
        .Q(key_in[67]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][4] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [4]),
        .Q(key_in[68]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][5] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [5]),
        .Q(key_in[69]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][6] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [6]),
        .Q(key_in[70]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][7] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [7]),
        .Q(key_in[71]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][8] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [8]),
        .Q(key_in[72]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[2].key_reg[1][9] 
       (.C(clk_i),
        .CE(\KR[2].key_reg[1][31]_0 ),
        .CLR(rst_i),
        .D(\KR[2].key_reg[1][31]_1 [9]),
        .Q(key_in[73]));
  (* SOFT_HLUTNM = "soft_lutpair235" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][0]_i_1 
       (.I0(key_in[96]),
        .I1(key_derivation_en),
        .I2(enable_i[0]),
        .O(\KR[3].key_host[0][0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][10]_i_1 
       (.I0(key_in[106]),
        .I1(key_derivation_en),
        .I2(enable_i[10]),
        .O(\KR[3].key_host[0][10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][11]_i_1 
       (.I0(key_in[107]),
        .I1(key_derivation_en),
        .I2(enable_i[11]),
        .O(\KR[3].key_host[0][11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][12]_i_1 
       (.I0(key_in[108]),
        .I1(key_derivation_en),
        .I2(enable_i[12]),
        .O(\KR[3].key_host[0][12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][13]_i_1 
       (.I0(key_in[109]),
        .I1(key_derivation_en),
        .I2(enable_i[13]),
        .O(\KR[3].key_host[0][13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][14]_i_1 
       (.I0(key_in[110]),
        .I1(key_derivation_en),
        .I2(enable_i[14]),
        .O(\KR[3].key_host[0][14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][15]_i_1 
       (.I0(key_in[111]),
        .I1(key_derivation_en),
        .I2(enable_i[15]),
        .O(\KR[3].key_host[0][15]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair237" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][16]_i_1 
       (.I0(key_in[112]),
        .I1(key_derivation_en),
        .I2(enable_i[16]),
        .O(\KR[3].key_host[0][16]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][17]_i_1 
       (.I0(key_in[113]),
        .I1(key_derivation_en),
        .I2(enable_i[17]),
        .O(\KR[3].key_host[0][17]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][18]_i_1 
       (.I0(key_in[114]),
        .I1(key_derivation_en),
        .I2(enable_i[18]),
        .O(\KR[3].key_host[0][18]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair243" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][19]_i_1 
       (.I0(key_in[115]),
        .I1(key_derivation_en),
        .I2(enable_i[19]),
        .O(\KR[3].key_host[0][19]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][1]_i_1 
       (.I0(key_in[97]),
        .I1(key_derivation_en),
        .I2(enable_i[1]),
        .O(\KR[3].key_host[0][1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair245" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][20]_i_1 
       (.I0(key_in[116]),
        .I1(key_derivation_en),
        .I2(enable_i[20]),
        .O(\KR[3].key_host[0][20]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair247" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][21]_i_1 
       (.I0(key_in[117]),
        .I1(key_derivation_en),
        .I2(enable_i[21]),
        .O(\KR[3].key_host[0][21]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair267" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][22]_i_1 
       (.I0(key_in[118]),
        .I1(key_derivation_en),
        .I2(enable_i[22]),
        .O(\KR[3].key_host[0][22]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair249" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][23]_i_1 
       (.I0(key_in[119]),
        .I1(key_derivation_en),
        .I2(enable_i[23]),
        .O(\KR[3].key_host[0][23]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair251" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][24]_i_1 
       (.I0(key_in[120]),
        .I1(key_derivation_en),
        .I2(enable_i[24]),
        .O(\KR[3].key_host[0][24]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair253" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][25]_i_1 
       (.I0(key_in[121]),
        .I1(key_derivation_en),
        .I2(enable_i[25]),
        .O(\KR[3].key_host[0][25]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair255" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][26]_i_1 
       (.I0(key_in[122]),
        .I1(key_derivation_en),
        .I2(enable_i[26]),
        .O(\KR[3].key_host[0][26]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair257" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][27]_i_1 
       (.I0(key_in[123]),
        .I1(key_derivation_en),
        .I2(enable_i[27]),
        .O(\KR[3].key_host[0][27]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair259" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][28]_i_1 
       (.I0(key_in[124]),
        .I1(key_derivation_en),
        .I2(enable_i[28]),
        .O(\KR[3].key_host[0][28]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair261" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][29]_i_1 
       (.I0(key_in[125]),
        .I1(key_derivation_en),
        .I2(enable_i[29]),
        .O(\KR[3].key_host[0][29]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][2]_i_1 
       (.I0(key_in[98]),
        .I1(key_derivation_en),
        .I2(enable_i[2]),
        .O(\KR[3].key_host[0][2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair263" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][30]_i_1 
       (.I0(key_in[126]),
        .I1(key_derivation_en),
        .I2(enable_i[30]),
        .O(\KR[3].key_host[0][30]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair265" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][31]_i_2 
       (.I0(key_in[127]),
        .I1(key_derivation_en),
        .I2(enable_i[31]),
        .O(\KR[3].key_host[0][31]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][3]_i_1 
       (.I0(key_in[99]),
        .I1(key_derivation_en),
        .I2(enable_i[3]),
        .O(\KR[3].key_host[0][3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][4]_i_1 
       (.I0(key_in[100]),
        .I1(key_derivation_en),
        .I2(enable_i[4]),
        .O(\KR[3].key_host[0][4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][5]_i_1 
       (.I0(key_in[101]),
        .I1(key_derivation_en),
        .I2(enable_i[5]),
        .O(\KR[3].key_host[0][5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][6]_i_1 
       (.I0(key_in[102]),
        .I1(key_derivation_en),
        .I2(enable_i[6]),
        .O(\KR[3].key_host[0][6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][7]_i_1 
       (.I0(key_in[103]),
        .I1(key_derivation_en),
        .I2(enable_i[7]),
        .O(\KR[3].key_host[0][7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][8]_i_1 
       (.I0(key_in[104]),
        .I1(key_derivation_en),
        .I2(enable_i[8]),
        .O(\KR[3].key_host[0][8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \KR[3].key_host[0][9]_i_1 
       (.I0(key_in[105]),
        .I1(key_derivation_en),
        .I2(enable_i[9]),
        .O(\KR[3].key_host[0][9]_i_1_n_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][0] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][0]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][10] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][10]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [10]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][11] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][11]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [11]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][12] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][12]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [12]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][13] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][13]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [13]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][14] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][14]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [14]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][15] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][15]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [15]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][16] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][16]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [16]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][17] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][17]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [17]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][18] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][18]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [18]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][19] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][19]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [19]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][1] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][1]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][20] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][20]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [20]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][21] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][21]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [21]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][22] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][22]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [22]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][23] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][23]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [23]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][24] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][24]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [24]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][25] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][25]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [25]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][26] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][26]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [26]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][27] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][27]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [27]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][28] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][28]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [28]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][29] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][29]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [29]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][2] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][2]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][30] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][30]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [30]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][31] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][31]_i_2_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [31]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][3] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][3]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][4] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][4]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][5] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][5]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][6] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][6]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][7] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][7]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [7]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][8] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][8]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [8]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_host_reg[0][9] 
       (.C(clk_i),
        .CE(\KR[3].key_host_reg[0][0]_0 ),
        .CLR(rst_i),
        .D(\KR[3].key_host[0][9]_i_1_n_0 ),
        .Q(\KR[3].key_host_reg[0]_3 [9]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][0] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_94),
        .Q(key_in[96]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][10] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_84),
        .Q(key_in[106]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][11] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_83),
        .Q(key_in[107]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][12] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_82),
        .Q(key_in[108]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][13] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_81),
        .Q(key_in[109]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][14] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_80),
        .Q(key_in[110]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][15] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_79),
        .Q(key_in[111]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][16] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_78),
        .Q(key_in[112]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][17] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_77),
        .Q(key_in[113]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][18] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_76),
        .Q(key_in[114]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][19] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_75),
        .Q(key_in[115]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][1] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_93),
        .Q(key_in[97]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][20] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_74),
        .Q(key_in[116]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][21] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_73),
        .Q(key_in[117]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][22] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_72),
        .Q(key_in[118]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][23] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_71),
        .Q(key_in[119]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][24] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_70),
        .Q(key_in[120]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][25] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_69),
        .Q(key_in[121]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][26] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_68),
        .Q(key_in[122]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][27] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_67),
        .Q(key_in[123]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][28] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_66),
        .Q(key_in[124]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][29] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_65),
        .Q(key_in[125]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][2] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_92),
        .Q(key_in[98]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][30] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_64),
        .Q(key_in[126]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][31] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_63),
        .Q(key_in[127]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][3] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_91),
        .Q(key_in[99]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][4] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_90),
        .Q(key_in[100]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][5] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_89),
        .Q(key_in[101]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][6] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_88),
        .Q(key_in[102]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][7] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_87),
        .Q(key_in[103]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][8] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_86),
        .Q(key_in[104]));
  FDCE #(
    .INIT(1'b0)) 
    \KR[3].key_reg[0][9] 
       (.C(clk_i),
        .CE(\KR[3].key_reg[0][31]_0 ),
        .CLR(rst_i),
        .D(SBOX_n_85),
        .Q(key_in[105]));
  switch_elements_sBox SBOX
       (.\CD[0].col[3][31]_i_14 (\CD[2].col_reg[1][31]_0 ),
        .\CD[0].col[3][31]_i_14_0 (\CD[1].col_reg[2][31]_0 ),
        .\CD[0].col[3][7]_i_9 (\CD[0].col[3][7]_i_9_0 ),
        .\CD[0].col[3][7]_i_9_0 (\CD[0].col[3][7]_i_9_1 ),
        .\CD[2].col_reg[1][0] (\CD[2].col_reg[1][0]_0 ),
        .\CD[2].col_reg[1][10] (SBOX_n_147),
        .\CD[2].col_reg[1][11] (SBOX_n_145),
        .\CD[2].col_reg[1][12] (SBOX_n_143),
        .\CD[2].col_reg[1][13] (\CD[2].col_reg[1][13]_0 ),
        .\CD[2].col_reg[1][14] (\CD[2].col_reg[1][14]_0 ),
        .\CD[2].col_reg[1][15] (SBOX_n_131),
        .\CD[2].col_reg[1][16] (\CD[2].col_reg[1][16]_0 ),
        .\CD[2].col_reg[1][17] (\CD[2].col_reg[1][17]_0 ),
        .\CD[2].col_reg[1][18] (SBOX_n_158),
        .\CD[2].col_reg[1][19] (SBOX_n_157),
        .\CD[2].col_reg[1][1] (\CD[2].col_reg[1][1]_0 ),
        .\CD[2].col_reg[1][20] (SBOX_n_156),
        .\CD[2].col_reg[1][21] (\CD[2].col_reg[1][21]_0 ),
        .\CD[2].col_reg[1][22] (\CD[2].col_reg[1][22]_0 ),
        .\CD[2].col_reg[1][23] (SBOX_n_153),
        .\CD[2].col_reg[1][24] (\CD[2].col_reg[1][24]_0 ),
        .\CD[2].col_reg[1][25] (\CD[2].col_reg[1][25]_0 ),
        .\CD[2].col_reg[1][26] (SBOX_n_148),
        .\CD[2].col_reg[1][27] (SBOX_n_146),
        .\CD[2].col_reg[1][28] (SBOX_n_144),
        .\CD[2].col_reg[1][29] (\CD[2].col_reg[1][29]_0 ),
        .\CD[2].col_reg[1][2] (SBOX_n_137),
        .\CD[2].col_reg[1][30] (\CD[2].col_reg[1][30]_0 ),
        .\CD[2].col_reg[1][31] (SBOX_n_132),
        .\CD[2].col_reg[1][3] (SBOX_n_141),
        .\CD[2].col_reg[1][4] (SBOX_n_142),
        .\CD[2].col_reg[1][5] (\CD[2].col_reg[1][5]_0 ),
        .\CD[2].col_reg[1][6] (\CD[2].col_reg[1][6]_0 ),
        .\CD[2].col_reg[1][7] (SBOX_n_130),
        .\CD[2].col_reg[1][8] (\CD[2].col_reg[1][8]_0 ),
        .\CD[2].col_reg[1][9] (\CD[2].col_reg[1][9]_0 ),
        .D({SBOX_n_6,SBOX_n_7,SBOX_n_8,SBOX_n_9,SBOX_n_10,SBOX_n_11,SBOX_n_12,SBOX_n_13,SBOX_n_14,SBOX_n_15,SBOX_n_16,SBOX_n_17,SBOX_n_18,SBOX_n_19,SBOX_n_20,SBOX_n_21,SBOX_n_22,SBOX_n_23,SBOX_n_24,SBOX_n_25,SBOX_n_26,SBOX_n_27,SBOX_n_28,SBOX_n_29,SBOX_n_30,SBOX_n_31,SBOX_n_32,SBOX_n_33,SBOX_n_34,SBOX_n_35,SBOX_n_36,SBOX_n_37}),
        .\KR[3].key_host_reg[0][31] ({SBOX_n_63,SBOX_n_64,SBOX_n_65,SBOX_n_66,SBOX_n_67,SBOX_n_68,SBOX_n_69,SBOX_n_70,SBOX_n_71,SBOX_n_72,SBOX_n_73,SBOX_n_74,SBOX_n_75,SBOX_n_76,SBOX_n_77,SBOX_n_78,SBOX_n_79,SBOX_n_80,SBOX_n_81,SBOX_n_82,SBOX_n_83,SBOX_n_84,SBOX_n_85,SBOX_n_86,SBOX_n_87,SBOX_n_88,SBOX_n_89,SBOX_n_90,SBOX_n_91,SBOX_n_92,SBOX_n_93,SBOX_n_94}),
        .\KR[3].key_reg[0][31] (\KR[3].key_host_reg[0]_3 ),
        .\KR[3].key_reg[0][31]_0 (key_in[127:96]),
        .Q(round_pp1),
        .\base_new_pp_reg[1] (p_86_in),
        .\base_new_pp_reg[1]_0 (p_86_in_5),
        .\base_new_pp_reg[1]_1 (p_86_in_11),
        .\base_new_pp_reg[2] (Q),
        .\base_new_pp_reg[3] (\base_new_pp_reg[3]_1 ),
        .\base_new_pp_reg[3]_0 (\base_new_pp_reg[3]_2 ),
        .\base_new_pp_reg[3]_1 (\base_new_pp_reg[3]_0 ),
        .\base_new_pp_reg[3]_2 (\base_new_pp_reg[3] ),
        .\base_new_pp_reg[4] (p_16_in),
        .\base_new_pp_reg[4]_0 (p_93_in),
        .\base_new_pp_reg[4]_1 (p_16_in_0),
        .\base_new_pp_reg[4]_2 (p_93_in_2),
        .\base_new_pp_reg[4]_3 (p_16_in_6),
        .\base_new_pp_reg[4]_4 (p_93_in_8),
        .\base_new_pp_reg[4]_5 (\base_new_pp_reg[4] ),
        .\base_new_pp_reg[4]_6 (\base_new_pp_reg[4]_2 ),
        .\base_new_pp_reg[4]_7 (\base_new_pp_reg[4]_3 ),
        .\base_new_pp_reg[4]_8 (\base_new_pp_reg[4]_1 ),
        .\base_new_pp_reg[4]_9 (\base_new_pp_reg[4]_0 ),
        .\base_new_pp_reg[6] (isomorphism_inv_return03_out),
        .\base_new_pp_reg[6]_0 (isomorphism_inv_return033_out),
        .\base_new_pp_reg[6]_1 (isomorphism_inv_return05_out),
        .\base_new_pp_reg[6]_2 (isomorphism_inv_return03_out_1),
        .\base_new_pp_reg[6]_3 (isomorphism_inv_return033_out_3),
        .\base_new_pp_reg[6]_4 (isomorphism_inv_return05_out_4),
        .\base_new_pp_reg[6]_5 (isomorphism_inv_return03_out_7),
        .\base_new_pp_reg[6]_6 (isomorphism_inv_return033_out_9),
        .\base_new_pp_reg[6]_7 (isomorphism_inv_return05_out_10),
        .clk_i(clk_i),
        .enable_i(enable_i),
        .enable_i_0_sp_1(enable_i_0_sn_1),
        .enc_dec_sbox(enc_dec_sbox),
        .g_func(g_func),
        .\info_o[28]_INST_0_i_7 (\info_o[28]_INST_0_i_7 ),
        .\info_o[28]_INST_0_i_7_0 (\info_o[28]_INST_0_i_7_0 ),
        .\info_o[31]_INST_0_i_11 (key_in[63:32]),
        .\info_o[31]_INST_0_i_11_0 (key_in[31:0]),
        .\info_o[31]_INST_0_i_9 (\CD[3].col_reg[0][31]_0 ),
        .isomorphism_return114_out(isomorphism_return114_out),
        .isomorphism_return114_out_13(isomorphism_return114_out_13),
        .isomorphism_return114_out_15(isomorphism_return114_out_15),
        .isomorphism_return114_out_17(isomorphism_return114_out_17),
        .isomorphism_return179_out(isomorphism_return179_out),
        .isomorphism_return179_out_12(isomorphism_return179_out_12),
        .isomorphism_return179_out_14(isomorphism_return179_out_14),
        .isomorphism_return179_out_16(isomorphism_return179_out_16),
        .key_en(key_en[0]),
        .key_sel_mux(key_sel_mux),
        .rc(\KEY_EXPANDER/rc ),
        .\round_pp1_reg[0] (\round_pp1_reg[0]_0 ),
        .\round_pp1_reg[0]_0 (\round_pp1_reg[0]_1 ),
        .\round_pp1_reg[0]_1 (\round_pp1_reg[0]_2 ),
        .\round_pp1_reg[3] (\round_pp1_reg[3]_0 ),
        .\round_pp1_reg[3]_0 (\round_pp1_reg[3]_1 ),
        .\round_pp1_reg[3]_1 (\round_pp1_reg[3]_2 ),
        .sbox_input(sbox_input),
        .sbox_out_enc(sbox_out_enc),
        .\sbox_pp2_reg[0] (key_out[0]),
        .\sbox_pp2_reg[10] (\KR[1].key_reg[2][10]_0 ),
        .\sbox_pp2_reg[11] (\KR[1].key_reg[2][11]_0 ),
        .\sbox_pp2_reg[12] (\KR[1].key_reg[2][12]_0 ),
        .\sbox_pp2_reg[13] (key_out[3]),
        .\sbox_pp2_reg[14] (key_out[4]),
        .\sbox_pp2_reg[15] (key_out[5]),
        .\sbox_pp2_reg[16] (key_out[6]),
        .\sbox_pp2_reg[17] (key_out[7]),
        .\sbox_pp2_reg[18] (key_out[8]),
        .\sbox_pp2_reg[19] (key_out[9]),
        .\sbox_pp2_reg[1] (\sbox_pp2[1]_i_3_n_0 ),
        .\sbox_pp2_reg[20] (key_out[10]),
        .\sbox_pp2_reg[21] (key_out[11]),
        .\sbox_pp2_reg[22] (key_out[12]),
        .\sbox_pp2_reg[23] (key_out[13]),
        .\sbox_pp2_reg[24] (key_out[14]),
        .\sbox_pp2_reg[25] (key_out[15]),
        .\sbox_pp2_reg[26] (key_out[16]),
        .\sbox_pp2_reg[27] (key_out[17]),
        .\sbox_pp2_reg[28] (key_out[18]),
        .\sbox_pp2_reg[29] (key_out[19]),
        .\sbox_pp2_reg[2] (\sbox_pp2[2]_i_3_n_0 ),
        .\sbox_pp2_reg[30] (key_out[20]),
        .\sbox_pp2_reg[31] (\sbox_pp2_reg[31]_0 ),
        .\sbox_pp2_reg[31]_0 (key_out[21]),
        .\sbox_pp2_reg[3] (\sbox_pp2[3]_i_2_n_0 ),
        .\sbox_pp2_reg[4] (\KR[1].key_reg[2][4]_0 ),
        .\sbox_pp2_reg[5] (\sbox_pp2[5]_i_3_n_0 ),
        .\sbox_pp2_reg[6] (\KR[1].key_reg[2][6]_0 ),
        .\sbox_pp2_reg[7] (key_out[1]),
        .\sbox_pp2_reg[8] (key_out[2]),
        .\sbox_pp2_reg[9] (\KR[1].key_reg[2][9]_0 ));
  switch_elements_data_swap SWAP_IN
       (.\IV_BKP_REGISTERS[3].bkp[3][31]_i_2 (\info_o[1] ),
        .bus_swap(bus_swap),
        .enable_i(enable_i));
  switch_elements_data_swap_0 SWAP_OUT
       (.\aes_cr_reg[2] (\aes_cr_reg[2]_0 ),
        .\aes_cr_reg[2]_0 (\aes_cr_reg[2] ),
        .col_out(col_out),
        .\info_o[1] (\info_o[1] ),
        .sbox_input(sbox_input));
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT5 #(
    .INIT(32'hFFFFBFFF)) 
    \aes_cr[10]_i_2 
       (.I0(enable_i[3]),
        .I1(enable_i[5]),
        .I2(enable_i[6]),
        .I3(enable_i[4]),
        .I4(enable_i[0]),
        .O(enable_i_3_sn_1));
  FDCE #(
    .INIT(1'b0)) 
    \col_en_cnt_unit_pp1_reg[0] 
       (.C(clk_i),
        .CE(\col_en_cnt_unit_pp1_reg[0]_0 ),
        .CLR(rst_i),
        .D(\col_en_cnt_unit_pp1_reg[3]_0 [0]),
        .Q(col_en_cnt_unit_pp1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \col_en_cnt_unit_pp1_reg[1] 
       (.C(clk_i),
        .CE(\col_en_cnt_unit_pp1_reg[0]_0 ),
        .CLR(rst_i),
        .D(\col_en_cnt_unit_pp1_reg[3]_0 [1]),
        .Q(col_en_cnt_unit_pp1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \col_en_cnt_unit_pp1_reg[2] 
       (.C(clk_i),
        .CE(\col_en_cnt_unit_pp1_reg[0]_0 ),
        .CLR(rst_i),
        .D(\col_en_cnt_unit_pp1_reg[3]_0 [2]),
        .Q(col_en_cnt_unit_pp1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \col_en_cnt_unit_pp1_reg[3] 
       (.C(clk_i),
        .CE(\col_en_cnt_unit_pp1_reg[0]_0 ),
        .CLR(rst_i),
        .D(\col_en_cnt_unit_pp1_reg[3]_0 [3]),
        .Q(col_en_cnt_unit_pp1[3]));
  FDCE #(
    .INIT(1'b0)) 
    \col_en_cnt_unit_pp2_reg[0] 
       (.C(clk_i),
        .CE(\col_en_cnt_unit_pp1_reg[0]_0 ),
        .CLR(rst_i),
        .D(col_en_cnt_unit_pp1[0]),
        .Q(\col_en_cnt_unit_pp2_reg[3]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \col_en_cnt_unit_pp2_reg[1] 
       (.C(clk_i),
        .CE(\col_en_cnt_unit_pp1_reg[0]_0 ),
        .CLR(rst_i),
        .D(col_en_cnt_unit_pp1[1]),
        .Q(\col_en_cnt_unit_pp2_reg[3]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \col_en_cnt_unit_pp2_reg[2] 
       (.C(clk_i),
        .CE(\col_en_cnt_unit_pp1_reg[0]_0 ),
        .CLR(rst_i),
        .D(col_en_cnt_unit_pp1[2]),
        .Q(\col_en_cnt_unit_pp2_reg[3]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \col_en_cnt_unit_pp2_reg[3] 
       (.C(clk_i),
        .CE(\col_en_cnt_unit_pp1_reg[0]_0 ),
        .CLR(rst_i),
        .D(col_en_cnt_unit_pp1[3]),
        .Q(\col_en_cnt_unit_pp2_reg[3]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \col_sel_pp1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\col_sel_pp1_reg[1]_0 [0]),
        .Q(col_sel_pp1[0]));
  FDPE #(
    .INIT(1'b1)) 
    \col_sel_pp1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\col_sel_pp1_reg[1]_0 [1]),
        .PRE(rst_i),
        .Q(col_sel_pp1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \col_sel_pp2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(col_sel_pp1[0]),
        .Q(\col_sel_pp2_reg[1]_0 [0]));
  FDPE #(
    .INIT(1'b1)) 
    \col_sel_pp2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(col_sel_pp1[1]),
        .PRE(rst_i),
        .Q(\col_sel_pp2_reg[1]_0 [1]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[0]_INST_0_i_2 
       (.I0(key_in[32]),
        .I1(key_in[0]),
        .I2(key_in[96]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[64]),
        .O(key_out[0]));
  LUT6 #(
    .INIT(64'hFF00F400F400F400)) 
    \info_o[0]_INST_0_i_4 
       (.I0(enable_i_0_sn_1),
        .I1(col_out),
        .I2(\info_o[0] ),
        .I3(\info_o[0]_0 ),
        .I4(\info_o[0]_1 ),
        .I5(\info_o[0]_2 ),
        .O(\aes_cr_reg[0] ));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[10]_INST_0_i_5 
       (.I0(key_in[42]),
        .I1(key_in[10]),
        .I2(key_in[106]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[74]),
        .O(\KR[1].key_reg[2][10]_0 ));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[11]_INST_0_i_5 
       (.I0(key_in[43]),
        .I1(key_in[11]),
        .I2(key_in[107]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[75]),
        .O(\KR[1].key_reg[2][11]_0 ));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[12]_INST_0_i_5 
       (.I0(key_in[44]),
        .I1(key_in[12]),
        .I2(key_in[108]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[76]),
        .O(\KR[1].key_reg[2][12]_0 ));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[13]_INST_0_i_2 
       (.I0(key_in[45]),
        .I1(key_in[13]),
        .I2(key_in[109]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[77]),
        .O(key_out[3]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[14]_INST_0_i_2 
       (.I0(key_in[46]),
        .I1(key_in[14]),
        .I2(key_in[110]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[78]),
        .O(key_out[4]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[15]_INST_0_i_2 
       (.I0(key_in[47]),
        .I1(key_in[15]),
        .I2(key_in[111]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[79]),
        .O(key_out[5]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[16]_INST_0_i_2 
       (.I0(key_in[48]),
        .I1(key_in[16]),
        .I2(key_in[112]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[80]),
        .O(key_out[6]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[17]_INST_0_i_2 
       (.I0(key_in[49]),
        .I1(key_in[17]),
        .I2(key_in[113]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[81]),
        .O(key_out[7]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[18]_INST_0_i_2 
       (.I0(key_in[50]),
        .I1(key_in[18]),
        .I2(key_in[114]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[82]),
        .O(key_out[8]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[19]_INST_0_i_2 
       (.I0(key_in[51]),
        .I1(key_in[19]),
        .I2(key_in[115]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[83]),
        .O(key_out[9]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[20]_INST_0_i_2 
       (.I0(key_in[52]),
        .I1(key_in[20]),
        .I2(key_in[116]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[84]),
        .O(key_out[10]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[21]_INST_0_i_2 
       (.I0(key_in[53]),
        .I1(key_in[21]),
        .I2(key_in[117]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[85]),
        .O(key_out[11]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[22]_INST_0_i_2 
       (.I0(key_in[54]),
        .I1(key_in[22]),
        .I2(key_in[118]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[86]),
        .O(key_out[12]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[23]_INST_0_i_2 
       (.I0(key_in[55]),
        .I1(key_in[23]),
        .I2(key_in[119]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[87]),
        .O(key_out[13]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[24]_INST_0_i_2 
       (.I0(key_in[56]),
        .I1(key_in[24]),
        .I2(key_in[120]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[88]),
        .O(key_out[14]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[25]_INST_0_i_2 
       (.I0(key_in[57]),
        .I1(key_in[25]),
        .I2(key_in[121]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[89]),
        .O(key_out[15]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[26]_INST_0_i_2 
       (.I0(key_in[58]),
        .I1(key_in[26]),
        .I2(key_in[122]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[90]),
        .O(key_out[16]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[27]_INST_0_i_2 
       (.I0(key_in[59]),
        .I1(key_in[27]),
        .I2(key_in[123]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[91]),
        .O(key_out[17]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[28]_INST_0_i_2 
       (.I0(key_in[60]),
        .I1(key_in[28]),
        .I2(key_in[124]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[92]),
        .O(key_out[18]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[29]_INST_0_i_2 
       (.I0(key_in[61]),
        .I1(key_in[29]),
        .I2(key_in[125]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[93]),
        .O(key_out[19]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[30]_INST_0_i_2 
       (.I0(key_in[62]),
        .I1(key_in[30]),
        .I2(key_in[126]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[94]),
        .O(key_out[20]));
  LUT6 #(
    .INIT(64'hFFFFFF00FFE2FFE2)) 
    \info_o[31]_INST_0_i_13 
       (.I0(key_out_sel_pp1),
        .I1(\sbox_pp2_reg[31]_0 ),
        .I2(key_out_sel_pp2),
        .I3(key_sel_rd),
        .I4(D[0]),
        .I5(bypass_key_en),
        .O(\info_o[31]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[31]_INST_0_i_4 
       (.I0(key_in[63]),
        .I1(key_in[31]),
        .I2(key_in[127]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[95]),
        .O(key_out[21]));
  LUT2 #(
    .INIT(4'hB)) 
    \info_o[31]_INST_0_i_41 
       (.I0(enable_i[2]),
        .I1(enable_i[1]),
        .O(enable_i_2_sn_1));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[4]_INST_0_i_5 
       (.I0(key_in[36]),
        .I1(key_in[4]),
        .I2(key_in[100]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[68]),
        .O(\KR[1].key_reg[2][4]_0 ));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[6]_INST_0_i_5 
       (.I0(key_in[38]),
        .I1(key_in[6]),
        .I2(key_in[102]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[70]),
        .O(\KR[1].key_reg[2][6]_0 ));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[7]_INST_0_i_2 
       (.I0(key_in[39]),
        .I1(key_in[7]),
        .I2(key_in[103]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[71]),
        .O(key_out[1]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[8]_INST_0_i_2 
       (.I0(key_in[40]),
        .I1(key_in[8]),
        .I2(key_in[104]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[72]),
        .O(key_out[2]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \info_o[9]_INST_0_i_5 
       (.I0(key_in[41]),
        .I1(key_in[9]),
        .I2(key_in[105]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[73]),
        .O(\KR[1].key_reg[2][9]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \key_en_pp1_reg[0] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\key_en_pp1_reg[3]_1 [0]),
        .Q(\key_en_pp1_reg[3]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \key_en_pp1_reg[1] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\key_en_pp1_reg[3]_1 [1]),
        .Q(\key_en_pp1_reg[3]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \key_en_pp1_reg[2] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\key_en_pp1_reg[3]_1 [2]),
        .Q(\key_en_pp1_reg[3]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \key_en_pp1_reg[3] 
       (.C(clk_i),
        .CE(E),
        .CLR(rst_i),
        .D(\key_en_pp1_reg[3]_1 [3]),
        .Q(\key_en_pp1_reg[3]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \key_out_sel_pp1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(D[0]),
        .Q(key_out_sel_pp1));
  FDCE #(
    .INIT(1'b0)) 
    \key_out_sel_pp1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(D[1]),
        .Q(\key_out_sel_pp1_reg[1]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    \key_out_sel_pp2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(key_out_sel_pp1),
        .Q(key_out_sel_pp2));
  FDCE #(
    .INIT(1'b0)) 
    \key_out_sel_pp2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\key_out_sel_pp1_reg[1]_0 ),
        .Q(\key_out_sel_pp2_reg[1]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    key_sel_pp1_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(key_sel),
        .Q(key_sel_pp1));
  FDPE #(
    .INIT(1'b1)) 
    last_round_pp1_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(last_round),
        .PRE(rst_i),
        .Q(last_round_pp1));
  FDCE #(
    .INIT(1'b0)) 
    last_round_pp2_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(last_round_pp1),
        .Q(last_round_pp2));
  FDPE #(
    .INIT(1'b1)) 
    rk_out_sel_pp1_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(rk_out_sel),
        .PRE(rst_i),
        .Q(rk_out_sel_pp1));
  FDPE #(
    .INIT(1'b1)) 
    rk_out_sel_pp2_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(rk_out_sel_pp1),
        .PRE(rst_i),
        .Q(rk_out_sel_pp2));
  FDCE #(
    .INIT(1'b0)) 
    \rk_sel_pp1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\rk_sel_pp1_reg[1]_0 [0]),
        .Q(rk_sel_pp1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rk_sel_pp1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\rk_sel_pp1_reg[1]_0 [1]),
        .Q(rk_sel_pp1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \rk_sel_pp2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(rk_sel_pp1[0]),
        .Q(rk_sel_pp2[0]));
  FDCE #(
    .INIT(1'b0)) 
    \rk_sel_pp2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(rk_sel_pp1[1]),
        .Q(rk_sel_pp2[1]));
  FDCE #(
    .INIT(1'b0)) 
    \round_pp1_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\round_pp1_reg[3]_3 [0]),
        .Q(round_pp1[0]));
  FDCE #(
    .INIT(1'b0)) 
    \round_pp1_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\round_pp1_reg[3]_3 [1]),
        .Q(round_pp1[1]));
  FDCE #(
    .INIT(1'b0)) 
    \round_pp1_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\round_pp1_reg[3]_3 [2]),
        .Q(round_pp1[2]));
  FDCE #(
    .INIT(1'b0)) 
    \round_pp1_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\round_pp1_reg[3]_3 [3]),
        .Q(round_pp1[3]));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \sbox_pp2[1]_i_3 
       (.I0(key_in[33]),
        .I1(key_in[1]),
        .I2(key_in[97]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[65]),
        .O(\sbox_pp2[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \sbox_pp2[2]_i_3 
       (.I0(key_in[34]),
        .I1(key_in[2]),
        .I2(key_in[98]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[66]),
        .O(\sbox_pp2[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \sbox_pp2[3]_i_2 
       (.I0(key_in[35]),
        .I1(key_in[3]),
        .I2(key_in[99]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[67]),
        .O(\sbox_pp2[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hCCFFAAF0CC00AAF0)) 
    \sbox_pp2[5]_i_3 
       (.I0(key_in[37]),
        .I1(key_in[5]),
        .I2(key_in[101]),
        .I3(\sbox_pp2_reg[5]_0 ),
        .I4(\info_o[31]_INST_0_i_13_n_0 ),
        .I5(key_in[69]),
        .O(\sbox_pp2[5]_i_3_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_37),
        .Q(sbox_pp2[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[10] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_27),
        .Q(sbox_pp2[10]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[11] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_26),
        .Q(sbox_pp2[11]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[12] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_25),
        .Q(sbox_pp2[12]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[13] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_24),
        .Q(sbox_pp2[13]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[14] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_23),
        .Q(sbox_pp2[14]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[15] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_22),
        .Q(sbox_pp2[15]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[16] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_21),
        .Q(sbox_pp2[16]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[17] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_20),
        .Q(sbox_pp2[17]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[18] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_19),
        .Q(sbox_pp2[18]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[19] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_18),
        .Q(sbox_pp2[19]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_36),
        .Q(sbox_pp2[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[20] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_17),
        .Q(sbox_pp2[20]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[21] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_16),
        .Q(sbox_pp2[21]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[22] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_15),
        .Q(sbox_pp2[22]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[23] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_14),
        .Q(sbox_pp2[23]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[24] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_13),
        .Q(sbox_pp2[24]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[25] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_12),
        .Q(sbox_pp2[25]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[26] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_11),
        .Q(sbox_pp2[26]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[27] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_10),
        .Q(sbox_pp2[27]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[28] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_9),
        .Q(sbox_pp2[28]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[29] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_8),
        .Q(sbox_pp2[29]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_35),
        .Q(sbox_pp2[2]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[30] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_7),
        .Q(sbox_pp2[30]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[31] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_6),
        .Q(sbox_pp2[31]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_34),
        .Q(sbox_pp2[3]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_33),
        .Q(sbox_pp2[4]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_32),
        .Q(sbox_pp2[5]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_31),
        .Q(sbox_pp2[6]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_30),
        .Q(sbox_pp2[7]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[8] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_29),
        .Q(sbox_pp2[8]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \sbox_pp2_reg[9] 
       (.C(clk_i),
        .CE(1'b1),
        .D(SBOX_n_28),
        .Q(sbox_pp2[9]),
        .R(1'b0));
endmodule

(* ORIG_REF_NAME = "host_interface" *) 
module switch_elements_host_interface
   (Q,
    ccf,
    first_block,
    info_o,
    \aes_cr_reg[7]_0 ,
    \aes_cr_reg[4]_0 ,
    \aes_cr_reg[0]_0 ,
    \aes_cr_reg[6]_0 ,
    \aes_cr_reg[7]_1 ,
    \aes_cr_reg[8]_0 ,
    \aes_cr_reg[9]_0 ,
    \aes_cr_reg[10]_0 ,
    \aes_cr_reg[4]_1 ,
    \aes_cr_reg[0]_1 ,
    \FSM_sequential_state_reg[0]_0 ,
    \aes_cr_reg[4]_2 ,
    \aes_cr_reg[5]_0 ,
    \FSM_sequential_state_reg[2]_0 ,
    \FSM_sequential_state_reg[2]_1 ,
    iv_en,
    enable_i_1_sp_1,
    key_en,
    \FSM_sequential_state_reg[0]_1 ,
    key_sel_rd,
    enable_i_2_sp_1,
    \enable_i[1]_0 ,
    \enable_i[2]_0 ,
    col_en_host,
    key_derivation_en,
    \FSM_sequential_state_reg[3] ,
    \aes_cr_reg[3]_0 ,
    \aes_cr_reg[0]_2 ,
    \FSM_sequential_state_reg[2]_2 ,
    \FSM_sequential_state_reg[2]_3 ,
    \aes_cr_reg[4]_3 ,
    \aes_cr_reg[6]_1 ,
    \aes_cr_reg[4]_4 ,
    enc_dec,
    \aes_cr_reg[6]_2 ,
    \FSM_sequential_state_reg[2]_4 ,
    \aes_cr_reg[4]_5 ,
    first_block_reg_0,
    \aes_cr_reg[4]_6 ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][0] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][0] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][0] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][0] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][1] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][1] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][1] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][1] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][2] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][2] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][2] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][2] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][3] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][3] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][3] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][3] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][4] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][4] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][4] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][4] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][5] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][5] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][5] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][5] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][6] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][6] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][6] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][6] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][7] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][7] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][7] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][7] ,
    \aes_cr_reg[5]_1 ,
    \aes_cr_reg[5]_2 ,
    \CD[2].col_reg[1][15] ,
    D,
    \aes_cr_reg[5]_3 ,
    \aes_cr_reg[5]_4 ,
    \aes_cr_reg[5]_5 ,
    \aes_cr_reg[5]_6 ,
    \aes_cr_reg[5]_7 ,
    \aes_cr_reg[5]_8 ,
    \aes_cr_reg[5]_9 ,
    \aes_cr_reg[5]_10 ,
    \aes_cr_reg[5]_11 ,
    \aes_cr_reg[5]_12 ,
    \aes_cr_reg[5]_13 ,
    \aes_cr_reg[5]_14 ,
    \aes_cr_reg[5]_15 ,
    \aes_cr_reg[5]_16 ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][16] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][16] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][16] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][16] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][17] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][17] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][17] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][17] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][18] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][18] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][18] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][18] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][19] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][19] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][19] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][19] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][20] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][20] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][20] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][20] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][21] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][21] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][21] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][21] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][22] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][22] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][22] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][22] ,
    \IV_BKP_REGISTERS[3].bkp_1_reg[3][23] ,
    \IV_BKP_REGISTERS[2].bkp_1_reg[2][23] ,
    \IV_BKP_REGISTERS[1].bkp_1_reg[1][23] ,
    \IV_BKP_REGISTERS[0].bkp_1_reg[0][23] ,
    \CD[1].col_reg[2][31] ,
    \CD[2].col_reg[1][31] ,
    \aes_cr_reg[5]_17 ,
    \aes_cr_reg[5]_18 ,
    \aes_cr_reg[5]_19 ,
    \aes_cr_reg[5]_20 ,
    \aes_cr_reg[5]_21 ,
    \aes_cr_reg[5]_22 ,
    \aes_cr_reg[5]_23 ,
    \aes_cr_reg[5]_24 ,
    \aes_cr_reg[5]_25 ,
    \aes_cr_reg[5]_26 ,
    \aes_cr_reg[5]_27 ,
    \aes_cr_reg[5]_28 ,
    \aes_cr_reg[5]_29 ,
    \aes_cr_reg[5]_30 ,
    \aes_cr_reg[5]_31 ,
    \aes_cr_reg[5]_32 ,
    E,
    \enable_i[4] ,
    \FSM_sequential_state_reg[2]_5 ,
    \enable_i[2]_1 ,
    first_block_reg_1,
    \col_en_cnt_unit_pp2_reg[3] ,
    rk_out_sel,
    \aes_cr_reg[5]_33 ,
    \col_en_cnt_unit_pp2_reg[3]_0 ,
    \col_en_cnt_unit_pp2_reg[2] ,
    \col_en_cnt_unit_pp2_reg[1] ,
    \col_en_cnt_unit_pp2_reg[0] ,
    \aes_cr_reg[5]_34 ,
    \aes_cr_reg[5]_35 ,
    clk_i,
    rst_i,
    ccf_reg_0,
    \info_o[3] ,
    info_o_1_sp_1,
    \info_o[3]_0 ,
    \info_o[12] ,
    \FSM_sequential_state_reg[0]_2 ,
    \cnt_reg[0]_0 ,
    enable_i,
    \FSM_sequential_state_reg[1]_0 ,
    \FSM_sequential_state_reg[1]_1 ,
    rk_out_sel_pp1_reg,
    \FSM_sequential_state_reg[1]_2 ,
    \FSM_sequential_state_reg[0]_3 ,
    \FSM_sequential_state_reg[0]_4 ,
    \aes_cr_reg[0]_3 ,
    \KR[1].key_host_reg[2][0] ,
    \info_o[0]_INST_0_i_4 ,
    info_o_2_sp_1,
    \info_o[31]_INST_0_i_15 ,
    \KR[0].key_host_reg[3][0] ,
    \IV_BKP_REGISTERS[3].iv_reg[3][0] ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][31] ,
    bus_swap,
    \IV_BKP_REGISTERS[2].bkp_reg[2][31] ,
    \IV_BKP_REGISTERS[1].bkp_reg[1][31] ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][31] ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 ,
    \IV_BKP_REGISTERS[0].bkp_reg[0][8] ,
    data_in,
    \IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 ,
    \IV_BKP_REGISTERS[3].bkp_reg[3][8] ,
    iv_mux_out16_out,
    \IV_BKP_REGISTERS[3].bkp_reg[3][0] ,
    bypass_rk,
    \CD[0].col[3][10]_i_12 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][0]_0 ,
    \IV_BKP_REGISTERS[3].iv_reg[3][0]_1 ,
    \IV_BKP_REGISTERS[2].bkp_reg[2][31]_2 );
  output [1:0]Q;
  output ccf;
  output first_block;
  output [2:0]info_o;
  output [6:0]\aes_cr_reg[7]_0 ;
  output \aes_cr_reg[4]_0 ;
  output \aes_cr_reg[0]_0 ;
  output \aes_cr_reg[6]_0 ;
  output \aes_cr_reg[7]_1 ;
  output \aes_cr_reg[8]_0 ;
  output \aes_cr_reg[9]_0 ;
  output \aes_cr_reg[10]_0 ;
  output \aes_cr_reg[4]_1 ;
  output \aes_cr_reg[0]_1 ;
  output \FSM_sequential_state_reg[0]_0 ;
  output [0:0]\aes_cr_reg[4]_2 ;
  output \aes_cr_reg[5]_0 ;
  output \FSM_sequential_state_reg[2]_0 ;
  output \FSM_sequential_state_reg[2]_1 ;
  output [2:0]iv_en;
  output enable_i_1_sp_1;
  output [3:0]key_en;
  output \FSM_sequential_state_reg[0]_1 ;
  output [0:0]key_sel_rd;
  output enable_i_2_sp_1;
  output \enable_i[1]_0 ;
  output \enable_i[2]_0 ;
  output [3:0]col_en_host;
  output key_derivation_en;
  output \FSM_sequential_state_reg[3] ;
  output \aes_cr_reg[3]_0 ;
  output \aes_cr_reg[0]_2 ;
  output \FSM_sequential_state_reg[2]_2 ;
  output \FSM_sequential_state_reg[2]_3 ;
  output \aes_cr_reg[4]_3 ;
  output \aes_cr_reg[6]_1 ;
  output \aes_cr_reg[4]_4 ;
  output enc_dec;
  output \aes_cr_reg[6]_2 ;
  output \FSM_sequential_state_reg[2]_4 ;
  output \aes_cr_reg[4]_5 ;
  output first_block_reg_0;
  output \aes_cr_reg[4]_6 ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][0] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][0] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][0] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][0] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][1] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][1] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][1] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][1] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][2] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][2] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][2] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][2] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][3] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][3] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][3] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][3] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][4] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][4] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][4] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][4] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][5] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][5] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][5] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][5] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][6] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][6] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][6] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][6] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][7] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][7] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][7] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][7] ;
  output \aes_cr_reg[5]_1 ;
  output \aes_cr_reg[5]_2 ;
  output [7:0]\CD[2].col_reg[1][15] ;
  output [7:0]D;
  output \aes_cr_reg[5]_3 ;
  output \aes_cr_reg[5]_4 ;
  output \aes_cr_reg[5]_5 ;
  output \aes_cr_reg[5]_6 ;
  output \aes_cr_reg[5]_7 ;
  output \aes_cr_reg[5]_8 ;
  output \aes_cr_reg[5]_9 ;
  output \aes_cr_reg[5]_10 ;
  output \aes_cr_reg[5]_11 ;
  output \aes_cr_reg[5]_12 ;
  output \aes_cr_reg[5]_13 ;
  output \aes_cr_reg[5]_14 ;
  output \aes_cr_reg[5]_15 ;
  output \aes_cr_reg[5]_16 ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][16] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][16] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][16] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][16] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][17] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][17] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][17] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][17] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][18] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][18] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][18] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][18] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][19] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][19] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][19] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][19] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][20] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][20] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][20] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][20] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][21] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][21] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][21] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][21] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][22] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][22] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][22] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][22] ;
  output \IV_BKP_REGISTERS[3].bkp_1_reg[3][23] ;
  output \IV_BKP_REGISTERS[2].bkp_1_reg[2][23] ;
  output \IV_BKP_REGISTERS[1].bkp_1_reg[1][23] ;
  output \IV_BKP_REGISTERS[0].bkp_1_reg[0][23] ;
  output [7:0]\CD[1].col_reg[2][31] ;
  output [7:0]\CD[2].col_reg[1][31] ;
  output \aes_cr_reg[5]_17 ;
  output \aes_cr_reg[5]_18 ;
  output \aes_cr_reg[5]_19 ;
  output \aes_cr_reg[5]_20 ;
  output \aes_cr_reg[5]_21 ;
  output \aes_cr_reg[5]_22 ;
  output \aes_cr_reg[5]_23 ;
  output \aes_cr_reg[5]_24 ;
  output \aes_cr_reg[5]_25 ;
  output \aes_cr_reg[5]_26 ;
  output \aes_cr_reg[5]_27 ;
  output \aes_cr_reg[5]_28 ;
  output \aes_cr_reg[5]_29 ;
  output \aes_cr_reg[5]_30 ;
  output \aes_cr_reg[5]_31 ;
  output \aes_cr_reg[5]_32 ;
  output [0:0]E;
  output [0:0]\enable_i[4] ;
  output [0:0]\FSM_sequential_state_reg[2]_5 ;
  output [0:0]\enable_i[2]_1 ;
  output first_block_reg_1;
  output \col_en_cnt_unit_pp2_reg[3] ;
  output rk_out_sel;
  output [0:0]\aes_cr_reg[5]_33 ;
  output [0:0]\col_en_cnt_unit_pp2_reg[3]_0 ;
  output [0:0]\col_en_cnt_unit_pp2_reg[2] ;
  output [0:0]\col_en_cnt_unit_pp2_reg[1] ;
  output [0:0]\col_en_cnt_unit_pp2_reg[0] ;
  output \aes_cr_reg[5]_34 ;
  output \aes_cr_reg[5]_35 ;
  input clk_i;
  input rst_i;
  input ccf_reg_0;
  input [2:0]\info_o[3] ;
  input info_o_1_sp_1;
  input \info_o[3]_0 ;
  input [5:0]\info_o[12] ;
  input \FSM_sequential_state_reg[0]_2 ;
  input \cnt_reg[0]_0 ;
  input [11:0]enable_i;
  input \FSM_sequential_state_reg[1]_0 ;
  input \FSM_sequential_state_reg[1]_1 ;
  input [3:0]rk_out_sel_pp1_reg;
  input \FSM_sequential_state_reg[1]_2 ;
  input [0:0]\FSM_sequential_state_reg[0]_3 ;
  input \FSM_sequential_state_reg[0]_4 ;
  input \aes_cr_reg[0]_3 ;
  input \KR[1].key_host_reg[2][0] ;
  input \info_o[0]_INST_0_i_4 ;
  input info_o_2_sp_1;
  input \info_o[31]_INST_0_i_15 ;
  input \KR[0].key_host_reg[3][0] ;
  input \IV_BKP_REGISTERS[3].iv_reg[3][0] ;
  input [31:0]\IV_BKP_REGISTERS[3].bkp_reg[3][31] ;
  input [31:0]bus_swap;
  input [31:0]\IV_BKP_REGISTERS[2].bkp_reg[2][31] ;
  input [31:0]\IV_BKP_REGISTERS[1].bkp_reg[1][31] ;
  input [31:0]\IV_BKP_REGISTERS[0].bkp_reg[0][31] ;
  input [31:0]\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 ;
  input \IV_BKP_REGISTERS[0].bkp_reg[0][8] ;
  input [15:0]data_in;
  input [15:0]\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 ;
  input \IV_BKP_REGISTERS[3].bkp_reg[3][8] ;
  input iv_mux_out16_out;
  input [3:0]\IV_BKP_REGISTERS[3].bkp_reg[3][0] ;
  input bypass_rk;
  input [0:0]\CD[0].col[3][10]_i_12 ;
  input \IV_BKP_REGISTERS[3].iv_reg[3][0]_0 ;
  input \IV_BKP_REGISTERS[3].iv_reg[3][0]_1 ;
  input \IV_BKP_REGISTERS[2].bkp_reg[2][31]_2 ;

  wire [0:0]\CD[0].col[3][10]_i_12 ;
  wire [7:0]\CD[1].col_reg[2][31] ;
  wire [7:0]\CD[2].col_reg[1][15] ;
  wire [7:0]\CD[2].col_reg[1][31] ;
  wire [7:0]D;
  wire [0:0]E;
  wire \FSM_sequential_state[0]_i_1_n_0 ;
  wire \FSM_sequential_state[0]_i_2__0_n_0 ;
  wire \FSM_sequential_state[0]_i_4__0_n_0 ;
  wire \FSM_sequential_state[1]_i_1_n_0 ;
  wire \FSM_sequential_state[1]_i_2__0_n_0 ;
  wire \FSM_sequential_state[1]_i_2_n_0 ;
  wire \FSM_sequential_state[1]_i_3_n_0 ;
  wire \FSM_sequential_state[1]_i_4_n_0 ;
  wire \FSM_sequential_state[1]_i_5__0_n_0 ;
  wire \FSM_sequential_state[1]_i_5_n_0 ;
  wire \FSM_sequential_state[1]_i_6__0_n_0 ;
  wire \FSM_sequential_state[1]_i_6_n_0 ;
  wire \FSM_sequential_state[2]_i_1_n_0 ;
  wire \FSM_sequential_state[2]_i_2_n_0 ;
  wire \FSM_sequential_state[2]_i_4_n_0 ;
  wire \FSM_sequential_state_reg[0]_0 ;
  wire \FSM_sequential_state_reg[0]_1 ;
  wire \FSM_sequential_state_reg[0]_2 ;
  wire [0:0]\FSM_sequential_state_reg[0]_3 ;
  wire \FSM_sequential_state_reg[0]_4 ;
  wire \FSM_sequential_state_reg[1]_0 ;
  wire \FSM_sequential_state_reg[1]_1 ;
  wire \FSM_sequential_state_reg[1]_2 ;
  wire \FSM_sequential_state_reg[2]_0 ;
  wire \FSM_sequential_state_reg[2]_1 ;
  wire \FSM_sequential_state_reg[2]_2 ;
  wire \FSM_sequential_state_reg[2]_3 ;
  wire \FSM_sequential_state_reg[2]_4 ;
  wire [0:0]\FSM_sequential_state_reg[2]_5 ;
  wire \FSM_sequential_state_reg[3] ;
  wire \IV_BKP_REGISTERS[0].bkp[0][10]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][11]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][12]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][13]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][14]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][15]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][8]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp[0][9]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][0] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][16] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][17] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][18] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][19] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][1] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][20] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][21] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][22] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][23] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][2] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][3] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][4] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][5] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][6] ;
  wire \IV_BKP_REGISTERS[0].bkp_1_reg[0][7] ;
  wire [31:0]\IV_BKP_REGISTERS[0].bkp_reg[0][31] ;
  wire \IV_BKP_REGISTERS[0].bkp_reg[0][8] ;
  wire \IV_BKP_REGISTERS[1].bkp[1][24]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][25]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][26]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][27]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][28]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][29]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][30]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp[1][31]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][0] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][16] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][17] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][18] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][19] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][1] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][20] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][21] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][22] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][23] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][2] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][3] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][4] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][5] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][6] ;
  wire \IV_BKP_REGISTERS[1].bkp_1_reg[1][7] ;
  wire [31:0]\IV_BKP_REGISTERS[1].bkp_reg[1][31] ;
  wire \IV_BKP_REGISTERS[2].bkp[2][24]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][24]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][25]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][25]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][26]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][26]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][27]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][27]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][28]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][28]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][29]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][29]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][30]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][30]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][31]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp[2][31]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][0] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][16] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][17] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][18] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][19] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][1] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][20] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][21] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][22] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][23] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][2] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][3] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][4] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][5] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][6] ;
  wire \IV_BKP_REGISTERS[2].bkp_1_reg[2][7] ;
  wire [31:0]\IV_BKP_REGISTERS[2].bkp_reg[2][31] ;
  wire [31:0]\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 ;
  wire [15:0]\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 ;
  wire \IV_BKP_REGISTERS[2].bkp_reg[2][31]_2 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][10]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][10]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][11]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][11]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][12]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][12]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][13]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][13]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][14]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][14]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][15]_i_5_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][15]_i_6_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][8]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][8]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][9]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp[3][9]_i_4_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_1[3][31]_i_2_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_1[3][31]_i_3_n_0 ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][0] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][16] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][17] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][18] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][19] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][1] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][20] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][21] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][22] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][23] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][2] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][3] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][4] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][5] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][6] ;
  wire \IV_BKP_REGISTERS[3].bkp_1_reg[3][7] ;
  wire [3:0]\IV_BKP_REGISTERS[3].bkp_reg[3][0] ;
  wire [31:0]\IV_BKP_REGISTERS[3].bkp_reg[3][31] ;
  wire \IV_BKP_REGISTERS[3].bkp_reg[3][8] ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][0] ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][0]_0 ;
  wire \IV_BKP_REGISTERS[3].iv_reg[3][0]_1 ;
  wire \KR[0].key_host_reg[3][0] ;
  wire \KR[1].key_host_reg[2][0] ;
  wire [1:0]Q;
  wire access_permission;
  wire aes_cr1;
  wire \aes_cr[0]_i_1_n_0 ;
  wire \aes_cr[0]_i_2_n_0 ;
  wire \aes_cr_reg[0]_0 ;
  wire \aes_cr_reg[0]_1 ;
  wire \aes_cr_reg[0]_2 ;
  wire \aes_cr_reg[0]_3 ;
  wire \aes_cr_reg[10]_0 ;
  wire \aes_cr_reg[3]_0 ;
  wire \aes_cr_reg[4]_0 ;
  wire \aes_cr_reg[4]_1 ;
  wire [0:0]\aes_cr_reg[4]_2 ;
  wire \aes_cr_reg[4]_3 ;
  wire \aes_cr_reg[4]_4 ;
  wire \aes_cr_reg[4]_5 ;
  wire \aes_cr_reg[4]_6 ;
  wire \aes_cr_reg[5]_0 ;
  wire \aes_cr_reg[5]_1 ;
  wire \aes_cr_reg[5]_10 ;
  wire \aes_cr_reg[5]_11 ;
  wire \aes_cr_reg[5]_12 ;
  wire \aes_cr_reg[5]_13 ;
  wire \aes_cr_reg[5]_14 ;
  wire \aes_cr_reg[5]_15 ;
  wire \aes_cr_reg[5]_16 ;
  wire \aes_cr_reg[5]_17 ;
  wire \aes_cr_reg[5]_18 ;
  wire \aes_cr_reg[5]_19 ;
  wire \aes_cr_reg[5]_2 ;
  wire \aes_cr_reg[5]_20 ;
  wire \aes_cr_reg[5]_21 ;
  wire \aes_cr_reg[5]_22 ;
  wire \aes_cr_reg[5]_23 ;
  wire \aes_cr_reg[5]_24 ;
  wire \aes_cr_reg[5]_25 ;
  wire \aes_cr_reg[5]_26 ;
  wire \aes_cr_reg[5]_27 ;
  wire \aes_cr_reg[5]_28 ;
  wire \aes_cr_reg[5]_29 ;
  wire \aes_cr_reg[5]_3 ;
  wire \aes_cr_reg[5]_30 ;
  wire \aes_cr_reg[5]_31 ;
  wire \aes_cr_reg[5]_32 ;
  wire [0:0]\aes_cr_reg[5]_33 ;
  wire \aes_cr_reg[5]_34 ;
  wire \aes_cr_reg[5]_35 ;
  wire \aes_cr_reg[5]_4 ;
  wire \aes_cr_reg[5]_5 ;
  wire \aes_cr_reg[5]_6 ;
  wire \aes_cr_reg[5]_7 ;
  wire \aes_cr_reg[5]_8 ;
  wire \aes_cr_reg[5]_9 ;
  wire \aes_cr_reg[6]_0 ;
  wire \aes_cr_reg[6]_1 ;
  wire \aes_cr_reg[6]_2 ;
  wire [6:0]\aes_cr_reg[7]_0 ;
  wire \aes_cr_reg[7]_1 ;
  wire \aes_cr_reg[8]_0 ;
  wire \aes_cr_reg[9]_0 ;
  wire [31:0]bus_swap;
  wire bypass_rk;
  wire ccf;
  wire ccf_reg_0;
  wire clk_i;
  wire \cnt[0]_i_1_n_0 ;
  wire \cnt[1]_i_1_n_0 ;
  wire \cnt[1]_i_2_n_0 ;
  wire \cnt[1]_i_3_n_0 ;
  wire \cnt[1]_i_4_n_0 ;
  wire \cnt_reg[0]_0 ;
  wire [0:0]\col_en_cnt_unit_pp2_reg[0] ;
  wire [0:0]\col_en_cnt_unit_pp2_reg[1] ;
  wire [0:0]\col_en_cnt_unit_pp2_reg[2] ;
  wire \col_en_cnt_unit_pp2_reg[3] ;
  wire [0:0]\col_en_cnt_unit_pp2_reg[3]_0 ;
  wire [3:0]col_en_host;
  wire [15:0]data_in;
  wire dma_in_en;
  wire dma_out_en;
  wire dma_req;
  wire [11:0]enable_i;
  wire \enable_i[1]_0 ;
  wire \enable_i[2]_0 ;
  wire [0:0]\enable_i[2]_1 ;
  wire [0:0]\enable_i[4] ;
  wire enable_i_1_sn_1;
  wire enable_i_2_sn_1;
  wire enc_dec;
  wire err_ie;
  wire first_block;
  wire first_block_i_1_n_0;
  wire first_block_reg_0;
  wire first_block_reg_1;
  wire [2:0]info_o;
  wire \info_o[0]_INST_0_i_4 ;
  wire [5:0]\info_o[12] ;
  wire \info_o[2]_INST_0_i_1_n_0 ;
  wire \info_o[2]_INST_0_i_2_n_0 ;
  wire \info_o[31]_INST_0_i_15 ;
  wire \info_o[31]_INST_0_i_44_n_0 ;
  wire [2:0]\info_o[3] ;
  wire \info_o[3]_0 ;
  wire \info_o[3]_INST_0_i_1_n_0 ;
  wire \info_o[3]_INST_0_i_4_n_0 ;
  wire info_o_1_sn_1;
  wire info_o_2_sn_1;
  wire [2:0]iv_en;
  wire iv_mux_out16_out;
  wire [3:3]iv_sel_rd;
  wire key_derivation_en;
  wire [3:0]key_en;
  wire [0:0]key_sel_rd;
  wire [3:3]p_1_in__0;
  wire rk_out_sel;
  wire [3:0]rk_out_sel_pp1_reg;
  wire rst_i;
  wire [2:0]state;
  wire wr_err;
  wire wr_err_en;
  wire wr_err_i_1_n_0;

  assign enable_i_1_sp_1 = enable_i_1_sn_1;
  assign enable_i_2_sp_1 = enable_i_2_sn_1;
  assign info_o_1_sn_1 = info_o_1_sp_1;
  assign info_o_2_sn_1 = info_o_2_sp_1;
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEEEFE)) 
    \CD[0].col[3][28]_i_18 
       (.I0(iv_sel_rd),
        .I1(col_en_host[3]),
        .I2(\IV_BKP_REGISTERS[3].bkp_reg[3][0] [3]),
        .I3(bypass_rk),
        .I4(\CD[0].col[3][10]_i_12 ),
        .I5(first_block_reg_0),
        .O(\col_en_cnt_unit_pp2_reg[3] ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \CD[0].col[3][28]_i_21 
       (.I0(enable_i[3]),
        .I1(enable_i[2]),
        .I2(access_permission),
        .I3(enable_i[1]),
        .I4(enable_i[0]),
        .O(iv_sel_rd));
  LUT3 #(
    .INIT(8'hB0)) 
    \CD[0].col[3][31]_i_21 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(first_block),
        .O(\aes_cr_reg[5]_35 ));
  (* SOFT_HLUTNM = "soft_lutpair294" *) 
  LUT4 #(
    .INIT(16'h5D00)) 
    \CD[0].col[3][31]_i_22 
       (.I0(first_block),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(iv_mux_out16_out),
        .O(first_block_reg_1));
  (* SOFT_HLUTNM = "soft_lutpair287" *) 
  LUT5 #(
    .INIT(32'hD5D500D5)) 
    \CD[0].col[3][31]_i_24 
       (.I0(\aes_cr_reg[7]_0 [3]),
        .I1(rk_out_sel_pp1_reg[1]),
        .I2(rk_out_sel_pp1_reg[2]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(\aes_cr_reg[7]_0 [4]),
        .O(\aes_cr_reg[4]_5 ));
  (* SOFT_HLUTNM = "soft_lutpair294" *) 
  LUT3 #(
    .INIT(8'hA2)) 
    \CD[0].col[3][31]_i_36 
       (.I0(first_block),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(\aes_cr_reg[7]_0 [4]),
        .O(first_block_reg_0));
  LUT6 #(
    .INIT(64'h2202020266666666)) 
    \CD[0].col[3][31]_i_9 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(\aes_cr_reg[7]_0 [3]),
        .I3(rk_out_sel_pp1_reg[1]),
        .I4(rk_out_sel_pp1_reg[2]),
        .I5(\IV_BKP_REGISTERS[3].iv_reg[3][0] ),
        .O(\aes_cr_reg[5]_34 ));
  LUT6 #(
    .INIT(64'h44FF444F00000000)) 
    \FSM_sequential_state[0]_i_1 
       (.I0(\FSM_sequential_state[0]_i_2__0_n_0 ),
        .I1(\FSM_sequential_state_reg[0]_0 ),
        .I2(\aes_cr_reg[4]_1 ),
        .I3(\FSM_sequential_state[0]_i_4__0_n_0 ),
        .I4(state[0]),
        .I5(\aes_cr_reg[0]_1 ),
        .O(\FSM_sequential_state[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair285" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \FSM_sequential_state[0]_i_2__0 
       (.I0(Q[0]),
        .I1(Q[1]),
        .O(\FSM_sequential_state[0]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    \FSM_sequential_state[0]_i_3 
       (.I0(state[0]),
        .I1(state[2]),
        .I2(state[1]),
        .I3(enable_i[2]),
        .I4(enable_i[1]),
        .I5(\aes_cr_reg[0]_3 ),
        .O(\FSM_sequential_state_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0000EFEF0000FF00)) 
    \FSM_sequential_state[0]_i_4 
       (.I0(state[2]),
        .I1(state[1]),
        .I2(state[0]),
        .I3(\FSM_sequential_state_reg[0]_3 ),
        .I4(\FSM_sequential_state_reg[0]_4 ),
        .I5(rk_out_sel_pp1_reg[0]),
        .O(\FSM_sequential_state_reg[2]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair292" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_state[0]_i_4__0 
       (.I0(state[1]),
        .I1(state[2]),
        .O(\FSM_sequential_state[0]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT5 #(
    .INIT(32'h20002020)) 
    \FSM_sequential_state[0]_i_8 
       (.I0(rk_out_sel_pp1_reg[3]),
        .I1(rk_out_sel_pp1_reg[2]),
        .I2(\aes_cr_reg[7]_0 [3]),
        .I3(\aes_cr_reg[7]_0 [4]),
        .I4(\aes_cr_reg[7]_0 [5]),
        .O(\FSM_sequential_state_reg[3] ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFAABAAA)) 
    \FSM_sequential_state[1]_i_1 
       (.I0(\FSM_sequential_state[1]_i_2__0_n_0 ),
        .I1(state[2]),
        .I2(\aes_cr_reg[4]_1 ),
        .I3(\aes_cr_reg[0]_1 ),
        .I4(state[0]),
        .I5(state[1]),
        .O(\FSM_sequential_state[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAAAABFAAAAAA)) 
    \FSM_sequential_state[1]_i_1__0 
       (.I0(\FSM_sequential_state[1]_i_2_n_0 ),
        .I1(\aes_cr_reg[5]_0 ),
        .I2(\aes_cr_reg[7]_0 [3]),
        .I3(\FSM_sequential_state_reg[1]_0 ),
        .I4(\aes_cr_reg[0]_1 ),
        .I5(\FSM_sequential_state_reg[1]_1 ),
        .O(\aes_cr_reg[4]_2 ));
  LUT6 #(
    .INIT(64'hFFFF000073400000)) 
    \FSM_sequential_state[1]_i_2 
       (.I0(\FSM_sequential_state_reg[2]_0 ),
        .I1(rk_out_sel_pp1_reg[0]),
        .I2(\FSM_sequential_state[1]_i_5_n_0 ),
        .I3(\FSM_sequential_state[1]_i_6__0_n_0 ),
        .I4(\aes_cr_reg[0]_1 ),
        .I5(\FSM_sequential_state_reg[1]_2 ),
        .O(\FSM_sequential_state[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAEAAAAA)) 
    \FSM_sequential_state[1]_i_2__0 
       (.I0(\FSM_sequential_state[1]_i_3_n_0 ),
        .I1(\aes_cr_reg[0]_1 ),
        .I2(state[1]),
        .I3(state[0]),
        .I4(\FSM_sequential_state[1]_i_4_n_0 ),
        .I5(\FSM_sequential_state[1]_i_5__0_n_0 ),
        .O(\FSM_sequential_state[1]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h000044000F000000)) 
    \FSM_sequential_state[1]_i_3 
       (.I0(state[0]),
        .I1(\FSM_sequential_state[1]_i_6_n_0 ),
        .I2(\FSM_sequential_state[2]_i_4_n_0 ),
        .I3(\aes_cr_reg[0]_1 ),
        .I4(state[2]),
        .I5(state[1]),
        .O(\FSM_sequential_state[1]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair285" *) 
  LUT5 #(
    .INIT(32'hFFFFBFFF)) 
    \FSM_sequential_state[1]_i_4 
       (.I0(enable_i[2]),
        .I1(enable_i[1]),
        .I2(Q[0]),
        .I3(Q[1]),
        .I4(\KR[1].key_host_reg[2][0] ),
        .O(\FSM_sequential_state[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h2FFF00002F2F0000)) 
    \FSM_sequential_state[1]_i_5 
       (.I0(\aes_cr_reg[7]_0 [5]),
        .I1(\aes_cr_reg[7]_0 [4]),
        .I2(\aes_cr_reg[7]_0 [3]),
        .I3(rk_out_sel_pp1_reg[3]),
        .I4(rk_out_sel_pp1_reg[2]),
        .I5(\aes_cr_reg[7]_0 [2]),
        .O(\FSM_sequential_state[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000808800000000)) 
    \FSM_sequential_state[1]_i_5__0 
       (.I0(state[2]),
        .I1(\aes_cr_reg[0]_1 ),
        .I2(enable_i[4]),
        .I3(enable_i[0]),
        .I4(state[0]),
        .I5(state[1]),
        .O(\FSM_sequential_state[1]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair288" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \FSM_sequential_state[1]_i_6 
       (.I0(enable_i[0]),
        .I1(enable_i[4]),
        .O(\FSM_sequential_state[1]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT5 #(
    .INIT(32'h10001010)) 
    \FSM_sequential_state[1]_i_6__0 
       (.I0(rk_out_sel_pp1_reg[3]),
        .I1(rk_out_sel_pp1_reg[2]),
        .I2(\aes_cr_reg[7]_0 [3]),
        .I3(\aes_cr_reg[7]_0 [4]),
        .I4(\aes_cr_reg[7]_0 [5]),
        .O(\FSM_sequential_state[1]_i_6__0_n_0 ));
  LUT5 #(
    .INIT(32'h337F3FFF)) 
    \FSM_sequential_state[2]_i_1 
       (.I0(\FSM_sequential_state_reg[0]_2 ),
        .I1(\aes_cr_reg[0]_1 ),
        .I2(state[0]),
        .I3(state[2]),
        .I4(state[1]),
        .O(\FSM_sequential_state[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hC000C000E0A00000)) 
    \FSM_sequential_state[2]_i_2 
       (.I0(\FSM_sequential_state[2]_i_4_n_0 ),
        .I1(\aes_cr_reg[4]_1 ),
        .I2(\aes_cr_reg[0]_1 ),
        .I3(state[0]),
        .I4(state[2]),
        .I5(state[1]),
        .O(\FSM_sequential_state[2]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hDFFF)) 
    \FSM_sequential_state[2]_i_4 
       (.I0(enable_i[5]),
        .I1(\cnt_reg[0]_0 ),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(\FSM_sequential_state[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h88000000C0000000)) 
    \FSM_sequential_state[2]_i_4__0 
       (.I0(\aes_cr_reg[7]_0 [3]),
        .I1(\aes_cr_reg[5]_0 ),
        .I2(\aes_cr_reg[7]_0 [2]),
        .I3(rk_out_sel_pp1_reg[0]),
        .I4(rk_out_sel_pp1_reg[2]),
        .I5(rk_out_sel_pp1_reg[3]),
        .O(\aes_cr_reg[4]_3 ));
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \FSM_sequential_state[2]_i_5 
       (.I0(\aes_cr_reg[7]_0 [3]),
        .I1(\aes_cr_reg[7]_0 [2]),
        .O(\aes_cr_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h00200020FFFF0000)) 
    \FSM_sequential_state[3]_i_3 
       (.I0(\aes_cr_reg[7]_0 [2]),
        .I1(\aes_cr_reg[7]_0 [3]),
        .I2(\aes_cr_reg[5]_0 ),
        .I3(\IV_BKP_REGISTERS[3].iv_reg[3][0] ),
        .I4(rk_out_sel_pp1_reg[0]),
        .I5(rk_out_sel_pp1_reg[1]),
        .O(\aes_cr_reg[3]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT5 #(
    .INIT(32'h2FFF0000)) 
    \FSM_sequential_state[3]_i_6 
       (.I0(\aes_cr_reg[7]_0 [5]),
        .I1(\aes_cr_reg[7]_0 [4]),
        .I2(\aes_cr_reg[7]_0 [3]),
        .I3(rk_out_sel_pp1_reg[0]),
        .I4(rk_out_sel_pp1_reg[1]),
        .O(\aes_cr_reg[6]_1 ));
  (* FSM_ENCODED_STATES = "WAIT:011,START:001,IDLE:000,OUTPUT:100,INPUT:010" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_state_reg[0] 
       (.C(clk_i),
        .CE(\FSM_sequential_state[2]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\FSM_sequential_state[0]_i_1_n_0 ),
        .Q(state[0]));
  (* FSM_ENCODED_STATES = "WAIT:011,START:001,IDLE:000,OUTPUT:100,INPUT:010" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_state_reg[1] 
       (.C(clk_i),
        .CE(\FSM_sequential_state[2]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\FSM_sequential_state[1]_i_1_n_0 ),
        .Q(state[1]));
  (* FSM_ENCODED_STATES = "WAIT:011,START:001,IDLE:000,OUTPUT:100,INPUT:010" *) 
  FDCE #(
    .INIT(1'b0)) 
    \FSM_sequential_state_reg[2] 
       (.C(clk_i),
        .CE(\FSM_sequential_state[2]_i_1_n_0 ),
        .CLR(rst_i),
        .D(\FSM_sequential_state[2]_i_2_n_0 ),
        .Q(state[2]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][0]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [0]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[0]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[0].bkp[0][10]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [18]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[2]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][10]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[0].bkp[0][10]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][15] [2]));
  (* SOFT_HLUTNM = "soft_lutpair311" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][10]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [10]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][10]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[0].bkp[0][11]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [19]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[3]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][11]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[0].bkp[0][11]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][15] [3]));
  (* SOFT_HLUTNM = "soft_lutpair311" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][11]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [11]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[0].bkp[0][12]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [20]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[4]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][12]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[0].bkp[0][12]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][15] [4]));
  (* SOFT_HLUTNM = "soft_lutpair310" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][12]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [12]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[0].bkp[0][13]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [21]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[5]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][13]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[0].bkp[0][13]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][15] [5]));
  (* SOFT_HLUTNM = "soft_lutpair310" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][13]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [13]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[0].bkp[0][14]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [22]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[6]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][14]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[0].bkp[0][14]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][15] [6]));
  (* SOFT_HLUTNM = "soft_lutpair309" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][14]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [14]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[0].bkp[0][15]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [23]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[7]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][15]_i_5_n_0 ),
        .I5(\IV_BKP_REGISTERS[0].bkp[0][15]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][15] [7]));
  (* SOFT_HLUTNM = "soft_lutpair309" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][15]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [15]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][15]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][16]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [16]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[16]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][16] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][17]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [17]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[17]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][17] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][18]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [18]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[18]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][18] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][19]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [19]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[19]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][19] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][1]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [1]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[1]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][1] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][20]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [20]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[20]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][20] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][21]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [21]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[21]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][21] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][22]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [22]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[22]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][22] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][23]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [23]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[23]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][23] ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[0].bkp[0][24]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[24]),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [24]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_17 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[0].bkp[0][25]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[25]),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [25]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_19 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[0].bkp[0][26]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[26]),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [26]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_21 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[0].bkp[0][27]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[27]),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [27]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_23 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[0].bkp[0][28]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[28]),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [28]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_25 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[0].bkp[0][29]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[29]),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [29]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_27 ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][2]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [2]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[2]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][2] ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[0].bkp[0][30]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[30]),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [30]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_29 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[0].bkp[0][31]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[31]),
        .I3(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [31]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_31 ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][3]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [3]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[3]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][3] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][4]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [4]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[4]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][4] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][5]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [5]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[5]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][5] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][6]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [6]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[6]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][6] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[0].bkp[0][7]_i_2 
       (.I0(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [7]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[7]),
        .O(\IV_BKP_REGISTERS[0].bkp_1_reg[0][7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[0].bkp[0][8]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [16]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[0]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][8]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[0].bkp[0][8]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][15] [0]));
  (* SOFT_HLUTNM = "soft_lutpair312" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][8]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [8]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[0].bkp[0][9]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [17]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][9]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[0].bkp[0][9]_i_2_n_0 ),
        .O(\CD[2].col_reg[1][15] [1]));
  (* SOFT_HLUTNM = "soft_lutpair312" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[0].bkp[0][9]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[0].bkp_reg[0][31] [9]),
        .O(\IV_BKP_REGISTERS[0].bkp[0][9]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h888F888888888888)) 
    \IV_BKP_REGISTERS[0].bkp_1[0][31]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][0] [0]),
        .I1(\IV_BKP_REGISTERS[3].bkp_1[3][31]_i_2_n_0 ),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\FSM_sequential_state_reg[0]_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_1[3][31]_i_3_n_0 ),
        .O(\col_en_cnt_unit_pp2_reg[0] ));
  (* SOFT_HLUTNM = "soft_lutpair279" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \IV_BKP_REGISTERS[0].iv[0][31]_i_1 
       (.I0(enable_i[5]),
        .I1(enable_i[6]),
        .I2(enable_i[0]),
        .I3(enable_i[4]),
        .I4(enable_i_2_sn_1),
        .O(iv_en[0]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][0]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [0]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[0]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][0] ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[1].bkp[1][10]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[10]),
        .I3(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [10]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_6 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[1].bkp[1][11]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[11]),
        .I3(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [11]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_8 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[1].bkp[1][12]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[12]),
        .I3(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [12]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_10 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[1].bkp[1][13]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[13]),
        .I3(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [13]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_12 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[1].bkp[1][14]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[14]),
        .I3(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [14]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_14 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[1].bkp[1][15]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[15]),
        .I3(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [15]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_16 ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][16]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [16]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[16]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][16] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][17]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [17]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[17]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][17] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][18]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [18]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[18]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][18] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][19]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [19]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[19]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][19] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][1]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [1]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[1]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][1] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][20]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [20]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[20]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][20] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][21]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [21]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[21]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][21] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][22]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [22]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[22]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][22] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][23]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [23]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[23]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][23] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[1].bkp[1][24]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [8]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[8]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][24]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[1].bkp[1][24]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [0]));
  (* SOFT_HLUTNM = "soft_lutpair308" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][24]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [24]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][24]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[1].bkp[1][25]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [9]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[9]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][25]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[1].bkp[1][25]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [1]));
  (* SOFT_HLUTNM = "soft_lutpair308" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][25]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [25]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][25]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[1].bkp[1][26]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [10]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[10]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][26]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[1].bkp[1][26]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [2]));
  (* SOFT_HLUTNM = "soft_lutpair307" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][26]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [26]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][26]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[1].bkp[1][27]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [11]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[11]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][27]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[1].bkp[1][27]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [3]));
  (* SOFT_HLUTNM = "soft_lutpair307" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][27]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [27]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[1].bkp[1][28]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [12]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[12]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][28]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[1].bkp[1][28]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [4]));
  (* SOFT_HLUTNM = "soft_lutpair306" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][28]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [28]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][28]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[1].bkp[1][29]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [13]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[13]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][29]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[1].bkp[1][29]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [5]));
  (* SOFT_HLUTNM = "soft_lutpair306" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][29]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [29]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][29]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][2]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [2]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[2]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[1].bkp[1][30]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [14]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[14]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][30]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[1].bkp[1][30]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [6]));
  (* SOFT_HLUTNM = "soft_lutpair305" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][30]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [30]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][30]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[1].bkp[1][31]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [15]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[15]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][31]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[1].bkp[1][31]_i_2_n_0 ),
        .O(\CD[1].col_reg[2][31] [7]));
  (* SOFT_HLUTNM = "soft_lutpair305" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[1].bkp[1][31]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [31]),
        .O(\IV_BKP_REGISTERS[1].bkp[1][31]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][3]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [3]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[3]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][3] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][4]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [4]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[4]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][4] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][5]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [5]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[5]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][5] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][6]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [6]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[6]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][6] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[1].bkp[1][7]_i_2 
       (.I0(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [7]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[7]),
        .O(\IV_BKP_REGISTERS[1].bkp_1_reg[1][7] ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[1].bkp[1][8]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[8]),
        .I3(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [8]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_2 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[1].bkp[1][9]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[9]),
        .I3(\IV_BKP_REGISTERS[1].bkp_reg[1][31] [9]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_4 ));
  LUT6 #(
    .INIT(64'h8F88888888888888)) 
    \IV_BKP_REGISTERS[1].bkp_1[1][31]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][0] [1]),
        .I1(\IV_BKP_REGISTERS[3].bkp_1[3][31]_i_2_n_0 ),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(\FSM_sequential_state_reg[0]_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_1[3][31]_i_3_n_0 ),
        .O(\col_en_cnt_unit_pp2_reg[1] ));
  (* SOFT_HLUTNM = "soft_lutpair279" *) 
  LUT5 #(
    .INIT(32'h40000000)) 
    \IV_BKP_REGISTERS[1].iv[1][31]_i_1 
       (.I0(enable_i[0]),
        .I1(enable_i[4]),
        .I2(enable_i[5]),
        .I3(enable_i[6]),
        .I4(enable_i_2_sn_1),
        .O(iv_en[1]));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \IV_BKP_REGISTERS[1].iv[1][31]_i_2 
       (.I0(enable_i[2]),
        .I1(enable_i[1]),
        .I2(enable_i[3]),
        .I3(state[0]),
        .I4(state[1]),
        .I5(state[2]),
        .O(enable_i_2_sn_1));
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][0]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [0]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[0]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][0] ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[2].bkp[2][10]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[10]),
        .I3(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [10]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_5 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[2].bkp[2][11]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[11]),
        .I3(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [11]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_7 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[2].bkp[2][12]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[12]),
        .I3(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [12]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_9 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[2].bkp[2][13]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[13]),
        .I3(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [13]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_11 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[2].bkp[2][14]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[14]),
        .I3(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [14]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_13 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[2].bkp[2][15]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[15]),
        .I3(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [15]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_15 ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][16]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [16]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[16]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][16] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][17]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [17]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[17]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][17] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][18]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [18]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[18]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][18] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][19]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [19]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[19]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][19] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][1]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [1]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[1]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][1] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][20]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [20]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[20]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][20] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][21]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [21]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[21]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][21] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][22]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [22]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[22]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][22] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][23]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [23]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[23]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][23] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][24]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [24]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[8]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][24]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[2].bkp[2][24]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [0]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][24]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [8]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[24]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][24]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair304" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][24]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [24]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][24]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][25]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [25]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[9]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][25]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[2].bkp[2][25]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [1]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][25]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [9]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[25]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][25]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair304" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][25]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [25]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][25]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][26]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [26]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[10]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][26]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[2].bkp[2][26]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [2]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][26]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [10]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[26]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][26]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair303" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][26]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [26]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][26]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][27]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [27]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[11]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][27]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[2].bkp[2][27]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [3]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][27]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [11]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[27]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][27]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair303" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][27]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [27]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][27]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][28]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [28]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[12]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][28]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[2].bkp[2][28]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [4]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][28]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [12]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[28]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][28]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair302" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][28]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [28]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][28]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][29]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [29]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[13]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][29]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[2].bkp[2][29]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [5]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][29]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [13]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[29]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][29]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair302" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][29]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [29]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][29]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][2]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [2]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[2]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][30]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [30]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[14]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][30]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[2].bkp[2][30]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [6]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][30]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [14]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[30]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][30]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair301" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][30]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [30]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][30]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[2].bkp[2][31]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [31]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[15]),
        .I4(\IV_BKP_REGISTERS[2].bkp[2][31]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[2].bkp[2][31]_i_4_n_0 ),
        .O(\CD[2].col_reg[1][31] [7]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][31]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [15]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[31]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][31]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair301" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[2].bkp[2][31]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [31]),
        .O(\IV_BKP_REGISTERS[2].bkp[2][31]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][3]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [3]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[3]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][3] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][4]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [4]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[4]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][4] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][5]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [5]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[5]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][5] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][6]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [6]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[6]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][6] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[2].bkp[2][7]_i_2 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [7]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[7]),
        .O(\IV_BKP_REGISTERS[2].bkp_1_reg[2][7] ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[2].bkp[2][8]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[8]),
        .I3(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [8]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_1 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[2].bkp[2][9]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[9]),
        .I3(\IV_BKP_REGISTERS[2].bkp_reg[2][31] [9]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_3 ));
  LUT6 #(
    .INIT(64'h8F88888888888888)) 
    \IV_BKP_REGISTERS[2].bkp_1[2][31]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][0] [2]),
        .I1(\IV_BKP_REGISTERS[3].bkp_1[3][31]_i_2_n_0 ),
        .I2(Q[0]),
        .I3(Q[1]),
        .I4(\FSM_sequential_state_reg[0]_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp_1[3][31]_i_3_n_0 ),
        .O(\col_en_cnt_unit_pp2_reg[2] ));
  (* SOFT_HLUTNM = "soft_lutpair288" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \IV_BKP_REGISTERS[2].iv[2][31]_i_1 
       (.I0(enable_i[5]),
        .I1(enable_i[6]),
        .I2(enable_i[0]),
        .I3(enable_i[4]),
        .I4(enable_i_1_sn_1),
        .O(iv_en[2]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][0]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [0]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[0]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[3].bkp[3][10]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [2]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[2]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][10]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp[3][10]_i_4_n_0 ),
        .O(D[2]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][10]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [2]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[10]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][10]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair300" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][10]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [10]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][10]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[3].bkp[3][11]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [3]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[3]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][11]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp[3][11]_i_4_n_0 ),
        .O(D[3]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][11]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [3]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[11]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][11]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair299" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][11]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [11]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][11]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[3].bkp[3][12]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [4]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[4]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][12]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp[3][12]_i_4_n_0 ),
        .O(D[4]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][12]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [4]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[12]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][12]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair298" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][12]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [12]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][12]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[3].bkp[3][13]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [5]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[5]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][13]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp[3][13]_i_4_n_0 ),
        .O(D[5]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][13]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [5]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[13]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][13]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair298" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][13]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [13]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[3].bkp[3][14]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [6]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[6]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][14]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp[3][14]_i_4_n_0 ),
        .O(D[6]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][14]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [6]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[14]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][14]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair297" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][14]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [14]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[3].bkp[3][15]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [7]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[7]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][15]_i_5_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp[3][15]_i_6_n_0 ),
        .O(D[7]));
  LUT6 #(
    .INIT(64'h2202020200000000)) 
    \IV_BKP_REGISTERS[3].bkp[3][15]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(\aes_cr_reg[7]_0 [3]),
        .I3(rk_out_sel_pp1_reg[1]),
        .I4(rk_out_sel_pp1_reg[2]),
        .I5(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_2 ),
        .O(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][15]_i_5 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [7]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[15]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][15]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair297" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][15]_i_6 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [15]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][15]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][16]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [16]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[16]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][16] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][17]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [17]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[17]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][17] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][18]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [18]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[18]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][18] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][19]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [19]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[19]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][19] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][1]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [1]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[1]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][1] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][20]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [20]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[20]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][20] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][21]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [21]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[21]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][21] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][22]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [22]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[22]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][22] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][23]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [23]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[23]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][23] ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[3].bkp[3][24]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[24]),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [24]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_18 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[3].bkp[3][25]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[25]),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [25]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_20 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[3].bkp[3][26]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[26]),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [26]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_22 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[3].bkp[3][27]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[27]),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [27]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_24 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[3].bkp[3][28]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[28]),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [28]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_26 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[3].bkp[3][29]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[29]),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [29]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_28 ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][2]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [2]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[2]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][2] ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[3].bkp[3][30]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[30]),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [30]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_30 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \IV_BKP_REGISTERS[3].bkp[3][31]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(bus_swap[31]),
        .I3(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [31]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .O(\aes_cr_reg[5]_32 ));
  (* SOFT_HLUTNM = "soft_lutpair286" *) 
  LUT5 #(
    .INIT(32'h008F0000)) 
    \IV_BKP_REGISTERS[3].bkp[3][31]_i_4 
       (.I0(rk_out_sel_pp1_reg[2]),
        .I1(rk_out_sel_pp1_reg[1]),
        .I2(\aes_cr_reg[7]_0 [3]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(\aes_cr_reg[7]_0 [4]),
        .O(\FSM_sequential_state_reg[2]_4 ));
  LUT5 #(
    .INIT(32'h9BBB9999)) 
    \IV_BKP_REGISTERS[3].bkp[3][31]_i_6 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(rk_out_sel_pp1_reg[2]),
        .I3(rk_out_sel_pp1_reg[1]),
        .I4(\aes_cr_reg[7]_0 [3]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][3]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [3]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[3]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][3] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][4]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [4]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[4]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][4] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][5]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [5]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[5]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][5] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][6]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [6]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[6]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][6] ));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][7]_i_2 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [7]),
        .I1(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[7]),
        .O(\IV_BKP_REGISTERS[3].bkp_1_reg[3][7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[3].bkp[3][8]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [0]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[0]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][8]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp[3][8]_i_4_n_0 ),
        .O(D[0]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][8]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [0]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[8]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][8]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair300" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][8]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [8]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][8]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \IV_BKP_REGISTERS[3].bkp[3][9]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][15]_i_2_n_0 ),
        .I1(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_0 [1]),
        .I2(\IV_BKP_REGISTERS[0].bkp_reg[0][8] ),
        .I3(data_in[1]),
        .I4(\IV_BKP_REGISTERS[3].bkp[3][9]_i_3_n_0 ),
        .I5(\IV_BKP_REGISTERS[3].bkp[3][9]_i_4_n_0 ),
        .O(D[1]));
  LUT5 #(
    .INIT(32'h8F888888)) 
    \IV_BKP_REGISTERS[3].bkp[3][9]_i_3 
       (.I0(\IV_BKP_REGISTERS[2].bkp_reg[2][31]_1 [1]),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][8] ),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(bus_swap[9]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][9]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair299" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \IV_BKP_REGISTERS[3].bkp[3][9]_i_4 
       (.I0(\IV_BKP_REGISTERS[3].bkp[3][31]_i_6_n_0 ),
        .I1(\IV_BKP_REGISTERS[3].bkp_reg[3][31] [9]),
        .O(\IV_BKP_REGISTERS[3].bkp[3][9]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF888888888888888)) 
    \IV_BKP_REGISTERS[3].bkp_1[3][31]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].bkp_reg[3][0] [3]),
        .I1(\IV_BKP_REGISTERS[3].bkp_1[3][31]_i_2_n_0 ),
        .I2(\FSM_sequential_state_reg[0]_0 ),
        .I3(Q[1]),
        .I4(Q[0]),
        .I5(\IV_BKP_REGISTERS[3].bkp_1[3][31]_i_3_n_0 ),
        .O(\col_en_cnt_unit_pp2_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0000000020002222)) 
    \IV_BKP_REGISTERS[3].bkp_1[3][31]_i_2 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(rk_out_sel_pp1_reg[2]),
        .I3(rk_out_sel_pp1_reg[1]),
        .I4(\aes_cr_reg[7]_0 [3]),
        .I5(\IV_BKP_REGISTERS[3].iv_reg[3][0] ),
        .O(\IV_BKP_REGISTERS[3].bkp_1[3][31]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair276" *) 
  LUT5 #(
    .INIT(32'h0070FF00)) 
    \IV_BKP_REGISTERS[3].bkp_1[3][31]_i_3 
       (.I0(rk_out_sel_pp1_reg[2]),
        .I1(rk_out_sel_pp1_reg[1]),
        .I2(\aes_cr_reg[7]_0 [3]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(\aes_cr_reg[7]_0 [4]),
        .O(\IV_BKP_REGISTERS[3].bkp_1[3][31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h88888F8888888888)) 
    \IV_BKP_REGISTERS[3].iv[3][31]_i_1 
       (.I0(\IV_BKP_REGISTERS[3].iv_reg[3][0]_0 ),
        .I1(enable_i_1_sn_1),
        .I2(\aes_cr_reg[7]_0 [4]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(\IV_BKP_REGISTERS[3].iv_reg[3][0] ),
        .I5(\IV_BKP_REGISTERS[3].iv_reg[3][0]_1 ),
        .O(\aes_cr_reg[5]_33 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \IV_BKP_REGISTERS[3].iv[3][31]_i_4 
       (.I0(enable_i[1]),
        .I1(state[2]),
        .I2(state[1]),
        .I3(state[0]),
        .I4(enable_i[2]),
        .I5(enable_i[3]),
        .O(enable_i_1_sn_1));
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \KR[0].key[3][31]_i_4 
       (.I0(state[2]),
        .I1(state[1]),
        .I2(state[0]),
        .O(\FSM_sequential_state_reg[2]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair295" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \KR[0].key_host[3][31]_i_1 
       (.I0(key_en[3]),
        .I1(key_derivation_en),
        .O(E));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \KR[0].key_host[3][31]_i_3 
       (.I0(\aes_cr_reg[0]_3 ),
        .I1(enable_i[2]),
        .I2(enable_i[1]),
        .I3(state[2]),
        .I4(state[1]),
        .I5(state[0]),
        .O(key_en[3]));
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    \KR[0].key_host[3][31]_i_4 
       (.I0(\aes_cr_reg[5]_0 ),
        .I1(\aes_cr_reg[7]_0 [3]),
        .I2(\aes_cr_reg[7]_0 [2]),
        .I3(\KR[0].key_host_reg[3][0] ),
        .I4(rk_out_sel_pp1_reg[3]),
        .I5(rk_out_sel_pp1_reg[2]),
        .O(key_derivation_en));
  (* SOFT_HLUTNM = "soft_lutpair296" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \KR[1].key_host[2][31]_i_1 
       (.I0(key_en[2]),
        .I1(key_derivation_en),
        .O(\enable_i[4] ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \KR[1].key_host[2][31]_i_3 
       (.I0(\KR[1].key_host_reg[2][0] ),
        .I1(enable_i[4]),
        .I2(enable_i[0]),
        .I3(enable_i[2]),
        .I4(enable_i[1]),
        .I5(access_permission),
        .O(key_en[2]));
  (* SOFT_HLUTNM = "soft_lutpair295" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \KR[2].key_host[1][31]_i_1 
       (.I0(key_en[1]),
        .I1(key_derivation_en),
        .O(\FSM_sequential_state_reg[2]_5 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \KR[2].key_host[1][31]_i_3 
       (.I0(state[2]),
        .I1(state[1]),
        .I2(state[0]),
        .I3(enable_i[1]),
        .I4(enable_i[2]),
        .I5(\aes_cr_reg[0]_3 ),
        .O(key_en[1]));
  (* SOFT_HLUTNM = "soft_lutpair296" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \KR[3].key_host[0][31]_i_1 
       (.I0(key_en[0]),
        .I1(key_derivation_en),
        .O(\enable_i[2]_1 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \KR[3].key_host[0][31]_i_3 
       (.I0(access_permission),
        .I1(enable_i[2]),
        .I2(enable_i[1]),
        .I3(enable_i[4]),
        .I4(enable_i[0]),
        .I5(\KR[1].key_host_reg[2][0] ),
        .O(key_en[0]));
  LUT6 #(
    .INIT(64'hCCCCCCC800000008)) 
    \aes_cr[0]_i_1 
       (.I0(enable_i[0]),
        .I1(\aes_cr[0]_i_2_n_0 ),
        .I2(enable_i[1]),
        .I3(enable_i[2]),
        .I4(\aes_cr_reg[0]_3 ),
        .I5(\aes_cr_reg[0]_1 ),
        .O(\aes_cr[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFDFFF)) 
    \aes_cr[0]_i_2 
       (.I0(state[1]),
        .I1(\aes_cr_reg[7]_0 [3]),
        .I2(\aes_cr_reg[7]_0 [2]),
        .I3(state[0]),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(state[2]),
        .O(\aes_cr[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \aes_cr[10]_i_1 
       (.I0(state[0]),
        .I1(state[1]),
        .I2(state[2]),
        .I3(enable_i[1]),
        .I4(enable_i[2]),
        .I5(\aes_cr_reg[0]_3 ),
        .O(aes_cr1));
  LUT4 #(
    .INIT(16'hDF00)) 
    \aes_cr[3]_i_1 
       (.I0(enable_i[6]),
        .I1(enable_i[5]),
        .I2(enable_i[4]),
        .I3(enable_i[3]),
        .O(p_1_in__0));
  FDCE #(
    .INIT(1'b0)) 
    \aes_cr_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(\aes_cr[0]_i_1_n_0 ),
        .Q(\aes_cr_reg[0]_1 ));
  FDCE #(
    .INIT(1'b0)) 
    \aes_cr_reg[10] 
       (.C(clk_i),
        .CE(aes_cr1),
        .CLR(rst_i),
        .D(enable_i[11]),
        .Q(dma_out_en));
  FDCE #(
    .INIT(1'b0)) 
    \aes_cr_reg[1] 
       (.C(clk_i),
        .CE(aes_cr1),
        .CLR(rst_i),
        .D(enable_i[1]),
        .Q(\aes_cr_reg[7]_0 [0]));
  FDCE #(
    .INIT(1'b0)) 
    \aes_cr_reg[2] 
       (.C(clk_i),
        .CE(aes_cr1),
        .CLR(rst_i),
        .D(enable_i[2]),
        .Q(\aes_cr_reg[7]_0 [1]));
  FDCE #(
    .INIT(1'b0)) 
    \aes_cr_reg[3] 
       (.C(clk_i),
        .CE(aes_cr1),
        .CLR(rst_i),
        .D(p_1_in__0),
        .Q(\aes_cr_reg[7]_0 [2]));
  FDCE #(
    .INIT(1'b0)) 
    \aes_cr_reg[4] 
       (.C(clk_i),
        .CE(aes_cr1),
        .CLR(rst_i),
        .D(enable_i[4]),
        .Q(\aes_cr_reg[7]_0 [3]));
  FDCE #(
    .INIT(1'b0)) 
    \aes_cr_reg[5] 
       (.C(clk_i),
        .CE(aes_cr1),
        .CLR(rst_i),
        .D(enable_i[5]),
        .Q(\aes_cr_reg[7]_0 [4]));
  FDCE #(
    .INIT(1'b0)) 
    \aes_cr_reg[6] 
       (.C(clk_i),
        .CE(aes_cr1),
        .CLR(rst_i),
        .D(enable_i[6]),
        .Q(\aes_cr_reg[7]_0 [5]));
  FDCE #(
    .INIT(1'b0)) 
    \aes_cr_reg[7] 
       (.C(clk_i),
        .CE(aes_cr1),
        .CLR(rst_i),
        .D(enable_i[8]),
        .Q(\aes_cr_reg[7]_0 [6]));
  FDCE #(
    .INIT(1'b0)) 
    \aes_cr_reg[8] 
       (.C(clk_i),
        .CE(aes_cr1),
        .CLR(rst_i),
        .D(enable_i[9]),
        .Q(err_ie));
  FDCE #(
    .INIT(1'b0)) 
    \aes_cr_reg[9] 
       (.C(clk_i),
        .CE(aes_cr1),
        .CLR(rst_i),
        .D(enable_i[10]),
        .Q(dma_in_en));
  (* SOFT_HLUTNM = "soft_lutpair276" *) 
  LUT5 #(
    .INIT(32'h8FFF8F8F)) 
    \base_new_pp[7]_i_10 
       (.I0(rk_out_sel_pp1_reg[2]),
        .I1(rk_out_sel_pp1_reg[1]),
        .I2(\aes_cr_reg[7]_0 [3]),
        .I3(\aes_cr_reg[7]_0 [4]),
        .I4(\aes_cr_reg[7]_0 [5]),
        .O(enc_dec));
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    ccf_i_3
       (.I0(\aes_cr_reg[0]_3 ),
        .I1(enable_i[2]),
        .I2(enable_i[1]),
        .O(\enable_i[2]_0 ));
  FDCE #(
    .INIT(1'b0)) 
    ccf_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(ccf_reg_0),
        .Q(ccf));
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT5 #(
    .INIT(32'h5755FFFF)) 
    \cnt[0]_i_1 
       (.I0(\aes_cr_reg[0]_1 ),
        .I1(state[2]),
        .I2(state[1]),
        .I3(state[0]),
        .I4(Q[0]),
        .O(\cnt[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFEFEFFFE)) 
    \cnt[1]_i_1 
       (.I0(\cnt[1]_i_3_n_0 ),
        .I1(\FSM_sequential_state_reg[0]_0 ),
        .I2(\cnt[1]_i_4_n_0 ),
        .I3(state[0]),
        .I4(\FSM_sequential_state_reg[0]_2 ),
        .I5(state[2]),
        .O(\cnt[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h6F6F6FFF6F6F6F6F)) 
    \cnt[1]_i_2 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(\aes_cr_reg[0]_1 ),
        .I3(state[2]),
        .I4(state[1]),
        .I5(state[0]),
        .O(\cnt[1]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT4 #(
    .INIT(16'h02FF)) 
    \cnt[1]_i_3 
       (.I0(state[0]),
        .I1(state[1]),
        .I2(state[2]),
        .I3(\aes_cr_reg[0]_1 ),
        .O(\cnt[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00FF000045454545)) 
    \cnt[1]_i_4 
       (.I0(state[1]),
        .I1(\aes_cr_reg[7]_0 [3]),
        .I2(\aes_cr_reg[7]_0 [2]),
        .I3(\cnt_reg[0]_0 ),
        .I4(enable_i[5]),
        .I5(state[2]),
        .O(\cnt[1]_i_4_n_0 ));
  FDPE #(
    .INIT(1'b1)) 
    \cnt_reg[0] 
       (.C(clk_i),
        .CE(\cnt[1]_i_1_n_0 ),
        .D(\cnt[0]_i_1_n_0 ),
        .PRE(rst_i),
        .Q(Q[0]));
  FDPE #(
    .INIT(1'b1)) 
    \cnt_reg[1] 
       (.C(clk_i),
        .CE(\cnt[1]_i_1_n_0 ),
        .D(\cnt[1]_i_2_n_0 ),
        .PRE(rst_i),
        .Q(Q[1]));
  (* SOFT_HLUTNM = "soft_lutpair287" *) 
  LUT3 #(
    .INIT(8'h2F)) 
    \col_en_cnt_unit_pp1[3]_i_3 
       (.I0(\aes_cr_reg[7]_0 [5]),
        .I1(\aes_cr_reg[7]_0 [4]),
        .I2(\aes_cr_reg[7]_0 [3]),
        .O(\aes_cr_reg[6]_2 ));
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT3 #(
    .INIT(8'h2C)) 
    \col_sel_pp1[1]_i_2 
       (.I0(\aes_cr_reg[7]_0 [3]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(\aes_cr_reg[7]_0 [4]),
        .O(\aes_cr_reg[4]_4 ));
  FDCE #(
    .INIT(1'b0)) 
    dma_req_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(Q[0]),
        .Q(dma_req));
  (* SOFT_HLUTNM = "soft_lutpair292" *) 
  LUT4 #(
    .INIT(16'hA8AB)) 
    first_block_i_1
       (.I0(first_block),
        .I1(state[0]),
        .I2(state[1]),
        .I3(state[2]),
        .O(first_block_i_1_n_0));
  FDPE #(
    .INIT(1'b1)) 
    first_block_reg
       (.C(clk_i),
        .CE(1'b1),
        .D(first_block_i_1_n_0),
        .PRE(rst_i),
        .Q(first_block));
  LUT5 #(
    .INIT(32'h00001011)) 
    \info_o[0]_INST_0_i_7 
       (.I0(enable_i[1]),
        .I1(enable_i[2]),
        .I2(ccf),
        .I3(enable_i[5]),
        .I4(\info_o[0]_INST_0_i_4 ),
        .O(\enable_i[1]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[10]_INST_0_i_3 
       (.I0(\info_o[12] [3]),
        .I1(\aes_cr_reg[0]_0 ),
        .I2(err_ie),
        .I3(\info_o[3]_0 ),
        .O(\aes_cr_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[11]_INST_0_i_3 
       (.I0(\info_o[12] [4]),
        .I1(\aes_cr_reg[0]_0 ),
        .I2(dma_in_en),
        .I3(\info_o[3]_0 ),
        .O(\aes_cr_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[12]_INST_0_i_3 
       (.I0(\info_o[12] [5]),
        .I1(\aes_cr_reg[0]_0 ),
        .I2(dma_out_en),
        .I3(\info_o[3]_0 ),
        .O(\aes_cr_reg[10]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair289" *) 
  LUT5 #(
    .INIT(32'hE0000000)) 
    \info_o[1]_INST_0 
       (.I0(state[0]),
        .I1(state[1]),
        .I2(\info_o[3] [0]),
        .I3(err_ie),
        .I4(info_o_1_sn_1),
        .O(info_o[0]));
  LUT4 #(
    .INIT(16'hA888)) 
    \info_o[2]_INST_0 
       (.I0(\info_o[2]_INST_0_i_1_n_0 ),
        .I1(\info_o[2]_INST_0_i_2_n_0 ),
        .I2(info_o_1_sn_1),
        .I3(\info_o[3] [1]),
        .O(info_o[1]));
  LUT6 #(
    .INIT(64'h0000100010000000)) 
    \info_o[2]_INST_0_i_1 
       (.I0(state[0]),
        .I1(state[2]),
        .I2(\aes_cr_reg[0]_1 ),
        .I3(dma_in_en),
        .I4(Q[0]),
        .I5(dma_req),
        .O(\info_o[2]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000AC)) 
    \info_o[2]_INST_0_i_2 
       (.I0(wr_err),
        .I1(\aes_cr_reg[7]_0 [1]),
        .I2(enable_i[0]),
        .I3(enable_i[1]),
        .I4(enable_i[2]),
        .I5(info_o_2_sn_1),
        .O(\info_o[2]_INST_0_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT5 #(
    .INIT(32'h00000004)) 
    \info_o[31]_INST_0_i_27 
       (.I0(enable_i[0]),
        .I1(enable_i[2]),
        .I2(state[0]),
        .I3(state[1]),
        .I4(state[2]),
        .O(key_sel_rd));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \info_o[31]_INST_0_i_29 
       (.I0(\aes_cr_reg[0]_3 ),
        .I1(\info_o[31]_INST_0_i_15 ),
        .I2(state[1]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(\FSM_sequential_state[0]_i_2__0_n_0 ),
        .O(col_en_host[3]));
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \info_o[31]_INST_0_i_3 
       (.I0(\aes_cr_reg[0]_1 ),
        .I1(enable_i[2]),
        .I2(enable_i[3]),
        .I3(enable_i[4]),
        .I4(enable_i[6]),
        .O(\aes_cr_reg[0]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \info_o[31]_INST_0_i_32 
       (.I0(state[2]),
        .I1(Q[0]),
        .I2(state[1]),
        .I3(state[0]),
        .O(\FSM_sequential_state_reg[2]_2 ));
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \info_o[31]_INST_0_i_34 
       (.I0(state[2]),
        .I1(Q[1]),
        .I2(state[1]),
        .I3(state[0]),
        .O(\FSM_sequential_state_reg[2]_3 ));
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \info_o[31]_INST_0_i_39 
       (.I0(state[0]),
        .I1(state[1]),
        .I2(state[2]),
        .I3(enable_i[1]),
        .O(\FSM_sequential_state_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \info_o[31]_INST_0_i_40 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(\aes_cr_reg[0]_3 ),
        .I3(\info_o[31]_INST_0_i_15 ),
        .I4(state[1]),
        .I5(\info_o[31]_INST_0_i_44_n_0 ),
        .O(col_en_host[2]));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \info_o[31]_INST_0_i_42 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(\aes_cr_reg[0]_3 ),
        .I3(\info_o[31]_INST_0_i_15 ),
        .I4(state[1]),
        .I5(\info_o[31]_INST_0_i_44_n_0 ),
        .O(col_en_host[1]));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \info_o[31]_INST_0_i_43 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(\aes_cr_reg[0]_3 ),
        .I3(\info_o[31]_INST_0_i_15 ),
        .I4(state[1]),
        .I5(\info_o[31]_INST_0_i_44_n_0 ),
        .O(col_en_host[0]));
  LUT2 #(
    .INIT(4'hE)) 
    \info_o[31]_INST_0_i_44 
       (.I0(state[0]),
        .I1(state[2]),
        .O(\info_o[31]_INST_0_i_44_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \info_o[31]_INST_0_i_6 
       (.I0(\aes_cr_reg[0]_1 ),
        .I1(enable_i[3]),
        .I2(enable_i[2]),
        .I3(enable_i[6]),
        .I4(enable_i[4]),
        .O(\aes_cr_reg[0]_2 ));
  LUT5 #(
    .INIT(32'hAA808080)) 
    \info_o[3]_INST_0 
       (.I0(\info_o[3]_INST_0_i_1_n_0 ),
        .I1(\info_o[3]_0 ),
        .I2(\aes_cr_reg[7]_0 [2]),
        .I3(info_o_1_sn_1),
        .I4(\info_o[3] [2]),
        .O(info_o[2]));
  LUT6 #(
    .INIT(64'h0000088000000000)) 
    \info_o[3]_INST_0_i_1 
       (.I0(state[2]),
        .I1(\aes_cr_reg[0]_1 ),
        .I2(dma_req),
        .I3(Q[0]),
        .I4(\info_o[3]_INST_0_i_4_n_0 ),
        .I5(dma_out_en),
        .O(\info_o[3]_INST_0_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair289" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \info_o[3]_INST_0_i_4 
       (.I0(state[0]),
        .I1(state[1]),
        .O(\info_o[3]_INST_0_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[4]_INST_0_i_3 
       (.I0(\info_o[12] [0]),
        .I1(\aes_cr_reg[0]_0 ),
        .I2(\aes_cr_reg[7]_0 [3]),
        .I3(\info_o[3]_0 ),
        .O(\aes_cr_reg[4]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[6]_INST_0_i_3 
       (.I0(\info_o[12] [1]),
        .I1(\aes_cr_reg[0]_0 ),
        .I2(\aes_cr_reg[7]_0 [5]),
        .I3(\info_o[3]_0 ),
        .O(\aes_cr_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[9]_INST_0_i_3 
       (.I0(\info_o[12] [2]),
        .I1(\aes_cr_reg[0]_0 ),
        .I2(\aes_cr_reg[7]_0 [6]),
        .I3(\info_o[3]_0 ),
        .O(\aes_cr_reg[7]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \key_en_pp1[3]_i_3 
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .O(\aes_cr_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hF4FFF4FF44FFFFFF)) 
    rk_out_sel_pp1_i_1
       (.I0(\aes_cr_reg[7]_0 [4]),
        .I1(\aes_cr_reg[7]_0 [5]),
        .I2(rk_out_sel_pp1_reg[1]),
        .I3(\aes_cr_reg[7]_0 [3]),
        .I4(rk_out_sel_pp1_reg[3]),
        .I5(rk_out_sel_pp1_reg[2]),
        .O(rk_out_sel));
  (* SOFT_HLUTNM = "soft_lutpair286" *) 
  LUT5 #(
    .INIT(32'hD5D5FFD5)) 
    \sbox_pp2[31]_i_5 
       (.I0(\aes_cr_reg[7]_0 [3]),
        .I1(rk_out_sel_pp1_reg[1]),
        .I2(rk_out_sel_pp1_reg[2]),
        .I3(\aes_cr_reg[7]_0 [5]),
        .I4(\aes_cr_reg[7]_0 [4]),
        .O(\aes_cr_reg[4]_6 ));
  LUT5 #(
    .INIT(32'hEFFFAAAA)) 
    wr_err_i_1
       (.I0(wr_err_en),
        .I1(\enable_i[2]_0 ),
        .I2(access_permission),
        .I3(enable_i[7]),
        .I4(wr_err),
        .O(wr_err_i_1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT5 #(
    .INIT(32'h04040400)) 
    wr_err_i_2
       (.I0(enable_i[2]),
        .I1(enable_i[1]),
        .I2(\aes_cr_reg[0]_3 ),
        .I3(state[2]),
        .I4(state[0]),
        .O(wr_err_en));
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT3 #(
    .INIT(8'h01)) 
    wr_err_i_3
       (.I0(state[2]),
        .I1(state[1]),
        .I2(state[0]),
        .O(access_permission));
  FDCE #(
    .INIT(1'b0)) 
    wr_err_reg
       (.C(clk_i),
        .CE(1'b1),
        .CLR(rst_i),
        .D(wr_err_i_1_n_0),
        .Q(wr_err));
endmodule

(* ORIG_REF_NAME = "sBox" *) 
module switch_elements_sBox
   (enable_i_0_sp_1,
    \round_pp1_reg[0] ,
    \round_pp1_reg[3] ,
    \round_pp1_reg[3]_0 ,
    \round_pp1_reg[0]_0 ,
    \round_pp1_reg[3]_1 ,
    D,
    \round_pp1_reg[0]_1 ,
    \base_new_pp_reg[4] ,
    sbox_out_enc,
    \base_new_pp_reg[6] ,
    \base_new_pp_reg[4]_0 ,
    \base_new_pp_reg[6]_0 ,
    \base_new_pp_reg[6]_1 ,
    \base_new_pp_reg[1] ,
    \base_new_pp_reg[4]_1 ,
    \base_new_pp_reg[6]_2 ,
    \base_new_pp_reg[4]_2 ,
    \base_new_pp_reg[6]_3 ,
    \base_new_pp_reg[6]_4 ,
    \base_new_pp_reg[1]_0 ,
    \base_new_pp_reg[4]_3 ,
    \base_new_pp_reg[6]_5 ,
    \base_new_pp_reg[4]_4 ,
    \base_new_pp_reg[6]_6 ,
    \base_new_pp_reg[6]_7 ,
    \base_new_pp_reg[1]_1 ,
    \KR[3].key_host_reg[0][31] ,
    g_func,
    sbox_input,
    \CD[2].col_reg[1][0] ,
    \CD[2].col_reg[1][7] ,
    \CD[2].col_reg[1][15] ,
    \CD[2].col_reg[1][31] ,
    \CD[2].col_reg[1][1] ,
    \CD[2].col_reg[1][6] ,
    \CD[2].col_reg[1][14] ,
    \CD[2].col_reg[1][30] ,
    \CD[2].col_reg[1][2] ,
    \CD[2].col_reg[1][5] ,
    \CD[2].col_reg[1][13] ,
    \CD[2].col_reg[1][29] ,
    \CD[2].col_reg[1][3] ,
    \CD[2].col_reg[1][4] ,
    \CD[2].col_reg[1][12] ,
    \CD[2].col_reg[1][28] ,
    \CD[2].col_reg[1][11] ,
    \CD[2].col_reg[1][27] ,
    \CD[2].col_reg[1][10] ,
    \CD[2].col_reg[1][26] ,
    \CD[2].col_reg[1][9] ,
    \CD[2].col_reg[1][25] ,
    \CD[2].col_reg[1][8] ,
    \CD[2].col_reg[1][24] ,
    \CD[2].col_reg[1][23] ,
    \CD[2].col_reg[1][22] ,
    \CD[2].col_reg[1][21] ,
    \CD[2].col_reg[1][20] ,
    \CD[2].col_reg[1][19] ,
    \CD[2].col_reg[1][18] ,
    \CD[2].col_reg[1][17] ,
    \CD[2].col_reg[1][16] ,
    enable_i,
    Q,
    enc_dec_sbox,
    \sbox_pp2_reg[30] ,
    \sbox_pp2_reg[31] ,
    \sbox_pp2_reg[26] ,
    \sbox_pp2_reg[28] ,
    \sbox_pp2_reg[27] ,
    \sbox_pp2_reg[24] ,
    \sbox_pp2_reg[25] ,
    \sbox_pp2_reg[31]_0 ,
    \sbox_pp2_reg[18] ,
    \sbox_pp2_reg[22] ,
    \sbox_pp2_reg[19] ,
    \sbox_pp2_reg[20] ,
    \sbox_pp2_reg[17] ,
    \sbox_pp2_reg[23] ,
    \sbox_pp2_reg[10] ,
    \sbox_pp2_reg[14] ,
    \sbox_pp2_reg[11] ,
    \sbox_pp2_reg[12] ,
    \sbox_pp2_reg[9] ,
    \sbox_pp2_reg[15] ,
    \sbox_pp2_reg[2] ,
    \sbox_pp2_reg[6] ,
    \sbox_pp2_reg[3] ,
    \sbox_pp2_reg[4] ,
    \sbox_pp2_reg[1] ,
    \sbox_pp2_reg[7] ,
    key_en,
    \KR[3].key_reg[0][31] ,
    key_sel_mux,
    \KR[3].key_reg[0][31]_0 ,
    \sbox_pp2_reg[29] ,
    \sbox_pp2_reg[21] ,
    \sbox_pp2_reg[16] ,
    \sbox_pp2_reg[13] ,
    \sbox_pp2_reg[8] ,
    \sbox_pp2_reg[5] ,
    \sbox_pp2_reg[0] ,
    \base_new_pp_reg[4]_5 ,
    \base_new_pp_reg[2] ,
    \info_o[31]_INST_0_i_9 ,
    \info_o[28]_INST_0_i_7 ,
    \info_o[31]_INST_0_i_11 ,
    \info_o[31]_INST_0_i_11_0 ,
    \info_o[28]_INST_0_i_7_0 ,
    \CD[0].col[3][31]_i_14 ,
    \CD[0].col[3][7]_i_9 ,
    \CD[0].col[3][31]_i_14_0 ,
    \CD[0].col[3][7]_i_9_0 ,
    rc,
    isomorphism_return179_out,
    isomorphism_return114_out,
    \base_new_pp_reg[4]_6 ,
    \base_new_pp_reg[3] ,
    isomorphism_return179_out_12,
    isomorphism_return114_out_13,
    \base_new_pp_reg[4]_7 ,
    \base_new_pp_reg[3]_0 ,
    isomorphism_return179_out_14,
    isomorphism_return114_out_15,
    \base_new_pp_reg[4]_8 ,
    \base_new_pp_reg[3]_1 ,
    isomorphism_return179_out_16,
    isomorphism_return114_out_17,
    \base_new_pp_reg[4]_9 ,
    \base_new_pp_reg[3]_2 ,
    clk_i);
  output enable_i_0_sp_1;
  output \round_pp1_reg[0] ;
  output \round_pp1_reg[3] ;
  output \round_pp1_reg[3]_0 ;
  output \round_pp1_reg[0]_0 ;
  output \round_pp1_reg[3]_1 ;
  output [31:0]D;
  output \round_pp1_reg[0]_1 ;
  output \base_new_pp_reg[4] ;
  output [5:0]sbox_out_enc;
  output \base_new_pp_reg[6] ;
  output \base_new_pp_reg[4]_0 ;
  output \base_new_pp_reg[6]_0 ;
  output \base_new_pp_reg[6]_1 ;
  output \base_new_pp_reg[1] ;
  output \base_new_pp_reg[4]_1 ;
  output \base_new_pp_reg[6]_2 ;
  output \base_new_pp_reg[4]_2 ;
  output \base_new_pp_reg[6]_3 ;
  output \base_new_pp_reg[6]_4 ;
  output \base_new_pp_reg[1]_0 ;
  output \base_new_pp_reg[4]_3 ;
  output \base_new_pp_reg[6]_5 ;
  output \base_new_pp_reg[4]_4 ;
  output \base_new_pp_reg[6]_6 ;
  output \base_new_pp_reg[6]_7 ;
  output \base_new_pp_reg[1]_1 ;
  output [31:0]\KR[3].key_host_reg[0][31] ;
  output [1:0]g_func;
  output [31:0]sbox_input;
  output \CD[2].col_reg[1][0] ;
  output \CD[2].col_reg[1][7] ;
  output \CD[2].col_reg[1][15] ;
  output \CD[2].col_reg[1][31] ;
  output \CD[2].col_reg[1][1] ;
  output \CD[2].col_reg[1][6] ;
  output \CD[2].col_reg[1][14] ;
  output \CD[2].col_reg[1][30] ;
  output \CD[2].col_reg[1][2] ;
  output \CD[2].col_reg[1][5] ;
  output \CD[2].col_reg[1][13] ;
  output \CD[2].col_reg[1][29] ;
  output \CD[2].col_reg[1][3] ;
  output \CD[2].col_reg[1][4] ;
  output \CD[2].col_reg[1][12] ;
  output \CD[2].col_reg[1][28] ;
  output \CD[2].col_reg[1][11] ;
  output \CD[2].col_reg[1][27] ;
  output \CD[2].col_reg[1][10] ;
  output \CD[2].col_reg[1][26] ;
  output \CD[2].col_reg[1][9] ;
  output \CD[2].col_reg[1][25] ;
  output \CD[2].col_reg[1][8] ;
  output \CD[2].col_reg[1][24] ;
  output \CD[2].col_reg[1][23] ;
  output \CD[2].col_reg[1][22] ;
  output \CD[2].col_reg[1][21] ;
  output \CD[2].col_reg[1][20] ;
  output \CD[2].col_reg[1][19] ;
  output \CD[2].col_reg[1][18] ;
  output \CD[2].col_reg[1][17] ;
  output \CD[2].col_reg[1][16] ;
  input [31:0]enable_i;
  input [3:0]Q;
  input enc_dec_sbox;
  input \sbox_pp2_reg[30] ;
  input \sbox_pp2_reg[31] ;
  input \sbox_pp2_reg[26] ;
  input \sbox_pp2_reg[28] ;
  input \sbox_pp2_reg[27] ;
  input \sbox_pp2_reg[24] ;
  input \sbox_pp2_reg[25] ;
  input \sbox_pp2_reg[31]_0 ;
  input \sbox_pp2_reg[18] ;
  input \sbox_pp2_reg[22] ;
  input \sbox_pp2_reg[19] ;
  input \sbox_pp2_reg[20] ;
  input \sbox_pp2_reg[17] ;
  input \sbox_pp2_reg[23] ;
  input \sbox_pp2_reg[10] ;
  input \sbox_pp2_reg[14] ;
  input \sbox_pp2_reg[11] ;
  input \sbox_pp2_reg[12] ;
  input \sbox_pp2_reg[9] ;
  input \sbox_pp2_reg[15] ;
  input \sbox_pp2_reg[2] ;
  input \sbox_pp2_reg[6] ;
  input \sbox_pp2_reg[3] ;
  input \sbox_pp2_reg[4] ;
  input \sbox_pp2_reg[1] ;
  input \sbox_pp2_reg[7] ;
  input [0:0]key_en;
  input [31:0]\KR[3].key_reg[0][31] ;
  input key_sel_mux;
  input [31:0]\KR[3].key_reg[0][31]_0 ;
  input \sbox_pp2_reg[29] ;
  input \sbox_pp2_reg[21] ;
  input \sbox_pp2_reg[16] ;
  input \sbox_pp2_reg[13] ;
  input \sbox_pp2_reg[8] ;
  input \sbox_pp2_reg[5] ;
  input \sbox_pp2_reg[0] ;
  input \base_new_pp_reg[4]_5 ;
  input [31:0]\base_new_pp_reg[2] ;
  input [31:0]\info_o[31]_INST_0_i_9 ;
  input \info_o[28]_INST_0_i_7 ;
  input [31:0]\info_o[31]_INST_0_i_11 ;
  input [31:0]\info_o[31]_INST_0_i_11_0 ;
  input \info_o[28]_INST_0_i_7_0 ;
  input [31:0]\CD[0].col[3][31]_i_14 ;
  input \CD[0].col[3][7]_i_9 ;
  input [31:0]\CD[0].col[3][31]_i_14_0 ;
  input \CD[0].col[3][7]_i_9_0 ;
  input [1:0]rc;
  input isomorphism_return179_out;
  input isomorphism_return114_out;
  input \base_new_pp_reg[4]_6 ;
  input \base_new_pp_reg[3] ;
  input isomorphism_return179_out_12;
  input isomorphism_return114_out_13;
  input \base_new_pp_reg[4]_7 ;
  input \base_new_pp_reg[3]_0 ;
  input isomorphism_return179_out_14;
  input isomorphism_return114_out_15;
  input \base_new_pp_reg[4]_8 ;
  input \base_new_pp_reg[3]_1 ;
  input isomorphism_return179_out_16;
  input isomorphism_return114_out_17;
  input \base_new_pp_reg[4]_9 ;
  input \base_new_pp_reg[3]_2 ;
  input clk_i;

  wire [31:0]\CD[0].col[3][31]_i_14 ;
  wire [31:0]\CD[0].col[3][31]_i_14_0 ;
  wire \CD[0].col[3][7]_i_9 ;
  wire \CD[0].col[3][7]_i_9_0 ;
  wire \CD[2].col_reg[1][0] ;
  wire \CD[2].col_reg[1][10] ;
  wire \CD[2].col_reg[1][11] ;
  wire \CD[2].col_reg[1][12] ;
  wire \CD[2].col_reg[1][13] ;
  wire \CD[2].col_reg[1][14] ;
  wire \CD[2].col_reg[1][15] ;
  wire \CD[2].col_reg[1][16] ;
  wire \CD[2].col_reg[1][17] ;
  wire \CD[2].col_reg[1][18] ;
  wire \CD[2].col_reg[1][19] ;
  wire \CD[2].col_reg[1][1] ;
  wire \CD[2].col_reg[1][20] ;
  wire \CD[2].col_reg[1][21] ;
  wire \CD[2].col_reg[1][22] ;
  wire \CD[2].col_reg[1][23] ;
  wire \CD[2].col_reg[1][24] ;
  wire \CD[2].col_reg[1][25] ;
  wire \CD[2].col_reg[1][26] ;
  wire \CD[2].col_reg[1][27] ;
  wire \CD[2].col_reg[1][28] ;
  wire \CD[2].col_reg[1][29] ;
  wire \CD[2].col_reg[1][2] ;
  wire \CD[2].col_reg[1][30] ;
  wire \CD[2].col_reg[1][31] ;
  wire \CD[2].col_reg[1][3] ;
  wire \CD[2].col_reg[1][4] ;
  wire \CD[2].col_reg[1][5] ;
  wire \CD[2].col_reg[1][6] ;
  wire \CD[2].col_reg[1][7] ;
  wire \CD[2].col_reg[1][8] ;
  wire \CD[2].col_reg[1][9] ;
  wire [31:0]D;
  wire [31:0]\KR[3].key_host_reg[0][31] ;
  wire [31:0]\KR[3].key_reg[0][31] ;
  wire [31:0]\KR[3].key_reg[0][31]_0 ;
  wire [3:0]Q;
  wire \base_new_pp_reg[1] ;
  wire \base_new_pp_reg[1]_0 ;
  wire \base_new_pp_reg[1]_1 ;
  wire [31:0]\base_new_pp_reg[2] ;
  wire \base_new_pp_reg[3] ;
  wire \base_new_pp_reg[3]_0 ;
  wire \base_new_pp_reg[3]_1 ;
  wire \base_new_pp_reg[3]_2 ;
  wire \base_new_pp_reg[4] ;
  wire \base_new_pp_reg[4]_0 ;
  wire \base_new_pp_reg[4]_1 ;
  wire \base_new_pp_reg[4]_2 ;
  wire \base_new_pp_reg[4]_3 ;
  wire \base_new_pp_reg[4]_4 ;
  wire \base_new_pp_reg[4]_5 ;
  wire \base_new_pp_reg[4]_6 ;
  wire \base_new_pp_reg[4]_7 ;
  wire \base_new_pp_reg[4]_8 ;
  wire \base_new_pp_reg[4]_9 ;
  wire \base_new_pp_reg[6] ;
  wire \base_new_pp_reg[6]_0 ;
  wire \base_new_pp_reg[6]_1 ;
  wire \base_new_pp_reg[6]_2 ;
  wire \base_new_pp_reg[6]_3 ;
  wire \base_new_pp_reg[6]_4 ;
  wire \base_new_pp_reg[6]_5 ;
  wire \base_new_pp_reg[6]_6 ;
  wire \base_new_pp_reg[6]_7 ;
  wire clk_i;
  wire [31:0]enable_i;
  wire enable_i_0_sn_1;
  wire enc_dec_sbox;
  wire [1:0]g_func;
  wire \info_o[28]_INST_0_i_7 ;
  wire \info_o[28]_INST_0_i_7_0 ;
  wire [31:0]\info_o[31]_INST_0_i_11 ;
  wire [31:0]\info_o[31]_INST_0_i_11_0 ;
  wire [31:0]\info_o[31]_INST_0_i_9 ;
  wire isomorphism_return114_out;
  wire isomorphism_return114_out_13;
  wire isomorphism_return114_out_15;
  wire isomorphism_return114_out_17;
  wire isomorphism_return179_out;
  wire isomorphism_return179_out_12;
  wire isomorphism_return179_out_14;
  wire isomorphism_return179_out_16;
  wire [0:0]key_en;
  wire key_sel_mux;
  wire [1:0]rc;
  wire \round_pp1_reg[0] ;
  wire \round_pp1_reg[0]_0 ;
  wire \round_pp1_reg[0]_1 ;
  wire \round_pp1_reg[3] ;
  wire \round_pp1_reg[3]_0 ;
  wire \round_pp1_reg[3]_1 ;
  wire [31:0]sbox_input;
  wire [5:0]sbox_out_enc;
  wire \sbox_pp2_reg[0] ;
  wire \sbox_pp2_reg[10] ;
  wire \sbox_pp2_reg[11] ;
  wire \sbox_pp2_reg[12] ;
  wire \sbox_pp2_reg[13] ;
  wire \sbox_pp2_reg[14] ;
  wire \sbox_pp2_reg[15] ;
  wire \sbox_pp2_reg[16] ;
  wire \sbox_pp2_reg[17] ;
  wire \sbox_pp2_reg[18] ;
  wire \sbox_pp2_reg[19] ;
  wire \sbox_pp2_reg[1] ;
  wire \sbox_pp2_reg[20] ;
  wire \sbox_pp2_reg[21] ;
  wire \sbox_pp2_reg[22] ;
  wire \sbox_pp2_reg[23] ;
  wire \sbox_pp2_reg[24] ;
  wire \sbox_pp2_reg[25] ;
  wire \sbox_pp2_reg[26] ;
  wire \sbox_pp2_reg[27] ;
  wire \sbox_pp2_reg[28] ;
  wire \sbox_pp2_reg[29] ;
  wire \sbox_pp2_reg[2] ;
  wire \sbox_pp2_reg[30] ;
  wire \sbox_pp2_reg[31] ;
  wire \sbox_pp2_reg[31]_0 ;
  wire \sbox_pp2_reg[3] ;
  wire \sbox_pp2_reg[4] ;
  wire \sbox_pp2_reg[5] ;
  wire \sbox_pp2_reg[6] ;
  wire \sbox_pp2_reg[7] ;
  wire \sbox_pp2_reg[8] ;
  wire \sbox_pp2_reg[9] ;

  assign enable_i_0_sp_1 = enable_i_0_sn_1;
  switch_elements_sBox_8 \SBOX[0] 
       (.\CD[0].col[3][7]_i_9 (\CD[0].col[3][31]_i_14 [7:0]),
        .\CD[0].col[3][7]_i_9_0 (\CD[0].col[3][7]_i_9 ),
        .\CD[0].col[3][7]_i_9_1 (\CD[0].col[3][31]_i_14_0 [7:0]),
        .\CD[0].col[3][7]_i_9_2 (\CD[0].col[3][7]_i_9_0 ),
        .\CD[0].col_reg[3][0] (sbox_input[0]),
        .\CD[0].col_reg[3][1] (sbox_input[1]),
        .\CD[0].col_reg[3][2] (sbox_input[2]),
        .\CD[0].col_reg[3][3] (sbox_input[3]),
        .\CD[0].col_reg[3][4] (sbox_input[4]),
        .\CD[0].col_reg[3][5] (sbox_input[5]),
        .\CD[0].col_reg[3][6] (sbox_input[6]),
        .\CD[0].col_reg[3][7] (sbox_input[7]),
        .\CD[2].col_reg[1][0] (\CD[2].col_reg[1][0] ),
        .\CD[2].col_reg[1][1] (\CD[2].col_reg[1][1] ),
        .\CD[2].col_reg[1][2] (\CD[2].col_reg[1][2] ),
        .\CD[2].col_reg[1][3] (\CD[2].col_reg[1][3] ),
        .\CD[2].col_reg[1][4] (\CD[2].col_reg[1][4] ),
        .\CD[2].col_reg[1][5] (\CD[2].col_reg[1][5] ),
        .\CD[2].col_reg[1][6] (\CD[2].col_reg[1][6] ),
        .\CD[2].col_reg[1][7] (\CD[2].col_reg[1][7] ),
        .D(D[7:0]),
        .\KR[3].key_host_reg[0][7] (\KR[3].key_host_reg[0][31] [7:0]),
        .\KR[3].key_reg[0][7] (\KR[3].key_reg[0][31] [7:0]),
        .\KR[3].key_reg[0][7]_0 (\KR[3].key_reg[0][31]_0 [7:0]),
        .\base_new_pp_reg[1]_0 (\base_new_pp_reg[1]_1 ),
        .\base_new_pp_reg[2]_0 (\base_new_pp_reg[2] [7:0]),
        .\base_new_pp_reg[3]_0 (\base_new_pp_reg[3]_2 ),
        .\base_new_pp_reg[4]_0 (\base_new_pp_reg[4]_3 ),
        .\base_new_pp_reg[4]_1 (\base_new_pp_reg[4]_4 ),
        .\base_new_pp_reg[4]_2 (\base_new_pp_reg[4]_5 ),
        .\base_new_pp_reg[4]_3 (\base_new_pp_reg[4]_9 ),
        .\base_new_pp_reg[6]_0 (\base_new_pp_reg[6]_5 ),
        .\base_new_pp_reg[6]_1 (\base_new_pp_reg[6]_6 ),
        .\base_new_pp_reg[6]_2 (\base_new_pp_reg[6]_7 ),
        .clk_i(clk_i),
        .enable_i(enable_i[7:0]),
        .enc_dec_sbox(enc_dec_sbox),
        .\info_o[28]_INST_0_i_7_0 (\info_o[28]_INST_0_i_7 ),
        .\info_o[28]_INST_0_i_7_1 (\info_o[28]_INST_0_i_7_0 ),
        .\info_o[31]_INST_0_i_11_0 (\info_o[31]_INST_0_i_9 [7:0]),
        .\info_o[31]_INST_0_i_11_1 (\info_o[31]_INST_0_i_11 [31:24]),
        .\info_o[31]_INST_0_i_11_2 (\info_o[31]_INST_0_i_11_0 [31:24]),
        .isomorphism_return114_out_17(isomorphism_return114_out_17),
        .isomorphism_return179_out_16(isomorphism_return179_out_16),
        .key_en(key_en),
        .key_sel_mux(key_sel_mux),
        .sbox_out_enc(sbox_out_enc[1:0]),
        .\sbox_pp2_reg[0] (\sbox_pp2_reg[0] ),
        .\sbox_pp2_reg[1] (\sbox_pp2_reg[1] ),
        .\sbox_pp2_reg[2] (\sbox_pp2_reg[2] ),
        .\sbox_pp2_reg[3] (\sbox_pp2_reg[3] ),
        .\sbox_pp2_reg[4] (\sbox_pp2_reg[4] ),
        .\sbox_pp2_reg[5] (\sbox_pp2_reg[5] ),
        .\sbox_pp2_reg[6] (\sbox_pp2_reg[6] ),
        .\sbox_pp2_reg[7] (\sbox_pp2_reg[31] ),
        .\sbox_pp2_reg[7]_0 (\sbox_pp2_reg[7] ));
  switch_elements_sBox_8_1 \SBOX[1] 
       (.\CD[0].col[3][15]_i_7 (\CD[0].col[3][31]_i_14 [15:8]),
        .\CD[0].col[3][15]_i_7_0 (\CD[0].col[3][7]_i_9 ),
        .\CD[0].col[3][15]_i_7_1 (\CD[0].col[3][31]_i_14_0 [15:8]),
        .\CD[0].col[3][15]_i_7_2 (\CD[0].col[3][7]_i_9_0 ),
        .\CD[0].col_reg[3][10] (sbox_input[10]),
        .\CD[0].col_reg[3][11] (sbox_input[11]),
        .\CD[0].col_reg[3][12] (sbox_input[12]),
        .\CD[0].col_reg[3][13] (sbox_input[13]),
        .\CD[0].col_reg[3][14] (sbox_input[14]),
        .\CD[0].col_reg[3][15] (sbox_input[15]),
        .\CD[0].col_reg[3][8] (sbox_input[8]),
        .\CD[0].col_reg[3][9] (sbox_input[9]),
        .\CD[2].col_reg[1][10] (\CD[2].col_reg[1][10] ),
        .\CD[2].col_reg[1][11] (\CD[2].col_reg[1][11] ),
        .\CD[2].col_reg[1][12] (\CD[2].col_reg[1][12] ),
        .\CD[2].col_reg[1][13] (\CD[2].col_reg[1][13] ),
        .\CD[2].col_reg[1][14] (\CD[2].col_reg[1][14] ),
        .\CD[2].col_reg[1][15] (\CD[2].col_reg[1][15] ),
        .\CD[2].col_reg[1][8] (\CD[2].col_reg[1][8] ),
        .\CD[2].col_reg[1][9] (\CD[2].col_reg[1][9] ),
        .D(D[15:8]),
        .\KR[3].key_host_reg[0][15] (\KR[3].key_host_reg[0][31] [15:8]),
        .\KR[3].key_reg[0][15] (\KR[3].key_reg[0][31] [15:8]),
        .\KR[3].key_reg[0][15]_0 (\KR[3].key_reg[0][31]_0 [15:8]),
        .\base_new_pp[4]_i_2__1_0 (\info_o[28]_INST_0_i_7 ),
        .\base_new_pp[4]_i_2__1_1 (\info_o[28]_INST_0_i_7_0 ),
        .\base_new_pp_reg[1]_0 (\base_new_pp_reg[1]_0 ),
        .\base_new_pp_reg[2]_0 (\base_new_pp_reg[2] [15:8]),
        .\base_new_pp_reg[3]_0 (\base_new_pp_reg[3]_1 ),
        .\base_new_pp_reg[4]_0 (\base_new_pp_reg[4]_1 ),
        .\base_new_pp_reg[4]_1 (\base_new_pp_reg[4]_2 ),
        .\base_new_pp_reg[4]_2 (\base_new_pp_reg[4]_5 ),
        .\base_new_pp_reg[4]_3 (\base_new_pp_reg[4]_8 ),
        .\base_new_pp_reg[6]_0 (\base_new_pp_reg[6]_2 ),
        .\base_new_pp_reg[6]_1 (\base_new_pp_reg[6]_3 ),
        .\base_new_pp_reg[6]_2 (\base_new_pp_reg[6]_4 ),
        .clk_i(clk_i),
        .enable_i(enable_i[15:8]),
        .enc_dec_sbox(enc_dec_sbox),
        .\info_o[31]_INST_0_i_8_0 (\info_o[31]_INST_0_i_9 [15:8]),
        .\info_o[31]_INST_0_i_8_1 (\info_o[31]_INST_0_i_11 [7:0]),
        .\info_o[31]_INST_0_i_8_2 (\info_o[31]_INST_0_i_11_0 [7:0]),
        .isomorphism_return114_out_15(isomorphism_return114_out_15),
        .isomorphism_return179_out_14(isomorphism_return179_out_14),
        .key_en(key_en),
        .key_sel_mux(key_sel_mux),
        .sbox_out_enc(sbox_out_enc[3:2]),
        .\sbox_pp2_reg[10] (\sbox_pp2_reg[10] ),
        .\sbox_pp2_reg[11] (\sbox_pp2_reg[11] ),
        .\sbox_pp2_reg[12] (\sbox_pp2_reg[12] ),
        .\sbox_pp2_reg[13] (\sbox_pp2_reg[13] ),
        .\sbox_pp2_reg[14] (\sbox_pp2_reg[14] ),
        .\sbox_pp2_reg[15] (\sbox_pp2_reg[31] ),
        .\sbox_pp2_reg[15]_0 (\sbox_pp2_reg[15] ),
        .\sbox_pp2_reg[8] (\sbox_pp2_reg[8] ),
        .\sbox_pp2_reg[9] (\sbox_pp2_reg[9] ));
  switch_elements_sBox_8_2 \SBOX[2] 
       (.\CD[0].col_reg[3][16] (sbox_input[16]),
        .\CD[0].col_reg[3][17] (sbox_input[17]),
        .\CD[0].col_reg[3][18] (sbox_input[18]),
        .\CD[0].col_reg[3][19] (sbox_input[19]),
        .\CD[0].col_reg[3][20] (sbox_input[20]),
        .\CD[0].col_reg[3][21] (sbox_input[21]),
        .\CD[0].col_reg[3][22] (sbox_input[22]),
        .\CD[0].col_reg[3][23] (sbox_input[23]),
        .\CD[1].col[2][23]_i_3 (\CD[0].col[3][31]_i_14 [23:16]),
        .\CD[1].col[2][23]_i_3_0 (\CD[0].col[3][7]_i_9 ),
        .\CD[1].col[2][23]_i_3_1 (\CD[0].col[3][31]_i_14_0 [23:16]),
        .\CD[1].col[2][23]_i_3_2 (\CD[0].col[3][7]_i_9_0 ),
        .\CD[2].col_reg[1][16] (\CD[2].col_reg[1][16] ),
        .\CD[2].col_reg[1][17] (\CD[2].col_reg[1][17] ),
        .\CD[2].col_reg[1][18] (\CD[2].col_reg[1][18] ),
        .\CD[2].col_reg[1][19] (\CD[2].col_reg[1][19] ),
        .\CD[2].col_reg[1][20] (\CD[2].col_reg[1][20] ),
        .\CD[2].col_reg[1][21] (\CD[2].col_reg[1][21] ),
        .\CD[2].col_reg[1][22] (\CD[2].col_reg[1][22] ),
        .\CD[2].col_reg[1][23] (\CD[2].col_reg[1][23] ),
        .D(D[23:16]),
        .\KR[3].key_host_reg[0][23] (\KR[3].key_host_reg[0][31] [23:16]),
        .\KR[3].key_reg[0][23] (\KR[3].key_reg[0][31] [23:16]),
        .\KR[3].key_reg[0][23]_0 (\KR[3].key_reg[0][31]_0 [23:16]),
        .\base_new_pp[4]_i_2__0_0 (\info_o[28]_INST_0_i_7 ),
        .\base_new_pp[4]_i_2__0_1 (\info_o[28]_INST_0_i_7_0 ),
        .\base_new_pp_reg[1]_0 (\base_new_pp_reg[1] ),
        .\base_new_pp_reg[2]_0 (\base_new_pp_reg[2] [23:16]),
        .\base_new_pp_reg[3]_0 (\base_new_pp_reg[3]_0 ),
        .\base_new_pp_reg[4]_0 (\base_new_pp_reg[4] ),
        .\base_new_pp_reg[4]_1 (\base_new_pp_reg[4]_0 ),
        .\base_new_pp_reg[4]_2 (\base_new_pp_reg[4]_5 ),
        .\base_new_pp_reg[4]_3 (\base_new_pp_reg[4]_7 ),
        .\base_new_pp_reg[6]_0 (\base_new_pp_reg[6] ),
        .\base_new_pp_reg[6]_1 (\base_new_pp_reg[6]_0 ),
        .\base_new_pp_reg[6]_2 (\base_new_pp_reg[6]_1 ),
        .clk_i(clk_i),
        .enable_i({enable_i[23:16],enable_i[6],enable_i[4:0]}),
        .enable_i_0_sp_1(enable_i_0_sn_1),
        .enc_dec_sbox(enc_dec_sbox),
        .\info_o[23]_INST_0_i_4_0 (\info_o[31]_INST_0_i_9 [23:16]),
        .\info_o[23]_INST_0_i_4_1 (\info_o[31]_INST_0_i_11 [15:8]),
        .\info_o[23]_INST_0_i_4_2 (\info_o[31]_INST_0_i_11_0 [15:8]),
        .isomorphism_return114_out_13(isomorphism_return114_out_13),
        .isomorphism_return179_out_12(isomorphism_return179_out_12),
        .key_en(key_en),
        .key_sel_mux(key_sel_mux),
        .sbox_out_enc(sbox_out_enc[5:4]),
        .\sbox_pp2_reg[16] (\sbox_pp2_reg[16] ),
        .\sbox_pp2_reg[17] (\sbox_pp2_reg[17] ),
        .\sbox_pp2_reg[18] (\sbox_pp2_reg[18] ),
        .\sbox_pp2_reg[19] (\sbox_pp2_reg[19] ),
        .\sbox_pp2_reg[20] (\sbox_pp2_reg[20] ),
        .\sbox_pp2_reg[21] (\sbox_pp2_reg[21] ),
        .\sbox_pp2_reg[22] (\sbox_pp2_reg[22] ),
        .\sbox_pp2_reg[23] (\sbox_pp2_reg[31] ),
        .\sbox_pp2_reg[23]_0 (\sbox_pp2_reg[23] ));
  switch_elements_sBox_8_3 \SBOX[3] 
       (.\CD[0].col[3][31]_i_14 (\CD[0].col[3][31]_i_14 [31:24]),
        .\CD[0].col[3][31]_i_14_0 (\CD[0].col[3][7]_i_9 ),
        .\CD[0].col[3][31]_i_14_1 (\CD[0].col[3][31]_i_14_0 [31:24]),
        .\CD[0].col[3][31]_i_14_2 (\CD[0].col[3][7]_i_9_0 ),
        .\CD[0].col_reg[3][24] (sbox_input[24]),
        .\CD[0].col_reg[3][25] (sbox_input[25]),
        .\CD[0].col_reg[3][26] (sbox_input[26]),
        .\CD[0].col_reg[3][27] (sbox_input[27]),
        .\CD[0].col_reg[3][28] (sbox_input[28]),
        .\CD[0].col_reg[3][29] (sbox_input[29]),
        .\CD[0].col_reg[3][30] (sbox_input[30]),
        .\CD[0].col_reg[3][31] (sbox_input[31]),
        .\CD[2].col_reg[1][24] (\CD[2].col_reg[1][24] ),
        .\CD[2].col_reg[1][25] (\CD[2].col_reg[1][25] ),
        .\CD[2].col_reg[1][26] (\CD[2].col_reg[1][26] ),
        .\CD[2].col_reg[1][27] (\CD[2].col_reg[1][27] ),
        .\CD[2].col_reg[1][28] (\CD[2].col_reg[1][28] ),
        .\CD[2].col_reg[1][29] (\CD[2].col_reg[1][29] ),
        .\CD[2].col_reg[1][30] (\CD[2].col_reg[1][30] ),
        .\CD[2].col_reg[1][31] (\CD[2].col_reg[1][31] ),
        .D(D[31:24]),
        .\KR[3].key_host_reg[0][31] (\KR[3].key_host_reg[0][31] [31:24]),
        .\KR[3].key_reg[0][31] (\KR[3].key_reg[0][31] [31:24]),
        .\KR[3].key_reg[0][31]_0 (\KR[3].key_reg[0][31]_0 [31:24]),
        .Q(Q),
        .\base_new_pp[4]_i_2_0 (\info_o[28]_INST_0_i_7 ),
        .\base_new_pp[4]_i_2_1 (\info_o[28]_INST_0_i_7_0 ),
        .\base_new_pp_reg[2]_0 (\base_new_pp_reg[2] [31:24]),
        .\base_new_pp_reg[3]_0 (\base_new_pp_reg[3] ),
        .\base_new_pp_reg[4]_0 (\base_new_pp_reg[4]_5 ),
        .\base_new_pp_reg[4]_1 (\base_new_pp_reg[4]_6 ),
        .clk_i(clk_i),
        .enable_i(enable_i[31:24]),
        .enc_dec_sbox(enc_dec_sbox),
        .g_func(g_func),
        .\info_o[31]_INST_0_i_9_0 (\info_o[31]_INST_0_i_9 [31:24]),
        .\info_o[31]_INST_0_i_9_1 (\info_o[31]_INST_0_i_11 [23:16]),
        .\info_o[31]_INST_0_i_9_2 (\info_o[31]_INST_0_i_11_0 [23:16]),
        .isomorphism_return114_out(isomorphism_return114_out),
        .isomorphism_return179_out(isomorphism_return179_out),
        .key_en(key_en),
        .key_sel_mux(key_sel_mux),
        .rc(rc),
        .\round_pp1_reg[0] (\round_pp1_reg[0] ),
        .\round_pp1_reg[0]_0 (\round_pp1_reg[0]_0 ),
        .\round_pp1_reg[0]_1 (\round_pp1_reg[0]_1 ),
        .\round_pp1_reg[3] (\round_pp1_reg[3] ),
        .\round_pp1_reg[3]_0 (\round_pp1_reg[3]_0 ),
        .\round_pp1_reg[3]_1 (\round_pp1_reg[3]_1 ),
        .\sbox_pp2_reg[24] (\sbox_pp2_reg[24] ),
        .\sbox_pp2_reg[25] (\sbox_pp2_reg[25] ),
        .\sbox_pp2_reg[26] (\sbox_pp2_reg[26] ),
        .\sbox_pp2_reg[27] (\sbox_pp2_reg[27] ),
        .\sbox_pp2_reg[28] (\sbox_pp2_reg[28] ),
        .\sbox_pp2_reg[29] (\sbox_pp2_reg[29] ),
        .\sbox_pp2_reg[30] (\sbox_pp2_reg[30] ),
        .\sbox_pp2_reg[31] (\sbox_pp2_reg[31] ),
        .\sbox_pp2_reg[31]_0 (\sbox_pp2_reg[31]_0 ));
endmodule

(* ORIG_REF_NAME = "sBox_8" *) 
module switch_elements_sBox_8
   (D,
    \base_new_pp_reg[4]_0 ,
    sbox_out_enc,
    \base_new_pp_reg[6]_0 ,
    \base_new_pp_reg[4]_1 ,
    \base_new_pp_reg[6]_1 ,
    \base_new_pp_reg[6]_2 ,
    \base_new_pp_reg[1]_0 ,
    \KR[3].key_host_reg[0][7] ,
    \CD[0].col_reg[3][0] ,
    \CD[2].col_reg[1][0] ,
    \CD[0].col_reg[3][7] ,
    \CD[2].col_reg[1][7] ,
    \CD[0].col_reg[3][1] ,
    \CD[2].col_reg[1][1] ,
    \CD[0].col_reg[3][6] ,
    \CD[2].col_reg[1][6] ,
    \CD[0].col_reg[3][2] ,
    \CD[2].col_reg[1][2] ,
    \CD[0].col_reg[3][5] ,
    \CD[2].col_reg[1][5] ,
    \CD[0].col_reg[3][3] ,
    \CD[2].col_reg[1][3] ,
    \CD[0].col_reg[3][4] ,
    \CD[2].col_reg[1][4] ,
    \sbox_pp2_reg[2] ,
    \sbox_pp2_reg[7] ,
    \sbox_pp2_reg[6] ,
    \sbox_pp2_reg[3] ,
    \sbox_pp2_reg[4] ,
    \sbox_pp2_reg[1] ,
    \sbox_pp2_reg[7]_0 ,
    key_en,
    \KR[3].key_reg[0][7] ,
    enable_i,
    key_sel_mux,
    \KR[3].key_reg[0][7]_0 ,
    \sbox_pp2_reg[5] ,
    \sbox_pp2_reg[0] ,
    \base_new_pp_reg[4]_2 ,
    \base_new_pp_reg[2]_0 ,
    \info_o[31]_INST_0_i_11_0 ,
    \info_o[28]_INST_0_i_7_0 ,
    enc_dec_sbox,
    \info_o[31]_INST_0_i_11_1 ,
    \info_o[31]_INST_0_i_11_2 ,
    \info_o[28]_INST_0_i_7_1 ,
    \CD[0].col[3][7]_i_9 ,
    \CD[0].col[3][7]_i_9_0 ,
    \CD[0].col[3][7]_i_9_1 ,
    \CD[0].col[3][7]_i_9_2 ,
    isomorphism_return179_out_16,
    isomorphism_return114_out_17,
    \base_new_pp_reg[4]_3 ,
    \base_new_pp_reg[3]_0 ,
    clk_i);
  output [7:0]D;
  output \base_new_pp_reg[4]_0 ;
  output [1:0]sbox_out_enc;
  output \base_new_pp_reg[6]_0 ;
  output \base_new_pp_reg[4]_1 ;
  output \base_new_pp_reg[6]_1 ;
  output \base_new_pp_reg[6]_2 ;
  output \base_new_pp_reg[1]_0 ;
  output [7:0]\KR[3].key_host_reg[0][7] ;
  output \CD[0].col_reg[3][0] ;
  output \CD[2].col_reg[1][0] ;
  output \CD[0].col_reg[3][7] ;
  output \CD[2].col_reg[1][7] ;
  output \CD[0].col_reg[3][1] ;
  output \CD[2].col_reg[1][1] ;
  output \CD[0].col_reg[3][6] ;
  output \CD[2].col_reg[1][6] ;
  output \CD[0].col_reg[3][2] ;
  output \CD[2].col_reg[1][2] ;
  output \CD[0].col_reg[3][5] ;
  output \CD[2].col_reg[1][5] ;
  output \CD[0].col_reg[3][3] ;
  output \CD[2].col_reg[1][3] ;
  output \CD[0].col_reg[3][4] ;
  output \CD[2].col_reg[1][4] ;
  input \sbox_pp2_reg[2] ;
  input \sbox_pp2_reg[7] ;
  input \sbox_pp2_reg[6] ;
  input \sbox_pp2_reg[3] ;
  input \sbox_pp2_reg[4] ;
  input \sbox_pp2_reg[1] ;
  input \sbox_pp2_reg[7]_0 ;
  input [0:0]key_en;
  input [7:0]\KR[3].key_reg[0][7] ;
  input [7:0]enable_i;
  input key_sel_mux;
  input [7:0]\KR[3].key_reg[0][7]_0 ;
  input \sbox_pp2_reg[5] ;
  input \sbox_pp2_reg[0] ;
  input \base_new_pp_reg[4]_2 ;
  input [7:0]\base_new_pp_reg[2]_0 ;
  input [7:0]\info_o[31]_INST_0_i_11_0 ;
  input \info_o[28]_INST_0_i_7_0 ;
  input enc_dec_sbox;
  input [7:0]\info_o[31]_INST_0_i_11_1 ;
  input [7:0]\info_o[31]_INST_0_i_11_2 ;
  input \info_o[28]_INST_0_i_7_1 ;
  input [7:0]\CD[0].col[3][7]_i_9 ;
  input \CD[0].col[3][7]_i_9_0 ;
  input [7:0]\CD[0].col[3][7]_i_9_1 ;
  input \CD[0].col[3][7]_i_9_2 ;
  input isomorphism_return179_out_16;
  input isomorphism_return114_out_17;
  input \base_new_pp_reg[4]_3 ;
  input \base_new_pp_reg[3]_0 ;
  input clk_i;

  wire [7:0]\CD[0].col[3][7]_i_9 ;
  wire \CD[0].col[3][7]_i_9_0 ;
  wire [7:0]\CD[0].col[3][7]_i_9_1 ;
  wire \CD[0].col[3][7]_i_9_2 ;
  wire \CD[0].col_reg[3][0] ;
  wire \CD[0].col_reg[3][1] ;
  wire \CD[0].col_reg[3][2] ;
  wire \CD[0].col_reg[3][3] ;
  wire \CD[0].col_reg[3][4] ;
  wire \CD[0].col_reg[3][5] ;
  wire \CD[0].col_reg[3][6] ;
  wire \CD[0].col_reg[3][7] ;
  wire \CD[2].col_reg[1][0] ;
  wire \CD[2].col_reg[1][1] ;
  wire \CD[2].col_reg[1][2] ;
  wire \CD[2].col_reg[1][3] ;
  wire \CD[2].col_reg[1][4] ;
  wire \CD[2].col_reg[1][5] ;
  wire \CD[2].col_reg[1][6] ;
  wire \CD[2].col_reg[1][7] ;
  wire [7:0]D;
  wire [7:0]\KR[3].key_host_reg[0][7] ;
  wire [7:0]\KR[3].key_reg[0][7] ;
  wire [7:0]\KR[3].key_reg[0][7]_0 ;
  wire \base_new_pp[0]_i_1__2_n_0 ;
  wire \base_new_pp[4]_i_1__2_n_0 ;
  wire \base_new_pp_reg[1]_0 ;
  wire [7:0]\base_new_pp_reg[2]_0 ;
  wire \base_new_pp_reg[3]_0 ;
  wire \base_new_pp_reg[4]_0 ;
  wire \base_new_pp_reg[4]_1 ;
  wire \base_new_pp_reg[4]_2 ;
  wire \base_new_pp_reg[4]_3 ;
  wire \base_new_pp_reg[6]_0 ;
  wire \base_new_pp_reg[6]_1 ;
  wire \base_new_pp_reg[6]_2 ;
  wire \base_new_pp_reg_n_0_[0] ;
  wire \base_new_pp_reg_n_0_[1] ;
  wire \base_new_pp_reg_n_0_[4] ;
  wire \base_new_pp_reg_n_0_[5] ;
  wire clk_i;
  wire [7:0]enable_i;
  wire enc_dec_sbox;
  wire [3:0]gf_inv_8_stage1_return;
  wire gf_inv_8_stage1_return1__0;
  wire gf_inv_8_stage1_return2__0;
  wire gf_inv_8_stage1_return349_in;
  wire gf_inv_8_stage1_return540_out;
  wire gf_inv_8_stage1_return542_out;
  wire gf_inv_8_stage1_return546_out;
  wire gf_inv_8_stage1_return547_out;
  wire [1:0]gf_inv_8_stage2_return013_out;
  wire [1:1]gf_inv_8_stage2_return0__3;
  wire [1:0]gf_muls_20_return__1;
  wire [1:0]gf_muls_scl_20_return;
  wire [1:0]gf_muls_scl_2_return;
  wire [1:0]in111_out;
  wire [1:0]in1__0;
  wire [1:0]in2;
  wire [1:0]in21_in;
  wire \info_o[28]_INST_0_i_13_n_0 ;
  wire \info_o[28]_INST_0_i_15_n_0 ;
  wire \info_o[28]_INST_0_i_7_0 ;
  wire \info_o[28]_INST_0_i_7_1 ;
  wire \info_o[29]_INST_0_i_13_n_0 ;
  wire \info_o[29]_INST_0_i_15_n_0 ;
  wire \info_o[30]_INST_0_i_13_n_0 ;
  wire \info_o[30]_INST_0_i_15_n_0 ;
  wire [7:0]\info_o[31]_INST_0_i_11_0 ;
  wire [7:0]\info_o[31]_INST_0_i_11_1 ;
  wire [7:0]\info_o[31]_INST_0_i_11_2 ;
  wire \info_o[31]_INST_0_i_22_n_0 ;
  wire \info_o[31]_INST_0_i_24_n_0 ;
  wire isomorphism_return076_out;
  wire isomorphism_return114_out_17;
  wire isomorphism_return179_out_16;
  wire isomorphism_return1__0;
  wire isomorphism_return277_out;
  wire [0:0]key_en;
  wire key_sel_mux;
  wire \out_gf_pp[1]_i_3__2_n_0 ;
  wire \out_gf_pp[1]_i_4__2_n_0 ;
  wire \out_gf_pp[2]_i_2__2_n_0 ;
  wire \out_gf_pp[2]_i_6__2_n_0 ;
  wire \out_gf_pp[2]_i_7__2_n_0 ;
  wire \out_gf_pp[3]_i_2__2_n_0 ;
  wire \out_gf_pp[3]_i_5__2_n_0 ;
  wire \out_gf_pp[3]_i_6__2_n_0 ;
  wire \out_gf_pp[3]_i_7__2_n_0 ;
  wire \out_gf_pp_reg_n_0_[0] ;
  wire \out_gf_pp_reg_n_0_[1] ;
  wire \out_gf_pp_reg_n_0_[2] ;
  wire \out_gf_pp_reg_n_0_[3] ;
  wire p_0_in;
  wire p_0_in2_in;
  wire p_0_in9_in;
  wire p_1_in;
  wire p_1_in10_in;
  wire p_1_in17_in;
  wire p_1_in18_in;
  wire p_1_in7_in;
  wire p_72_in;
  wire [0:0]sbox_out_dec;
  wire [1:0]sbox_out_enc;
  wire \sbox_pp2_reg[0] ;
  wire \sbox_pp2_reg[1] ;
  wire \sbox_pp2_reg[2] ;
  wire \sbox_pp2_reg[3] ;
  wire \sbox_pp2_reg[4] ;
  wire \sbox_pp2_reg[5] ;
  wire \sbox_pp2_reg[6] ;
  wire \sbox_pp2_reg[7] ;
  wire \sbox_pp2_reg[7]_0 ;

  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \KR[2].key[1][0]_i_3 
       (.I0(p_0_in2_in),
        .I1(gf_inv_8_stage2_return013_out[0]),
        .I2(gf_inv_8_stage2_return0__3),
        .O(\base_new_pp_reg[1]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \KR[2].key[1][1]_i_3 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(p_1_in),
        .I2(p_0_in2_in),
        .O(\base_new_pp_reg[4]_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \KR[2].key[1][2]_i_3 
       (.I0(\base_new_pp_reg[6]_2 ),
        .I1(sbox_out_dec),
        .I2(\base_new_pp_reg[4]_1 ),
        .O(sbox_out_enc[0]));
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \KR[2].key[1][3]_i_3 
       (.I0(p_0_in2_in),
        .I1(gf_inv_8_stage2_return013_out[0]),
        .I2(\base_new_pp_reg[6]_0 ),
        .O(sbox_out_enc[1]));
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \KR[2].key[1][4]_i_3 
       (.I0(\base_new_pp_reg[6]_1 ),
        .I1(p_1_in),
        .O(\base_new_pp_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h96A59955695A66AA)) 
    \KR[2].key[1][5]_i_3 
       (.I0(gf_muls_scl_20_return[0]),
        .I1(\base_new_pp_reg_n_0_[4] ),
        .I2(gf_muls_20_return__1[0]),
        .I3(gf_muls_20_return__1[1]),
        .I4(\base_new_pp_reg_n_0_[5] ),
        .I5(gf_inv_8_stage2_return013_out[0]),
        .O(\base_new_pp_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h609F9F6060606060)) 
    \KR[2].key[1][5]_i_4 
       (.I0(\base_new_pp_reg_n_0_[5] ),
        .I1(in2[1]),
        .I2(in111_out[1]),
        .I3(\base_new_pp_reg_n_0_[4] ),
        .I4(in2[0]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_20_return[0]));
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT4 #(
    .INIT(16'hBE22)) 
    \KR[2].key[1][5]_i_5 
       (.I0(\out_gf_pp_reg_n_0_[2] ),
        .I1(\out_gf_pp_reg_n_0_[0] ),
        .I2(\out_gf_pp_reg_n_0_[1] ),
        .I3(\out_gf_pp_reg_n_0_[3] ),
        .O(gf_muls_20_return__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT4 #(
    .INIT(16'hDD82)) 
    \KR[2].key[1][5]_i_6 
       (.I0(\out_gf_pp_reg_n_0_[3] ),
        .I1(\out_gf_pp_reg_n_0_[1] ),
        .I2(\out_gf_pp_reg_n_0_[0] ),
        .I3(\out_gf_pp_reg_n_0_[2] ),
        .O(gf_muls_20_return__1[1]));
  LUT6 #(
    .INIT(64'hE4281BD71BD7E428)) 
    \KR[2].key[1][6]_i_3 
       (.I0(in2[0]),
        .I1(in1__0[0]),
        .I2(in1__0[1]),
        .I3(in2[1]),
        .I4(gf_muls_scl_20_return[1]),
        .I5(gf_inv_8_stage2_return013_out[1]),
        .O(\base_new_pp_reg[6]_1 ));
  LUT6 #(
    .INIT(64'h1BD7E428E4281BD7)) 
    \KR[2].key[1][7]_i_3 
       (.I0(in2[0]),
        .I1(in1__0[0]),
        .I2(in1__0[1]),
        .I3(in2[1]),
        .I4(gf_muls_scl_20_return[1]),
        .I5(p_1_in),
        .O(\base_new_pp_reg[6]_2 ));
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT4 #(
    .INIT(16'hB2E2)) 
    \KR[2].key[1][7]_i_4 
       (.I0(\out_gf_pp_reg_n_0_[0] ),
        .I1(\out_gf_pp_reg_n_0_[2] ),
        .I2(\out_gf_pp_reg_n_0_[1] ),
        .I3(\out_gf_pp_reg_n_0_[3] ),
        .O(in1__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT4 #(
    .INIT(16'hE4C6)) 
    \KR[2].key[1][7]_i_5 
       (.I0(\out_gf_pp_reg_n_0_[1] ),
        .I1(\out_gf_pp_reg_n_0_[0] ),
        .I2(\out_gf_pp_reg_n_0_[3] ),
        .I3(\out_gf_pp_reg_n_0_[2] ),
        .O(in1__0[1]));
  LUT6 #(
    .INIT(64'h0FF0666669960000)) 
    \KR[2].key[1][7]_i_6 
       (.I0(in2[1]),
        .I1(\base_new_pp_reg_n_0_[5] ),
        .I2(in2[0]),
        .I3(\base_new_pp_reg_n_0_[4] ),
        .I4(in111_out[1]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_20_return[1]));
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT4 #(
    .INIT(16'h23D6)) 
    \KR[2].key[1][7]_i_7 
       (.I0(\out_gf_pp_reg_n_0_[2] ),
        .I1(\out_gf_pp_reg_n_0_[3] ),
        .I2(\out_gf_pp_reg_n_0_[0] ),
        .I3(\out_gf_pp_reg_n_0_[1] ),
        .O(in111_out[1]));
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT4 #(
    .INIT(16'h6DB0)) 
    \KR[2].key[1][7]_i_8 
       (.I0(\out_gf_pp_reg_n_0_[3] ),
        .I1(\out_gf_pp_reg_n_0_[1] ),
        .I2(\out_gf_pp_reg_n_0_[2] ),
        .I3(\out_gf_pp_reg_n_0_[0] ),
        .O(in111_out[0]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][0]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][7] [0]),
        .I2(enable_i[0]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[1]_0 ),
        .I5(\KR[3].key_reg[0][7]_0 [0]),
        .O(\KR[3].key_host_reg[0][7] [0]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][1]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][7] [1]),
        .I2(enable_i[1]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[4]_0 ),
        .I5(\KR[3].key_reg[0][7]_0 [1]),
        .O(\KR[3].key_host_reg[0][7] [1]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][2]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][7] [2]),
        .I2(enable_i[2]),
        .I3(key_sel_mux),
        .I4(sbox_out_enc[0]),
        .I5(\KR[3].key_reg[0][7]_0 [2]),
        .O(\KR[3].key_host_reg[0][7] [2]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][3]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][7] [3]),
        .I2(enable_i[3]),
        .I3(key_sel_mux),
        .I4(sbox_out_enc[1]),
        .I5(\KR[3].key_reg[0][7]_0 [3]),
        .O(\KR[3].key_host_reg[0][7] [3]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][4]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][7] [4]),
        .I2(enable_i[4]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[6]_0 ),
        .I5(\KR[3].key_reg[0][7]_0 [4]),
        .O(\KR[3].key_host_reg[0][7] [4]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][5]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][7] [5]),
        .I2(enable_i[5]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[4]_1 ),
        .I5(\KR[3].key_reg[0][7]_0 [5]),
        .O(\KR[3].key_host_reg[0][7] [5]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][6]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][7] [6]),
        .I2(enable_i[6]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[6]_1 ),
        .I5(\KR[3].key_reg[0][7]_0 [6]),
        .O(\KR[3].key_host_reg[0][7] [6]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][7]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][7] [7]),
        .I2(enable_i[7]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[6]_2 ),
        .I5(\KR[3].key_reg[0][7]_0 [7]),
        .O(\KR[3].key_host_reg[0][7] [7]));
  LUT5 #(
    .INIT(32'h66F0660F)) 
    \base_new_pp[0]_i_1__2 
       (.I0(\CD[0].col_reg[3][2] ),
        .I1(isomorphism_return1__0),
        .I2(\CD[0].col_reg[3][1] ),
        .I3(enc_dec_sbox),
        .I4(isomorphism_return076_out),
        .O(\base_new_pp[0]_i_1__2_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \base_new_pp[0]_i_2__2 
       (.I0(\CD[0].col_reg[3][1] ),
        .I1(\CD[0].col_reg[3][0] ),
        .I2(\CD[0].col_reg[3][6] ),
        .I3(\CD[0].col_reg[3][3] ),
        .O(isomorphism_return1__0));
  LUT4 #(
    .INIT(16'h9669)) 
    \base_new_pp[0]_i_3__2 
       (.I0(\CD[0].col_reg[3][5] ),
        .I1(\CD[0].col_reg[3][0] ),
        .I2(\CD[0].col_reg[3][6] ),
        .I3(\CD[0].col_reg[3][4] ),
        .O(isomorphism_return076_out));
  LUT6 #(
    .INIT(64'hF00F0FF066996699)) 
    \base_new_pp[1]_i_1__2 
       (.I0(\CD[0].col_reg[3][4] ),
        .I1(\CD[0].col_reg[3][3] ),
        .I2(\CD[0].col_reg[3][6] ),
        .I3(\CD[0].col_reg[3][0] ),
        .I4(\CD[0].col_reg[3][5] ),
        .I5(enc_dec_sbox),
        .O(p_0_in));
  LUT5 #(
    .INIT(32'h8BB8B88B)) 
    \base_new_pp[2]_i_1__2 
       (.I0(\CD[0].col_reg[3][0] ),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][2] ),
        .I3(\CD[0].col_reg[3][5] ),
        .I4(\CD[0].col_reg[3][7] ),
        .O(p_0_in9_in));
  LUT6 #(
    .INIT(64'h1DD1E22EE22E1DD1)) 
    \base_new_pp[3]_i_1__2 
       (.I0(\CD[0].col_reg[3][6] ),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][1] ),
        .I3(p_72_in),
        .I4(\CD[0].col_reg[3][7] ),
        .I5(\CD[0].col_reg[3][4] ),
        .O(p_1_in17_in));
  LUT6 #(
    .INIT(64'h011101110111FEEE)) 
    \base_new_pp[3]_i_2__2 
       (.I0(\CD[2].col_reg[1][0] ),
        .I1(\info_o[31]_INST_0_i_22_n_0 ),
        .I2(\base_new_pp_reg[2]_0 [0]),
        .I3(\base_new_pp_reg[4]_2 ),
        .I4(\CD[2].col_reg[1][3] ),
        .I5(\base_new_pp_reg[3]_0 ),
        .O(p_72_in));
  LUT6 #(
    .INIT(64'hF00F66660FF09999)) 
    \base_new_pp[4]_i_1__2 
       (.I0(\CD[0].col_reg[3][3] ),
        .I1(\CD[0].col_reg[3][1] ),
        .I2(\CD[0].col_reg[3][5] ),
        .I3(\CD[0].col_reg[3][7] ),
        .I4(enc_dec_sbox),
        .I5(isomorphism_return277_out),
        .O(\base_new_pp[4]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'h011101110111FEEE)) 
    \base_new_pp[4]_i_2__2 
       (.I0(\CD[2].col_reg[1][0] ),
        .I1(\info_o[31]_INST_0_i_22_n_0 ),
        .I2(\base_new_pp_reg[2]_0 [0]),
        .I3(\base_new_pp_reg[4]_2 ),
        .I4(\CD[2].col_reg[1][6] ),
        .I5(\base_new_pp_reg[4]_3 ),
        .O(isomorphism_return277_out));
  LUT6 #(
    .INIT(64'h69966996FF0000FF)) 
    \base_new_pp[5]_i_1__2 
       (.I0(\CD[0].col_reg[3][1] ),
        .I1(\CD[0].col_reg[3][5] ),
        .I2(\CD[0].col_reg[3][0] ),
        .I3(\CD[0].col_reg[3][6] ),
        .I4(\CD[0].col_reg[3][4] ),
        .I5(enc_dec_sbox),
        .O(p_1_in7_in));
  LUT6 #(
    .INIT(64'h3CC3C33CA55A5AA5)) 
    \base_new_pp[6]_i_1__2 
       (.I0(\CD[0].col_reg[3][1] ),
        .I1(\CD[0].col_reg[3][5] ),
        .I2(\CD[0].col_reg[3][0] ),
        .I3(\CD[0].col_reg[3][6] ),
        .I4(\CD[0].col_reg[3][4] ),
        .I5(enc_dec_sbox),
        .O(p_1_in10_in));
  LUT6 #(
    .INIT(64'h3CC36666C33C6666)) 
    \base_new_pp[7]_i_1__2 
       (.I0(\CD[0].col_reg[3][4] ),
        .I1(\CD[0].col_reg[3][7] ),
        .I2(\CD[0].col_reg[3][5] ),
        .I3(\CD[0].col_reg[3][2] ),
        .I4(enc_dec_sbox),
        .I5(isomorphism_return179_out_16),
        .O(p_1_in18_in));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\base_new_pp[0]_i_1__2_n_0 ),
        .Q(\base_new_pp_reg_n_0_[0] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in),
        .Q(\base_new_pp_reg_n_0_[1] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in9_in),
        .Q(in21_in[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in17_in),
        .Q(in21_in[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\base_new_pp[4]_i_1__2_n_0 ),
        .Q(\base_new_pp_reg_n_0_[4] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in7_in),
        .Q(\base_new_pp_reg_n_0_[5] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in10_in),
        .Q(in2[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in18_in),
        .Q(in2[1]),
        .R(1'b0));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[28]_INST_0_i_13 
       (.I0(\info_o[31]_INST_0_i_11_0 [3]),
        .I1(\info_o[28]_INST_0_i_7_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_11_1 [3]),
        .I4(\info_o[31]_INST_0_i_11_2 [3]),
        .I5(\info_o[28]_INST_0_i_7_1 ),
        .O(\info_o[28]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[28]_INST_0_i_14 
       (.I0(\CD[0].col[3][7]_i_9 [3]),
        .I1(\CD[0].col[3][7]_i_9_0 ),
        .I2(\CD[0].col[3][7]_i_9_1 [3]),
        .I3(\CD[0].col[3][7]_i_9_2 ),
        .O(\CD[2].col_reg[1][3] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[28]_INST_0_i_15 
       (.I0(\info_o[31]_INST_0_i_11_0 [4]),
        .I1(\info_o[28]_INST_0_i_7_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_11_1 [4]),
        .I4(\info_o[31]_INST_0_i_11_2 [4]),
        .I5(\info_o[28]_INST_0_i_7_1 ),
        .O(\info_o[28]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[28]_INST_0_i_16 
       (.I0(\CD[0].col[3][7]_i_9 [4]),
        .I1(\CD[0].col[3][7]_i_9_0 ),
        .I2(\CD[0].col[3][7]_i_9_1 [4]),
        .I3(\CD[0].col[3][7]_i_9_2 ),
        .O(\CD[2].col_reg[1][4] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[28]_INST_0_i_6 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [3]),
        .I2(\info_o[28]_INST_0_i_13_n_0 ),
        .I3(\CD[2].col_reg[1][3] ),
        .O(\CD[0].col_reg[3][3] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[28]_INST_0_i_7 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [4]),
        .I2(\info_o[28]_INST_0_i_15_n_0 ),
        .I3(\CD[2].col_reg[1][4] ),
        .O(\CD[0].col_reg[3][4] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[29]_INST_0_i_13 
       (.I0(\info_o[31]_INST_0_i_11_0 [2]),
        .I1(\info_o[28]_INST_0_i_7_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_11_1 [2]),
        .I4(\info_o[31]_INST_0_i_11_2 [2]),
        .I5(\info_o[28]_INST_0_i_7_1 ),
        .O(\info_o[29]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[29]_INST_0_i_14 
       (.I0(\CD[0].col[3][7]_i_9 [2]),
        .I1(\CD[0].col[3][7]_i_9_0 ),
        .I2(\CD[0].col[3][7]_i_9_1 [2]),
        .I3(\CD[0].col[3][7]_i_9_2 ),
        .O(\CD[2].col_reg[1][2] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[29]_INST_0_i_15 
       (.I0(\info_o[31]_INST_0_i_11_0 [5]),
        .I1(\info_o[28]_INST_0_i_7_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_11_1 [5]),
        .I4(\info_o[31]_INST_0_i_11_2 [5]),
        .I5(\info_o[28]_INST_0_i_7_1 ),
        .O(\info_o[29]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[29]_INST_0_i_16 
       (.I0(\CD[0].col[3][7]_i_9 [5]),
        .I1(\CD[0].col[3][7]_i_9_0 ),
        .I2(\CD[0].col[3][7]_i_9_1 [5]),
        .I3(\CD[0].col[3][7]_i_9_2 ),
        .O(\CD[2].col_reg[1][5] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[29]_INST_0_i_6 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [2]),
        .I2(\info_o[29]_INST_0_i_13_n_0 ),
        .I3(\CD[2].col_reg[1][2] ),
        .O(\CD[0].col_reg[3][2] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[29]_INST_0_i_7 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [5]),
        .I2(\info_o[29]_INST_0_i_15_n_0 ),
        .I3(\CD[2].col_reg[1][5] ),
        .O(\CD[0].col_reg[3][5] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[30]_INST_0_i_13 
       (.I0(\info_o[31]_INST_0_i_11_0 [1]),
        .I1(\info_o[28]_INST_0_i_7_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_11_1 [1]),
        .I4(\info_o[31]_INST_0_i_11_2 [1]),
        .I5(\info_o[28]_INST_0_i_7_1 ),
        .O(\info_o[30]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[30]_INST_0_i_14 
       (.I0(\CD[0].col[3][7]_i_9 [1]),
        .I1(\CD[0].col[3][7]_i_9_0 ),
        .I2(\CD[0].col[3][7]_i_9_1 [1]),
        .I3(\CD[0].col[3][7]_i_9_2 ),
        .O(\CD[2].col_reg[1][1] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[30]_INST_0_i_15 
       (.I0(\info_o[31]_INST_0_i_11_0 [6]),
        .I1(\info_o[28]_INST_0_i_7_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_11_1 [6]),
        .I4(\info_o[31]_INST_0_i_11_2 [6]),
        .I5(\info_o[28]_INST_0_i_7_1 ),
        .O(\info_o[30]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[30]_INST_0_i_16 
       (.I0(\CD[0].col[3][7]_i_9 [6]),
        .I1(\CD[0].col[3][7]_i_9_0 ),
        .I2(\CD[0].col[3][7]_i_9_1 [6]),
        .I3(\CD[0].col[3][7]_i_9_2 ),
        .O(\CD[2].col_reg[1][6] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[30]_INST_0_i_6 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [1]),
        .I2(\info_o[30]_INST_0_i_13_n_0 ),
        .I3(\CD[2].col_reg[1][1] ),
        .O(\CD[0].col_reg[3][1] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[30]_INST_0_i_7 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [6]),
        .I2(\info_o[30]_INST_0_i_15_n_0 ),
        .I3(\CD[2].col_reg[1][6] ),
        .O(\CD[0].col_reg[3][6] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[31]_INST_0_i_10 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [0]),
        .I2(\info_o[31]_INST_0_i_22_n_0 ),
        .I3(\CD[2].col_reg[1][0] ),
        .O(\CD[0].col_reg[3][0] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[31]_INST_0_i_11 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [7]),
        .I2(\info_o[31]_INST_0_i_24_n_0 ),
        .I3(\CD[2].col_reg[1][7] ),
        .O(\CD[0].col_reg[3][7] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[31]_INST_0_i_22 
       (.I0(\info_o[31]_INST_0_i_11_0 [0]),
        .I1(\info_o[28]_INST_0_i_7_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_11_1 [0]),
        .I4(\info_o[31]_INST_0_i_11_2 [0]),
        .I5(\info_o[28]_INST_0_i_7_1 ),
        .O(\info_o[31]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[31]_INST_0_i_23 
       (.I0(\CD[0].col[3][7]_i_9 [0]),
        .I1(\CD[0].col[3][7]_i_9_0 ),
        .I2(\CD[0].col[3][7]_i_9_1 [0]),
        .I3(\CD[0].col[3][7]_i_9_2 ),
        .O(\CD[2].col_reg[1][0] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[31]_INST_0_i_24 
       (.I0(\info_o[31]_INST_0_i_11_0 [7]),
        .I1(\info_o[28]_INST_0_i_7_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_11_1 [7]),
        .I4(\info_o[31]_INST_0_i_11_2 [7]),
        .I5(\info_o[28]_INST_0_i_7_1 ),
        .O(\info_o[31]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[31]_INST_0_i_25 
       (.I0(\CD[0].col[3][7]_i_9 [7]),
        .I1(\CD[0].col[3][7]_i_9_0 ),
        .I2(\CD[0].col[3][7]_i_9_1 [7]),
        .I3(\CD[0].col[3][7]_i_9_2 ),
        .O(\CD[2].col_reg[1][7] ));
  LUT6 #(
    .INIT(64'hA9A69A955659656A)) 
    \out_gf_pp[0]_i_1__2 
       (.I0(gf_inv_8_stage1_return2__0),
        .I1(p_1_in7_in),
        .I2(p_0_in),
        .I3(\base_new_pp[4]_i_1__2_n_0 ),
        .I4(\base_new_pp[0]_i_1__2_n_0 ),
        .I5(gf_inv_8_stage1_return1__0),
        .O(gf_inv_8_stage1_return[0]));
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT4 #(
    .INIT(16'hF99F)) 
    \out_gf_pp[0]_i_2__2 
       (.I0(p_1_in18_in),
        .I1(p_1_in7_in),
        .I2(p_1_in17_in),
        .I3(p_0_in),
        .O(gf_inv_8_stage1_return2__0));
  LUT6 #(
    .INIT(64'h9999969699666996)) 
    \out_gf_pp[1]_i_1__2 
       (.I0(gf_inv_8_stage1_return1__0),
        .I1(gf_inv_8_stage1_return349_in),
        .I2(\out_gf_pp[1]_i_3__2_n_0 ),
        .I3(\out_gf_pp[3]_i_5__2_n_0 ),
        .I4(\out_gf_pp[3]_i_6__2_n_0 ),
        .I5(\out_gf_pp[1]_i_4__2_n_0 ),
        .O(gf_inv_8_stage1_return[1]));
  LUT6 #(
    .INIT(64'hF5C5FFCFFFCFFACA)) 
    \out_gf_pp[1]_i_2__2 
       (.I0(\CD[0].col_reg[3][6] ),
        .I1(\CD[0].col_reg[3][1] ),
        .I2(enc_dec_sbox),
        .I3(isomorphism_return114_out_17),
        .I4(p_72_in),
        .I5(\CD[0].col_reg[3][4] ),
        .O(gf_inv_8_stage1_return349_in));
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[1]_i_3__2 
       (.I0(\base_new_pp[4]_i_1__2_n_0 ),
        .I1(p_1_in7_in),
        .O(\out_gf_pp[1]_i_3__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[1]_i_4__2 
       (.I0(p_1_in18_in),
        .I1(p_1_in10_in),
        .O(\out_gf_pp[1]_i_4__2_n_0 ));
  LUT6 #(
    .INIT(64'h6A6A6A959595956A)) 
    \out_gf_pp[2]_i_1__2 
       (.I0(\out_gf_pp[2]_i_2__2_n_0 ),
        .I1(p_1_in10_in),
        .I2(p_0_in9_in),
        .I3(gf_inv_8_stage1_return542_out),
        .I4(gf_inv_8_stage1_return540_out),
        .I5(gf_inv_8_stage1_return1__0),
        .O(gf_inv_8_stage1_return[2]));
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT4 #(
    .INIT(16'hF99F)) 
    \out_gf_pp[2]_i_2__2 
       (.I0(p_0_in9_in),
        .I1(p_1_in17_in),
        .I2(p_1_in10_in),
        .I3(p_1_in18_in),
        .O(\out_gf_pp[2]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[2]_i_3__2 
       (.I0(p_1_in7_in),
        .I1(p_1_in18_in),
        .O(gf_inv_8_stage1_return542_out));
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[2]_i_4__2 
       (.I0(p_0_in),
        .I1(p_1_in17_in),
        .O(gf_inv_8_stage1_return540_out));
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT5 #(
    .INIT(32'hF9F9F99F)) 
    \out_gf_pp[2]_i_5__2 
       (.I0(p_1_in10_in),
        .I1(\base_new_pp[4]_i_1__2_n_0 ),
        .I2(p_0_in9_in),
        .I3(\out_gf_pp[2]_i_6__2_n_0 ),
        .I4(\out_gf_pp[2]_i_7__2_n_0 ),
        .O(gf_inv_8_stage1_return1__0));
  LUT6 #(
    .INIT(64'h9669000069960000)) 
    \out_gf_pp[2]_i_6__2 
       (.I0(\CD[0].col_reg[3][1] ),
        .I1(\CD[0].col_reg[3][0] ),
        .I2(\CD[0].col_reg[3][6] ),
        .I3(\CD[0].col_reg[3][3] ),
        .I4(enc_dec_sbox),
        .I5(\CD[0].col_reg[3][2] ),
        .O(\out_gf_pp[2]_i_6__2_n_0 ));
  LUT6 #(
    .INIT(64'h0000966900006996)) 
    \out_gf_pp[2]_i_7__2 
       (.I0(\CD[0].col_reg[3][5] ),
        .I1(\CD[0].col_reg[3][0] ),
        .I2(\CD[0].col_reg[3][6] ),
        .I3(\CD[0].col_reg[3][4] ),
        .I4(enc_dec_sbox),
        .I5(\CD[0].col_reg[3][1] ),
        .O(\out_gf_pp[2]_i_7__2_n_0 ));
  LUT6 #(
    .INIT(64'h5656565656A9A956)) 
    \out_gf_pp[3]_i_1__2 
       (.I0(\out_gf_pp[3]_i_2__2_n_0 ),
        .I1(gf_inv_8_stage1_return547_out),
        .I2(gf_inv_8_stage1_return546_out),
        .I3(\out_gf_pp[3]_i_5__2_n_0 ),
        .I4(\out_gf_pp[3]_i_6__2_n_0 ),
        .I5(\out_gf_pp[3]_i_7__2_n_0 ),
        .O(gf_inv_8_stage1_return[3]));
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT4 #(
    .INIT(16'hA6C0)) 
    \out_gf_pp[3]_i_2__2 
       (.I0(p_1_in18_in),
        .I1(p_1_in10_in),
        .I2(p_1_in17_in),
        .I3(p_0_in9_in),
        .O(\out_gf_pp[3]_i_2__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[3]_i_3__2 
       (.I0(\base_new_pp[4]_i_1__2_n_0 ),
        .I1(p_1_in10_in),
        .O(gf_inv_8_stage1_return547_out));
  LUT6 #(
    .INIT(64'hDE1212DE21EDED21)) 
    \out_gf_pp[3]_i_4__2 
       (.I0(isomorphism_return076_out),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][1] ),
        .I3(isomorphism_return1__0),
        .I4(\CD[0].col_reg[3][2] ),
        .I5(p_0_in9_in),
        .O(gf_inv_8_stage1_return546_out));
  LUT6 #(
    .INIT(64'hDE1212DE21EDED21)) 
    \out_gf_pp[3]_i_5__2 
       (.I0(isomorphism_return076_out),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][1] ),
        .I3(isomorphism_return1__0),
        .I4(\CD[0].col_reg[3][2] ),
        .I5(p_0_in),
        .O(\out_gf_pp[3]_i_5__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[3]_i_6__2 
       (.I0(p_1_in17_in),
        .I1(p_0_in9_in),
        .O(\out_gf_pp[3]_i_6__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \out_gf_pp[3]_i_7__2 
       (.I0(p_1_in10_in),
        .I1(p_1_in18_in),
        .I2(p_1_in7_in),
        .I3(\base_new_pp[4]_i_1__2_n_0 ),
        .O(\out_gf_pp[3]_i_7__2_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[0]),
        .Q(\out_gf_pp_reg_n_0_[0] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[1]),
        .Q(\out_gf_pp_reg_n_0_[1] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[2]),
        .Q(\out_gf_pp_reg_n_0_[2] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[3]),
        .Q(\out_gf_pp_reg_n_0_[3] ),
        .R(1'b0));
  LUT4 #(
    .INIT(16'h0F66)) 
    \sbox_pp2[0]_i_1 
       (.I0(sbox_out_dec),
        .I1(\sbox_pp2_reg[0] ),
        .I2(\base_new_pp_reg[1]_0 ),
        .I3(\sbox_pp2_reg[7] ),
        .O(D[0]));
  LUT5 #(
    .INIT(32'h00FF9696)) 
    \sbox_pp2[1]_i_1 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(p_1_in),
        .I2(\sbox_pp2_reg[1] ),
        .I3(\base_new_pp_reg[4]_0 ),
        .I4(\sbox_pp2_reg[7] ),
        .O(D[1]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[1]_i_2 
       (.I0(\base_new_pp_reg_n_0_[0] ),
        .I1(gf_muls_20_return__1[0]),
        .I2(gf_muls_20_return__1[1]),
        .I3(\base_new_pp_reg_n_0_[1] ),
        .I4(gf_muls_scl_2_return[1]),
        .O(p_1_in));
  LUT5 #(
    .INIT(32'hFF960096)) 
    \sbox_pp2[2]_i_1 
       (.I0(\base_new_pp_reg[4]_0 ),
        .I1(gf_inv_8_stage2_return013_out[1]),
        .I2(\sbox_pp2_reg[2] ),
        .I3(\sbox_pp2_reg[7] ),
        .I4(sbox_out_enc[0]),
        .O(D[2]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[2]_i_2 
       (.I0(in21_in[0]),
        .I1(in1__0[0]),
        .I2(in1__0[1]),
        .I3(in21_in[1]),
        .I4(gf_muls_scl_2_return[1]),
        .O(gf_inv_8_stage2_return013_out[1]));
  LUT6 #(
    .INIT(64'h0FF0666669960000)) 
    \sbox_pp2[2]_i_4 
       (.I0(in21_in[1]),
        .I1(\base_new_pp_reg_n_0_[1] ),
        .I2(in21_in[0]),
        .I3(\base_new_pp_reg_n_0_[0] ),
        .I4(in111_out[1]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_2_return[1]));
  LUT6 #(
    .INIT(64'hFFFF966900009669)) 
    \sbox_pp2[3]_i_1 
       (.I0(\base_new_pp_reg[6]_2 ),
        .I1(sbox_out_dec),
        .I2(\base_new_pp_reg[1]_0 ),
        .I3(\sbox_pp2_reg[3] ),
        .I4(\sbox_pp2_reg[7] ),
        .I5(sbox_out_enc[1]),
        .O(D[3]));
  LUT5 #(
    .INIT(32'h00FF9696)) 
    \sbox_pp2[4]_i_1 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(gf_inv_8_stage2_return013_out[0]),
        .I2(\sbox_pp2_reg[4] ),
        .I3(\base_new_pp_reg[6]_0 ),
        .I4(\sbox_pp2_reg[7] ),
        .O(D[4]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[4]_i_2 
       (.I0(in21_in[1]),
        .I1(in1__0[1]),
        .I2(in1__0[0]),
        .I3(in21_in[0]),
        .I4(gf_muls_scl_2_return[0]),
        .O(gf_inv_8_stage2_return013_out[0]));
  LUT5 #(
    .INIT(32'h00FF9669)) 
    \sbox_pp2[5]_i_1 
       (.I0(\base_new_pp_reg[6]_0 ),
        .I1(sbox_out_dec),
        .I2(\sbox_pp2_reg[5] ),
        .I3(\base_new_pp_reg[4]_1 ),
        .I4(\sbox_pp2_reg[7] ),
        .O(D[5]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[5]_i_2 
       (.I0(in2[1]),
        .I1(in1__0[1]),
        .I2(in1__0[0]),
        .I3(in2[0]),
        .I4(gf_muls_scl_20_return[0]),
        .O(sbox_out_dec));
  LUT6 #(
    .INIT(64'h0000FFFF96699669)) 
    \sbox_pp2[6]_i_1 
       (.I0(\base_new_pp_reg[6]_0 ),
        .I1(\base_new_pp_reg[4]_1 ),
        .I2(gf_inv_8_stage2_return0__3),
        .I3(\sbox_pp2_reg[6] ),
        .I4(\base_new_pp_reg[6]_1 ),
        .I5(\sbox_pp2_reg[7] ),
        .O(D[6]));
  LUT5 #(
    .INIT(32'h00FF9696)) 
    \sbox_pp2[7]_i_1 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(p_0_in2_in),
        .I2(\sbox_pp2_reg[7]_0 ),
        .I3(\base_new_pp_reg[6]_2 ),
        .I4(\sbox_pp2_reg[7] ),
        .O(D[7]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[7]_i_2 
       (.I0(\base_new_pp_reg_n_0_[4] ),
        .I1(gf_muls_20_return__1[0]),
        .I2(gf_muls_20_return__1[1]),
        .I3(\base_new_pp_reg_n_0_[5] ),
        .I4(gf_muls_scl_20_return[1]),
        .O(gf_inv_8_stage2_return0__3));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[7]_i_3 
       (.I0(\base_new_pp_reg_n_0_[1] ),
        .I1(gf_muls_20_return__1[1]),
        .I2(gf_muls_20_return__1[0]),
        .I3(\base_new_pp_reg_n_0_[0] ),
        .I4(gf_muls_scl_2_return[0]),
        .O(p_0_in2_in));
  LUT6 #(
    .INIT(64'h609F9F6060606060)) 
    \sbox_pp2[7]_i_4 
       (.I0(\base_new_pp_reg_n_0_[1] ),
        .I1(in21_in[1]),
        .I2(in111_out[1]),
        .I3(\base_new_pp_reg_n_0_[0] ),
        .I4(in21_in[0]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_2_return[0]));
endmodule

(* ORIG_REF_NAME = "sBox_8" *) 
module switch_elements_sBox_8_1
   (D,
    \base_new_pp_reg[4]_0 ,
    sbox_out_enc,
    \base_new_pp_reg[6]_0 ,
    \base_new_pp_reg[4]_1 ,
    \base_new_pp_reg[6]_1 ,
    \base_new_pp_reg[6]_2 ,
    \base_new_pp_reg[1]_0 ,
    \KR[3].key_host_reg[0][15] ,
    \CD[0].col_reg[3][15] ,
    \CD[2].col_reg[1][15] ,
    \CD[0].col_reg[3][14] ,
    \CD[2].col_reg[1][14] ,
    \CD[0].col_reg[3][13] ,
    \CD[2].col_reg[1][13] ,
    \CD[0].col_reg[3][12] ,
    \CD[2].col_reg[1][12] ,
    \CD[0].col_reg[3][11] ,
    \CD[2].col_reg[1][11] ,
    \CD[0].col_reg[3][10] ,
    \CD[2].col_reg[1][10] ,
    \CD[0].col_reg[3][9] ,
    \CD[2].col_reg[1][9] ,
    \CD[0].col_reg[3][8] ,
    \CD[2].col_reg[1][8] ,
    \sbox_pp2_reg[10] ,
    \sbox_pp2_reg[15] ,
    \sbox_pp2_reg[14] ,
    \sbox_pp2_reg[11] ,
    \sbox_pp2_reg[12] ,
    \sbox_pp2_reg[9] ,
    \sbox_pp2_reg[15]_0 ,
    key_en,
    \KR[3].key_reg[0][15] ,
    enable_i,
    key_sel_mux,
    \KR[3].key_reg[0][15]_0 ,
    \sbox_pp2_reg[13] ,
    \sbox_pp2_reg[8] ,
    \base_new_pp_reg[4]_2 ,
    \base_new_pp_reg[2]_0 ,
    \info_o[31]_INST_0_i_8_0 ,
    \base_new_pp[4]_i_2__1_0 ,
    enc_dec_sbox,
    \info_o[31]_INST_0_i_8_1 ,
    \info_o[31]_INST_0_i_8_2 ,
    \base_new_pp[4]_i_2__1_1 ,
    \CD[0].col[3][15]_i_7 ,
    \CD[0].col[3][15]_i_7_0 ,
    \CD[0].col[3][15]_i_7_1 ,
    \CD[0].col[3][15]_i_7_2 ,
    isomorphism_return179_out_14,
    isomorphism_return114_out_15,
    \base_new_pp_reg[4]_3 ,
    \base_new_pp_reg[3]_0 ,
    clk_i);
  output [7:0]D;
  output \base_new_pp_reg[4]_0 ;
  output [1:0]sbox_out_enc;
  output \base_new_pp_reg[6]_0 ;
  output \base_new_pp_reg[4]_1 ;
  output \base_new_pp_reg[6]_1 ;
  output \base_new_pp_reg[6]_2 ;
  output \base_new_pp_reg[1]_0 ;
  output [7:0]\KR[3].key_host_reg[0][15] ;
  output \CD[0].col_reg[3][15] ;
  output \CD[2].col_reg[1][15] ;
  output \CD[0].col_reg[3][14] ;
  output \CD[2].col_reg[1][14] ;
  output \CD[0].col_reg[3][13] ;
  output \CD[2].col_reg[1][13] ;
  output \CD[0].col_reg[3][12] ;
  output \CD[2].col_reg[1][12] ;
  output \CD[0].col_reg[3][11] ;
  output \CD[2].col_reg[1][11] ;
  output \CD[0].col_reg[3][10] ;
  output \CD[2].col_reg[1][10] ;
  output \CD[0].col_reg[3][9] ;
  output \CD[2].col_reg[1][9] ;
  output \CD[0].col_reg[3][8] ;
  output \CD[2].col_reg[1][8] ;
  input \sbox_pp2_reg[10] ;
  input \sbox_pp2_reg[15] ;
  input \sbox_pp2_reg[14] ;
  input \sbox_pp2_reg[11] ;
  input \sbox_pp2_reg[12] ;
  input \sbox_pp2_reg[9] ;
  input \sbox_pp2_reg[15]_0 ;
  input [0:0]key_en;
  input [7:0]\KR[3].key_reg[0][15] ;
  input [7:0]enable_i;
  input key_sel_mux;
  input [7:0]\KR[3].key_reg[0][15]_0 ;
  input \sbox_pp2_reg[13] ;
  input \sbox_pp2_reg[8] ;
  input \base_new_pp_reg[4]_2 ;
  input [7:0]\base_new_pp_reg[2]_0 ;
  input [7:0]\info_o[31]_INST_0_i_8_0 ;
  input \base_new_pp[4]_i_2__1_0 ;
  input enc_dec_sbox;
  input [7:0]\info_o[31]_INST_0_i_8_1 ;
  input [7:0]\info_o[31]_INST_0_i_8_2 ;
  input \base_new_pp[4]_i_2__1_1 ;
  input [7:0]\CD[0].col[3][15]_i_7 ;
  input \CD[0].col[3][15]_i_7_0 ;
  input [7:0]\CD[0].col[3][15]_i_7_1 ;
  input \CD[0].col[3][15]_i_7_2 ;
  input isomorphism_return179_out_14;
  input isomorphism_return114_out_15;
  input \base_new_pp_reg[4]_3 ;
  input \base_new_pp_reg[3]_0 ;
  input clk_i;

  wire [7:0]\CD[0].col[3][15]_i_7 ;
  wire \CD[0].col[3][15]_i_7_0 ;
  wire [7:0]\CD[0].col[3][15]_i_7_1 ;
  wire \CD[0].col[3][15]_i_7_2 ;
  wire \CD[0].col_reg[3][10] ;
  wire \CD[0].col_reg[3][11] ;
  wire \CD[0].col_reg[3][12] ;
  wire \CD[0].col_reg[3][13] ;
  wire \CD[0].col_reg[3][14] ;
  wire \CD[0].col_reg[3][15] ;
  wire \CD[0].col_reg[3][8] ;
  wire \CD[0].col_reg[3][9] ;
  wire \CD[2].col_reg[1][10] ;
  wire \CD[2].col_reg[1][11] ;
  wire \CD[2].col_reg[1][12] ;
  wire \CD[2].col_reg[1][13] ;
  wire \CD[2].col_reg[1][14] ;
  wire \CD[2].col_reg[1][15] ;
  wire \CD[2].col_reg[1][8] ;
  wire \CD[2].col_reg[1][9] ;
  wire [7:0]D;
  wire [7:0]\KR[3].key_host_reg[0][15] ;
  wire [7:0]\KR[3].key_reg[0][15] ;
  wire [7:0]\KR[3].key_reg[0][15]_0 ;
  wire \base_new_pp[0]_i_1__1_n_0 ;
  wire \base_new_pp[4]_i_1__1_n_0 ;
  wire \base_new_pp[4]_i_2__1_0 ;
  wire \base_new_pp[4]_i_2__1_1 ;
  wire \base_new_pp_reg[1]_0 ;
  wire [7:0]\base_new_pp_reg[2]_0 ;
  wire \base_new_pp_reg[3]_0 ;
  wire \base_new_pp_reg[4]_0 ;
  wire \base_new_pp_reg[4]_1 ;
  wire \base_new_pp_reg[4]_2 ;
  wire \base_new_pp_reg[4]_3 ;
  wire \base_new_pp_reg[6]_0 ;
  wire \base_new_pp_reg[6]_1 ;
  wire \base_new_pp_reg[6]_2 ;
  wire \base_new_pp_reg_n_0_[0] ;
  wire \base_new_pp_reg_n_0_[1] ;
  wire \base_new_pp_reg_n_0_[4] ;
  wire \base_new_pp_reg_n_0_[5] ;
  wire clk_i;
  wire [7:0]enable_i;
  wire enc_dec_sbox;
  wire [3:0]gf_inv_8_stage1_return;
  wire gf_inv_8_stage1_return1__0;
  wire gf_inv_8_stage1_return2__0;
  wire gf_inv_8_stage1_return349_in;
  wire gf_inv_8_stage1_return540_out;
  wire gf_inv_8_stage1_return542_out;
  wire gf_inv_8_stage1_return546_out;
  wire gf_inv_8_stage1_return547_out;
  wire [1:0]gf_inv_8_stage2_return013_out;
  wire [1:1]gf_inv_8_stage2_return0__3;
  wire [1:0]gf_muls_20_return__1;
  wire [1:0]gf_muls_scl_20_return;
  wire [1:0]gf_muls_scl_2_return;
  wire [1:0]in111_out;
  wire [1:0]in1__0;
  wire [1:0]in2;
  wire [1:0]in21_in;
  wire \info_o[24]_INST_0_i_7_n_0 ;
  wire \info_o[25]_INST_0_i_7_n_0 ;
  wire \info_o[26]_INST_0_i_7_n_0 ;
  wire \info_o[27]_INST_0_i_7_n_0 ;
  wire \info_o[28]_INST_0_i_9_n_0 ;
  wire \info_o[29]_INST_0_i_9_n_0 ;
  wire \info_o[30]_INST_0_i_9_n_0 ;
  wire \info_o[31]_INST_0_i_18_n_0 ;
  wire [7:0]\info_o[31]_INST_0_i_8_0 ;
  wire [7:0]\info_o[31]_INST_0_i_8_1 ;
  wire [7:0]\info_o[31]_INST_0_i_8_2 ;
  wire isomorphism_return076_out;
  wire isomorphism_return114_out_15;
  wire isomorphism_return179_out_14;
  wire isomorphism_return1__0;
  wire isomorphism_return277_out;
  wire [0:0]key_en;
  wire key_sel_mux;
  wire \out_gf_pp[1]_i_3__1_n_0 ;
  wire \out_gf_pp[1]_i_4__1_n_0 ;
  wire \out_gf_pp[2]_i_2__1_n_0 ;
  wire \out_gf_pp[2]_i_6__1_n_0 ;
  wire \out_gf_pp[2]_i_7__1_n_0 ;
  wire \out_gf_pp[3]_i_2__1_n_0 ;
  wire \out_gf_pp[3]_i_5__1_n_0 ;
  wire \out_gf_pp[3]_i_6__1_n_0 ;
  wire \out_gf_pp[3]_i_7__1_n_0 ;
  wire \out_gf_pp_reg_n_0_[0] ;
  wire \out_gf_pp_reg_n_0_[1] ;
  wire \out_gf_pp_reg_n_0_[2] ;
  wire \out_gf_pp_reg_n_0_[3] ;
  wire p_0_in;
  wire p_0_in2_in;
  wire p_0_in9_in;
  wire p_1_in;
  wire p_1_in10_in;
  wire p_1_in17_in;
  wire p_1_in18_in;
  wire p_1_in7_in;
  wire p_72_in;
  wire [8:8]sbox_out_dec;
  wire [1:0]sbox_out_enc;
  wire \sbox_pp2_reg[10] ;
  wire \sbox_pp2_reg[11] ;
  wire \sbox_pp2_reg[12] ;
  wire \sbox_pp2_reg[13] ;
  wire \sbox_pp2_reg[14] ;
  wire \sbox_pp2_reg[15] ;
  wire \sbox_pp2_reg[15]_0 ;
  wire \sbox_pp2_reg[8] ;
  wire \sbox_pp2_reg[9] ;

  LUT3 #(
    .INIT(8'h69)) 
    \KR[2].key[1][10]_i_3 
       (.I0(\base_new_pp_reg[6]_2 ),
        .I1(sbox_out_dec),
        .I2(\base_new_pp_reg[4]_1 ),
        .O(sbox_out_enc[0]));
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \KR[2].key[1][11]_i_3 
       (.I0(p_0_in2_in),
        .I1(gf_inv_8_stage2_return013_out[0]),
        .I2(\base_new_pp_reg[6]_0 ),
        .O(sbox_out_enc[1]));
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \KR[2].key[1][12]_i_3 
       (.I0(\base_new_pp_reg[6]_1 ),
        .I1(p_1_in),
        .O(\base_new_pp_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h96A59955695A66AA)) 
    \KR[2].key[1][13]_i_3 
       (.I0(gf_muls_scl_20_return[0]),
        .I1(\base_new_pp_reg_n_0_[4] ),
        .I2(gf_muls_20_return__1[0]),
        .I3(gf_muls_20_return__1[1]),
        .I4(\base_new_pp_reg_n_0_[5] ),
        .I5(gf_inv_8_stage2_return013_out[0]),
        .O(\base_new_pp_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h609F9F6060606060)) 
    \KR[2].key[1][13]_i_4 
       (.I0(\base_new_pp_reg_n_0_[5] ),
        .I1(in2[1]),
        .I2(in111_out[1]),
        .I3(\base_new_pp_reg_n_0_[4] ),
        .I4(in2[0]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_20_return[0]));
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT4 #(
    .INIT(16'hBE22)) 
    \KR[2].key[1][13]_i_5 
       (.I0(\out_gf_pp_reg_n_0_[2] ),
        .I1(\out_gf_pp_reg_n_0_[0] ),
        .I2(\out_gf_pp_reg_n_0_[1] ),
        .I3(\out_gf_pp_reg_n_0_[3] ),
        .O(gf_muls_20_return__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT4 #(
    .INIT(16'hDD82)) 
    \KR[2].key[1][13]_i_6 
       (.I0(\out_gf_pp_reg_n_0_[3] ),
        .I1(\out_gf_pp_reg_n_0_[1] ),
        .I2(\out_gf_pp_reg_n_0_[0] ),
        .I3(\out_gf_pp_reg_n_0_[2] ),
        .O(gf_muls_20_return__1[1]));
  LUT6 #(
    .INIT(64'hE4281BD71BD7E428)) 
    \KR[2].key[1][14]_i_3 
       (.I0(in2[0]),
        .I1(in1__0[0]),
        .I2(in1__0[1]),
        .I3(in2[1]),
        .I4(gf_muls_scl_20_return[1]),
        .I5(gf_inv_8_stage2_return013_out[1]),
        .O(\base_new_pp_reg[6]_1 ));
  LUT6 #(
    .INIT(64'h1BD7E428E4281BD7)) 
    \KR[2].key[1][15]_i_3 
       (.I0(in2[0]),
        .I1(in1__0[0]),
        .I2(in1__0[1]),
        .I3(in2[1]),
        .I4(gf_muls_scl_20_return[1]),
        .I5(p_1_in),
        .O(\base_new_pp_reg[6]_2 ));
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT4 #(
    .INIT(16'hB2E2)) 
    \KR[2].key[1][15]_i_4 
       (.I0(\out_gf_pp_reg_n_0_[0] ),
        .I1(\out_gf_pp_reg_n_0_[2] ),
        .I2(\out_gf_pp_reg_n_0_[1] ),
        .I3(\out_gf_pp_reg_n_0_[3] ),
        .O(in1__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT4 #(
    .INIT(16'hE4C6)) 
    \KR[2].key[1][15]_i_5 
       (.I0(\out_gf_pp_reg_n_0_[1] ),
        .I1(\out_gf_pp_reg_n_0_[0] ),
        .I2(\out_gf_pp_reg_n_0_[3] ),
        .I3(\out_gf_pp_reg_n_0_[2] ),
        .O(in1__0[1]));
  LUT6 #(
    .INIT(64'h0FF0666669960000)) 
    \KR[2].key[1][15]_i_6 
       (.I0(in2[1]),
        .I1(\base_new_pp_reg_n_0_[5] ),
        .I2(in2[0]),
        .I3(\base_new_pp_reg_n_0_[4] ),
        .I4(in111_out[1]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_20_return[1]));
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT4 #(
    .INIT(16'h23D6)) 
    \KR[2].key[1][15]_i_7 
       (.I0(\out_gf_pp_reg_n_0_[2] ),
        .I1(\out_gf_pp_reg_n_0_[3] ),
        .I2(\out_gf_pp_reg_n_0_[0] ),
        .I3(\out_gf_pp_reg_n_0_[1] ),
        .O(in111_out[1]));
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT4 #(
    .INIT(16'h6DB0)) 
    \KR[2].key[1][15]_i_8 
       (.I0(\out_gf_pp_reg_n_0_[3] ),
        .I1(\out_gf_pp_reg_n_0_[1] ),
        .I2(\out_gf_pp_reg_n_0_[2] ),
        .I3(\out_gf_pp_reg_n_0_[0] ),
        .O(in111_out[0]));
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \KR[2].key[1][8]_i_3 
       (.I0(p_0_in2_in),
        .I1(gf_inv_8_stage2_return013_out[0]),
        .I2(gf_inv_8_stage2_return0__3),
        .O(\base_new_pp_reg[1]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \KR[2].key[1][9]_i_3 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(p_1_in),
        .I2(p_0_in2_in),
        .O(\base_new_pp_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][10]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][15] [2]),
        .I2(enable_i[2]),
        .I3(key_sel_mux),
        .I4(sbox_out_enc[0]),
        .I5(\KR[3].key_reg[0][15]_0 [2]),
        .O(\KR[3].key_host_reg[0][15] [2]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][11]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][15] [3]),
        .I2(enable_i[3]),
        .I3(key_sel_mux),
        .I4(sbox_out_enc[1]),
        .I5(\KR[3].key_reg[0][15]_0 [3]),
        .O(\KR[3].key_host_reg[0][15] [3]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][12]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][15] [4]),
        .I2(enable_i[4]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[6]_0 ),
        .I5(\KR[3].key_reg[0][15]_0 [4]),
        .O(\KR[3].key_host_reg[0][15] [4]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][13]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][15] [5]),
        .I2(enable_i[5]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[4]_1 ),
        .I5(\KR[3].key_reg[0][15]_0 [5]),
        .O(\KR[3].key_host_reg[0][15] [5]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][14]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][15] [6]),
        .I2(enable_i[6]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[6]_1 ),
        .I5(\KR[3].key_reg[0][15]_0 [6]),
        .O(\KR[3].key_host_reg[0][15] [6]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][15]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][15] [7]),
        .I2(enable_i[7]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[6]_2 ),
        .I5(\KR[3].key_reg[0][15]_0 [7]),
        .O(\KR[3].key_host_reg[0][15] [7]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][8]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][15] [0]),
        .I2(enable_i[0]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[1]_0 ),
        .I5(\KR[3].key_reg[0][15]_0 [0]),
        .O(\KR[3].key_host_reg[0][15] [0]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][9]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][15] [1]),
        .I2(enable_i[1]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[4]_0 ),
        .I5(\KR[3].key_reg[0][15]_0 [1]),
        .O(\KR[3].key_host_reg[0][15] [1]));
  LUT5 #(
    .INIT(32'h66F0660F)) 
    \base_new_pp[0]_i_1__1 
       (.I0(\CD[0].col_reg[3][10] ),
        .I1(isomorphism_return1__0),
        .I2(\CD[0].col_reg[3][9] ),
        .I3(enc_dec_sbox),
        .I4(isomorphism_return076_out),
        .O(\base_new_pp[0]_i_1__1_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \base_new_pp[0]_i_2__1 
       (.I0(\CD[0].col_reg[3][9] ),
        .I1(\CD[0].col_reg[3][8] ),
        .I2(\CD[0].col_reg[3][14] ),
        .I3(\CD[0].col_reg[3][11] ),
        .O(isomorphism_return1__0));
  LUT4 #(
    .INIT(16'h9669)) 
    \base_new_pp[0]_i_3__1 
       (.I0(\CD[0].col_reg[3][13] ),
        .I1(\CD[0].col_reg[3][8] ),
        .I2(\CD[0].col_reg[3][14] ),
        .I3(\CD[0].col_reg[3][12] ),
        .O(isomorphism_return076_out));
  LUT6 #(
    .INIT(64'hF00F0FF066996699)) 
    \base_new_pp[1]_i_1__1 
       (.I0(\CD[0].col_reg[3][12] ),
        .I1(\CD[0].col_reg[3][11] ),
        .I2(\CD[0].col_reg[3][14] ),
        .I3(\CD[0].col_reg[3][8] ),
        .I4(\CD[0].col_reg[3][13] ),
        .I5(enc_dec_sbox),
        .O(p_0_in));
  LUT5 #(
    .INIT(32'h8BB8B88B)) 
    \base_new_pp[2]_i_1__1 
       (.I0(\CD[0].col_reg[3][8] ),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][10] ),
        .I3(\CD[0].col_reg[3][13] ),
        .I4(\CD[0].col_reg[3][15] ),
        .O(p_0_in9_in));
  LUT6 #(
    .INIT(64'h1DD1E22EE22E1DD1)) 
    \base_new_pp[3]_i_1__1 
       (.I0(\CD[0].col_reg[3][14] ),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][9] ),
        .I3(p_72_in),
        .I4(\CD[0].col_reg[3][15] ),
        .I5(\CD[0].col_reg[3][12] ),
        .O(p_1_in17_in));
  LUT6 #(
    .INIT(64'h011101110111FEEE)) 
    \base_new_pp[3]_i_2__1 
       (.I0(\CD[2].col_reg[1][8] ),
        .I1(\info_o[24]_INST_0_i_7_n_0 ),
        .I2(\base_new_pp_reg[2]_0 [0]),
        .I3(\base_new_pp_reg[4]_2 ),
        .I4(\CD[2].col_reg[1][11] ),
        .I5(\base_new_pp_reg[3]_0 ),
        .O(p_72_in));
  LUT6 #(
    .INIT(64'hF00F66660FF09999)) 
    \base_new_pp[4]_i_1__1 
       (.I0(\CD[0].col_reg[3][11] ),
        .I1(\CD[0].col_reg[3][9] ),
        .I2(\CD[0].col_reg[3][13] ),
        .I3(\CD[0].col_reg[3][15] ),
        .I4(enc_dec_sbox),
        .I5(isomorphism_return277_out),
        .O(\base_new_pp[4]_i_1__1_n_0 ));
  LUT6 #(
    .INIT(64'h011101110111FEEE)) 
    \base_new_pp[4]_i_2__1 
       (.I0(\CD[2].col_reg[1][8] ),
        .I1(\info_o[24]_INST_0_i_7_n_0 ),
        .I2(\base_new_pp_reg[2]_0 [0]),
        .I3(\base_new_pp_reg[4]_2 ),
        .I4(\CD[2].col_reg[1][14] ),
        .I5(\base_new_pp_reg[4]_3 ),
        .O(isomorphism_return277_out));
  LUT6 #(
    .INIT(64'h69966996FF0000FF)) 
    \base_new_pp[5]_i_1__1 
       (.I0(\CD[0].col_reg[3][9] ),
        .I1(\CD[0].col_reg[3][13] ),
        .I2(\CD[0].col_reg[3][8] ),
        .I3(\CD[0].col_reg[3][14] ),
        .I4(\CD[0].col_reg[3][12] ),
        .I5(enc_dec_sbox),
        .O(p_1_in7_in));
  LUT6 #(
    .INIT(64'h3CC3C33CA55A5AA5)) 
    \base_new_pp[6]_i_1__1 
       (.I0(\CD[0].col_reg[3][9] ),
        .I1(\CD[0].col_reg[3][13] ),
        .I2(\CD[0].col_reg[3][8] ),
        .I3(\CD[0].col_reg[3][14] ),
        .I4(\CD[0].col_reg[3][12] ),
        .I5(enc_dec_sbox),
        .O(p_1_in10_in));
  LUT6 #(
    .INIT(64'h3CC36666C33C6666)) 
    \base_new_pp[7]_i_1__1 
       (.I0(\CD[0].col_reg[3][12] ),
        .I1(\CD[0].col_reg[3][15] ),
        .I2(\CD[0].col_reg[3][13] ),
        .I3(\CD[0].col_reg[3][10] ),
        .I4(enc_dec_sbox),
        .I5(isomorphism_return179_out_14),
        .O(p_1_in18_in));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\base_new_pp[0]_i_1__1_n_0 ),
        .Q(\base_new_pp_reg_n_0_[0] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in),
        .Q(\base_new_pp_reg_n_0_[1] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in9_in),
        .Q(in21_in[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in17_in),
        .Q(in21_in[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\base_new_pp[4]_i_1__1_n_0 ),
        .Q(\base_new_pp_reg_n_0_[4] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in7_in),
        .Q(\base_new_pp_reg_n_0_[5] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in10_in),
        .Q(in2[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in18_in),
        .Q(in2[1]),
        .R(1'b0));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[24]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [0]),
        .I2(\info_o[24]_INST_0_i_7_n_0 ),
        .I3(\CD[2].col_reg[1][8] ),
        .O(\CD[0].col_reg[3][8] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[24]_INST_0_i_7 
       (.I0(\info_o[31]_INST_0_i_8_0 [0]),
        .I1(\base_new_pp[4]_i_2__1_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_8_1 [0]),
        .I4(\info_o[31]_INST_0_i_8_2 [0]),
        .I5(\base_new_pp[4]_i_2__1_1 ),
        .O(\info_o[24]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[24]_INST_0_i_8 
       (.I0(\CD[0].col[3][15]_i_7 [0]),
        .I1(\CD[0].col[3][15]_i_7_0 ),
        .I2(\CD[0].col[3][15]_i_7_1 [0]),
        .I3(\CD[0].col[3][15]_i_7_2 ),
        .O(\CD[2].col_reg[1][8] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[25]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [1]),
        .I2(\info_o[25]_INST_0_i_7_n_0 ),
        .I3(\CD[2].col_reg[1][9] ),
        .O(\CD[0].col_reg[3][9] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[25]_INST_0_i_7 
       (.I0(\info_o[31]_INST_0_i_8_0 [1]),
        .I1(\base_new_pp[4]_i_2__1_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_8_1 [1]),
        .I4(\info_o[31]_INST_0_i_8_2 [1]),
        .I5(\base_new_pp[4]_i_2__1_1 ),
        .O(\info_o[25]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[25]_INST_0_i_8 
       (.I0(\CD[0].col[3][15]_i_7 [1]),
        .I1(\CD[0].col[3][15]_i_7_0 ),
        .I2(\CD[0].col[3][15]_i_7_1 [1]),
        .I3(\CD[0].col[3][15]_i_7_2 ),
        .O(\CD[2].col_reg[1][9] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[26]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [2]),
        .I2(\info_o[26]_INST_0_i_7_n_0 ),
        .I3(\CD[2].col_reg[1][10] ),
        .O(\CD[0].col_reg[3][10] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[26]_INST_0_i_7 
       (.I0(\info_o[31]_INST_0_i_8_0 [2]),
        .I1(\base_new_pp[4]_i_2__1_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_8_1 [2]),
        .I4(\info_o[31]_INST_0_i_8_2 [2]),
        .I5(\base_new_pp[4]_i_2__1_1 ),
        .O(\info_o[26]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[26]_INST_0_i_8 
       (.I0(\CD[0].col[3][15]_i_7 [2]),
        .I1(\CD[0].col[3][15]_i_7_0 ),
        .I2(\CD[0].col[3][15]_i_7_1 [2]),
        .I3(\CD[0].col[3][15]_i_7_2 ),
        .O(\CD[2].col_reg[1][10] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[27]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [3]),
        .I2(\info_o[27]_INST_0_i_7_n_0 ),
        .I3(\CD[2].col_reg[1][11] ),
        .O(\CD[0].col_reg[3][11] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[27]_INST_0_i_7 
       (.I0(\info_o[31]_INST_0_i_8_0 [3]),
        .I1(\base_new_pp[4]_i_2__1_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_8_1 [3]),
        .I4(\info_o[31]_INST_0_i_8_2 [3]),
        .I5(\base_new_pp[4]_i_2__1_1 ),
        .O(\info_o[27]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[27]_INST_0_i_8 
       (.I0(\CD[0].col[3][15]_i_7 [3]),
        .I1(\CD[0].col[3][15]_i_7_0 ),
        .I2(\CD[0].col[3][15]_i_7_1 [3]),
        .I3(\CD[0].col[3][15]_i_7_2 ),
        .O(\CD[2].col_reg[1][11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[28]_INST_0_i_10 
       (.I0(\CD[0].col[3][15]_i_7 [4]),
        .I1(\CD[0].col[3][15]_i_7_0 ),
        .I2(\CD[0].col[3][15]_i_7_1 [4]),
        .I3(\CD[0].col[3][15]_i_7_2 ),
        .O(\CD[2].col_reg[1][12] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[28]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [4]),
        .I2(\info_o[28]_INST_0_i_9_n_0 ),
        .I3(\CD[2].col_reg[1][12] ),
        .O(\CD[0].col_reg[3][12] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[28]_INST_0_i_9 
       (.I0(\info_o[31]_INST_0_i_8_0 [4]),
        .I1(\base_new_pp[4]_i_2__1_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_8_1 [4]),
        .I4(\info_o[31]_INST_0_i_8_2 [4]),
        .I5(\base_new_pp[4]_i_2__1_1 ),
        .O(\info_o[28]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[29]_INST_0_i_10 
       (.I0(\CD[0].col[3][15]_i_7 [5]),
        .I1(\CD[0].col[3][15]_i_7_0 ),
        .I2(\CD[0].col[3][15]_i_7_1 [5]),
        .I3(\CD[0].col[3][15]_i_7_2 ),
        .O(\CD[2].col_reg[1][13] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[29]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [5]),
        .I2(\info_o[29]_INST_0_i_9_n_0 ),
        .I3(\CD[2].col_reg[1][13] ),
        .O(\CD[0].col_reg[3][13] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[29]_INST_0_i_9 
       (.I0(\info_o[31]_INST_0_i_8_0 [5]),
        .I1(\base_new_pp[4]_i_2__1_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_8_1 [5]),
        .I4(\info_o[31]_INST_0_i_8_2 [5]),
        .I5(\base_new_pp[4]_i_2__1_1 ),
        .O(\info_o[29]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[30]_INST_0_i_10 
       (.I0(\CD[0].col[3][15]_i_7 [6]),
        .I1(\CD[0].col[3][15]_i_7_0 ),
        .I2(\CD[0].col[3][15]_i_7_1 [6]),
        .I3(\CD[0].col[3][15]_i_7_2 ),
        .O(\CD[2].col_reg[1][14] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[30]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [6]),
        .I2(\info_o[30]_INST_0_i_9_n_0 ),
        .I3(\CD[2].col_reg[1][14] ),
        .O(\CD[0].col_reg[3][14] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[30]_INST_0_i_9 
       (.I0(\info_o[31]_INST_0_i_8_0 [6]),
        .I1(\base_new_pp[4]_i_2__1_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_8_1 [6]),
        .I4(\info_o[31]_INST_0_i_8_2 [6]),
        .I5(\base_new_pp[4]_i_2__1_1 ),
        .O(\info_o[30]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[31]_INST_0_i_18 
       (.I0(\info_o[31]_INST_0_i_8_0 [7]),
        .I1(\base_new_pp[4]_i_2__1_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_8_1 [7]),
        .I4(\info_o[31]_INST_0_i_8_2 [7]),
        .I5(\base_new_pp[4]_i_2__1_1 ),
        .O(\info_o[31]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[31]_INST_0_i_19 
       (.I0(\CD[0].col[3][15]_i_7 [7]),
        .I1(\CD[0].col[3][15]_i_7_0 ),
        .I2(\CD[0].col[3][15]_i_7_1 [7]),
        .I3(\CD[0].col[3][15]_i_7_2 ),
        .O(\CD[2].col_reg[1][15] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[31]_INST_0_i_8 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [7]),
        .I2(\info_o[31]_INST_0_i_18_n_0 ),
        .I3(\CD[2].col_reg[1][15] ),
        .O(\CD[0].col_reg[3][15] ));
  LUT6 #(
    .INIT(64'hA9A69A955659656A)) 
    \out_gf_pp[0]_i_1__1 
       (.I0(gf_inv_8_stage1_return2__0),
        .I1(p_1_in7_in),
        .I2(p_0_in),
        .I3(\base_new_pp[4]_i_1__1_n_0 ),
        .I4(\base_new_pp[0]_i_1__1_n_0 ),
        .I5(gf_inv_8_stage1_return1__0),
        .O(gf_inv_8_stage1_return[0]));
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT4 #(
    .INIT(16'hF99F)) 
    \out_gf_pp[0]_i_2__1 
       (.I0(p_1_in18_in),
        .I1(p_1_in7_in),
        .I2(p_1_in17_in),
        .I3(p_0_in),
        .O(gf_inv_8_stage1_return2__0));
  LUT6 #(
    .INIT(64'h9999969699666996)) 
    \out_gf_pp[1]_i_1__1 
       (.I0(gf_inv_8_stage1_return1__0),
        .I1(gf_inv_8_stage1_return349_in),
        .I2(\out_gf_pp[1]_i_3__1_n_0 ),
        .I3(\out_gf_pp[3]_i_5__1_n_0 ),
        .I4(\out_gf_pp[3]_i_6__1_n_0 ),
        .I5(\out_gf_pp[1]_i_4__1_n_0 ),
        .O(gf_inv_8_stage1_return[1]));
  LUT6 #(
    .INIT(64'hF5C5FFCFFFCFFACA)) 
    \out_gf_pp[1]_i_2__1 
       (.I0(\CD[0].col_reg[3][14] ),
        .I1(\CD[0].col_reg[3][9] ),
        .I2(enc_dec_sbox),
        .I3(isomorphism_return114_out_15),
        .I4(p_72_in),
        .I5(\CD[0].col_reg[3][12] ),
        .O(gf_inv_8_stage1_return349_in));
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[1]_i_3__1 
       (.I0(\base_new_pp[4]_i_1__1_n_0 ),
        .I1(p_1_in7_in),
        .O(\out_gf_pp[1]_i_3__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[1]_i_4__1 
       (.I0(p_1_in18_in),
        .I1(p_1_in10_in),
        .O(\out_gf_pp[1]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h6A6A6A959595956A)) 
    \out_gf_pp[2]_i_1__1 
       (.I0(\out_gf_pp[2]_i_2__1_n_0 ),
        .I1(p_1_in10_in),
        .I2(p_0_in9_in),
        .I3(gf_inv_8_stage1_return542_out),
        .I4(gf_inv_8_stage1_return540_out),
        .I5(gf_inv_8_stage1_return1__0),
        .O(gf_inv_8_stage1_return[2]));
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT4 #(
    .INIT(16'hF99F)) 
    \out_gf_pp[2]_i_2__1 
       (.I0(p_0_in9_in),
        .I1(p_1_in17_in),
        .I2(p_1_in10_in),
        .I3(p_1_in18_in),
        .O(\out_gf_pp[2]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[2]_i_3__1 
       (.I0(p_1_in7_in),
        .I1(p_1_in18_in),
        .O(gf_inv_8_stage1_return542_out));
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[2]_i_4__1 
       (.I0(p_0_in),
        .I1(p_1_in17_in),
        .O(gf_inv_8_stage1_return540_out));
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT5 #(
    .INIT(32'hF9F9F99F)) 
    \out_gf_pp[2]_i_5__1 
       (.I0(p_1_in10_in),
        .I1(\base_new_pp[4]_i_1__1_n_0 ),
        .I2(p_0_in9_in),
        .I3(\out_gf_pp[2]_i_6__1_n_0 ),
        .I4(\out_gf_pp[2]_i_7__1_n_0 ),
        .O(gf_inv_8_stage1_return1__0));
  LUT6 #(
    .INIT(64'h9669000069960000)) 
    \out_gf_pp[2]_i_6__1 
       (.I0(\CD[0].col_reg[3][9] ),
        .I1(\CD[0].col_reg[3][8] ),
        .I2(\CD[0].col_reg[3][14] ),
        .I3(\CD[0].col_reg[3][11] ),
        .I4(enc_dec_sbox),
        .I5(\CD[0].col_reg[3][10] ),
        .O(\out_gf_pp[2]_i_6__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000966900006996)) 
    \out_gf_pp[2]_i_7__1 
       (.I0(\CD[0].col_reg[3][13] ),
        .I1(\CD[0].col_reg[3][8] ),
        .I2(\CD[0].col_reg[3][14] ),
        .I3(\CD[0].col_reg[3][12] ),
        .I4(enc_dec_sbox),
        .I5(\CD[0].col_reg[3][9] ),
        .O(\out_gf_pp[2]_i_7__1_n_0 ));
  LUT6 #(
    .INIT(64'h5656565656A9A956)) 
    \out_gf_pp[3]_i_1__1 
       (.I0(\out_gf_pp[3]_i_2__1_n_0 ),
        .I1(gf_inv_8_stage1_return547_out),
        .I2(gf_inv_8_stage1_return546_out),
        .I3(\out_gf_pp[3]_i_5__1_n_0 ),
        .I4(\out_gf_pp[3]_i_6__1_n_0 ),
        .I5(\out_gf_pp[3]_i_7__1_n_0 ),
        .O(gf_inv_8_stage1_return[3]));
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT4 #(
    .INIT(16'hA6C0)) 
    \out_gf_pp[3]_i_2__1 
       (.I0(p_1_in18_in),
        .I1(p_1_in10_in),
        .I2(p_1_in17_in),
        .I3(p_0_in9_in),
        .O(\out_gf_pp[3]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[3]_i_3__1 
       (.I0(\base_new_pp[4]_i_1__1_n_0 ),
        .I1(p_1_in10_in),
        .O(gf_inv_8_stage1_return547_out));
  LUT6 #(
    .INIT(64'hDE1212DE21EDED21)) 
    \out_gf_pp[3]_i_4__1 
       (.I0(isomorphism_return076_out),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][9] ),
        .I3(isomorphism_return1__0),
        .I4(\CD[0].col_reg[3][10] ),
        .I5(p_0_in9_in),
        .O(gf_inv_8_stage1_return546_out));
  LUT6 #(
    .INIT(64'hDE1212DE21EDED21)) 
    \out_gf_pp[3]_i_5__1 
       (.I0(isomorphism_return076_out),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][9] ),
        .I3(isomorphism_return1__0),
        .I4(\CD[0].col_reg[3][10] ),
        .I5(p_0_in),
        .O(\out_gf_pp[3]_i_5__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[3]_i_6__1 
       (.I0(p_1_in17_in),
        .I1(p_0_in9_in),
        .O(\out_gf_pp[3]_i_6__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \out_gf_pp[3]_i_7__1 
       (.I0(p_1_in10_in),
        .I1(p_1_in18_in),
        .I2(p_1_in7_in),
        .I3(\base_new_pp[4]_i_1__1_n_0 ),
        .O(\out_gf_pp[3]_i_7__1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[0]),
        .Q(\out_gf_pp_reg_n_0_[0] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[1]),
        .Q(\out_gf_pp_reg_n_0_[1] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[2]),
        .Q(\out_gf_pp_reg_n_0_[2] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[3]),
        .Q(\out_gf_pp_reg_n_0_[3] ),
        .R(1'b0));
  LUT5 #(
    .INIT(32'hFF960096)) 
    \sbox_pp2[10]_i_1 
       (.I0(\base_new_pp_reg[4]_0 ),
        .I1(gf_inv_8_stage2_return013_out[1]),
        .I2(\sbox_pp2_reg[10] ),
        .I3(\sbox_pp2_reg[15] ),
        .I4(sbox_out_enc[0]),
        .O(D[2]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[10]_i_2 
       (.I0(in21_in[0]),
        .I1(in1__0[0]),
        .I2(in1__0[1]),
        .I3(in21_in[1]),
        .I4(gf_muls_scl_2_return[1]),
        .O(gf_inv_8_stage2_return013_out[1]));
  LUT6 #(
    .INIT(64'h0FF0666669960000)) 
    \sbox_pp2[10]_i_3 
       (.I0(in21_in[1]),
        .I1(\base_new_pp_reg_n_0_[1] ),
        .I2(in21_in[0]),
        .I3(\base_new_pp_reg_n_0_[0] ),
        .I4(in111_out[1]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_2_return[1]));
  LUT6 #(
    .INIT(64'hFFFF966900009669)) 
    \sbox_pp2[11]_i_1 
       (.I0(\base_new_pp_reg[6]_2 ),
        .I1(sbox_out_dec),
        .I2(\base_new_pp_reg[1]_0 ),
        .I3(\sbox_pp2_reg[11] ),
        .I4(\sbox_pp2_reg[15] ),
        .I5(sbox_out_enc[1]),
        .O(D[3]));
  LUT5 #(
    .INIT(32'h00FF9696)) 
    \sbox_pp2[12]_i_1 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(gf_inv_8_stage2_return013_out[0]),
        .I2(\sbox_pp2_reg[12] ),
        .I3(\base_new_pp_reg[6]_0 ),
        .I4(\sbox_pp2_reg[15] ),
        .O(D[4]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[12]_i_2 
       (.I0(in21_in[1]),
        .I1(in1__0[1]),
        .I2(in1__0[0]),
        .I3(in21_in[0]),
        .I4(gf_muls_scl_2_return[0]),
        .O(gf_inv_8_stage2_return013_out[0]));
  LUT5 #(
    .INIT(32'h00FF9669)) 
    \sbox_pp2[13]_i_1 
       (.I0(\base_new_pp_reg[6]_0 ),
        .I1(sbox_out_dec),
        .I2(\sbox_pp2_reg[13] ),
        .I3(\base_new_pp_reg[4]_1 ),
        .I4(\sbox_pp2_reg[15] ),
        .O(D[5]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[13]_i_2 
       (.I0(in2[1]),
        .I1(in1__0[1]),
        .I2(in1__0[0]),
        .I3(in2[0]),
        .I4(gf_muls_scl_20_return[0]),
        .O(sbox_out_dec));
  LUT6 #(
    .INIT(64'h0000FFFF96699669)) 
    \sbox_pp2[14]_i_1 
       (.I0(\base_new_pp_reg[6]_0 ),
        .I1(\base_new_pp_reg[4]_1 ),
        .I2(gf_inv_8_stage2_return0__3),
        .I3(\sbox_pp2_reg[14] ),
        .I4(\base_new_pp_reg[6]_1 ),
        .I5(\sbox_pp2_reg[15] ),
        .O(D[6]));
  LUT5 #(
    .INIT(32'h00FF9696)) 
    \sbox_pp2[15]_i_1 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(p_0_in2_in),
        .I2(\sbox_pp2_reg[15]_0 ),
        .I3(\base_new_pp_reg[6]_2 ),
        .I4(\sbox_pp2_reg[15] ),
        .O(D[7]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[15]_i_2 
       (.I0(\base_new_pp_reg_n_0_[4] ),
        .I1(gf_muls_20_return__1[0]),
        .I2(gf_muls_20_return__1[1]),
        .I3(\base_new_pp_reg_n_0_[5] ),
        .I4(gf_muls_scl_20_return[1]),
        .O(gf_inv_8_stage2_return0__3));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[15]_i_3 
       (.I0(\base_new_pp_reg_n_0_[1] ),
        .I1(gf_muls_20_return__1[1]),
        .I2(gf_muls_20_return__1[0]),
        .I3(\base_new_pp_reg_n_0_[0] ),
        .I4(gf_muls_scl_2_return[0]),
        .O(p_0_in2_in));
  LUT6 #(
    .INIT(64'h609F9F6060606060)) 
    \sbox_pp2[15]_i_4 
       (.I0(\base_new_pp_reg_n_0_[1] ),
        .I1(in21_in[1]),
        .I2(in111_out[1]),
        .I3(\base_new_pp_reg_n_0_[0] ),
        .I4(in21_in[0]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_2_return[0]));
  LUT4 #(
    .INIT(16'h0F66)) 
    \sbox_pp2[8]_i_1 
       (.I0(sbox_out_dec),
        .I1(\sbox_pp2_reg[8] ),
        .I2(\base_new_pp_reg[1]_0 ),
        .I3(\sbox_pp2_reg[15] ),
        .O(D[0]));
  LUT5 #(
    .INIT(32'h00FF9696)) 
    \sbox_pp2[9]_i_1 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(p_1_in),
        .I2(\sbox_pp2_reg[9] ),
        .I3(\base_new_pp_reg[4]_0 ),
        .I4(\sbox_pp2_reg[15] ),
        .O(D[1]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[9]_i_2 
       (.I0(\base_new_pp_reg_n_0_[0] ),
        .I1(gf_muls_20_return__1[0]),
        .I2(gf_muls_20_return__1[1]),
        .I3(\base_new_pp_reg_n_0_[1] ),
        .I4(gf_muls_scl_2_return[1]),
        .O(p_1_in));
endmodule

(* ORIG_REF_NAME = "sBox_8" *) 
module switch_elements_sBox_8_2
   (enable_i_0_sp_1,
    D,
    \base_new_pp_reg[4]_0 ,
    sbox_out_enc,
    \base_new_pp_reg[6]_0 ,
    \base_new_pp_reg[4]_1 ,
    \base_new_pp_reg[6]_1 ,
    \base_new_pp_reg[6]_2 ,
    \base_new_pp_reg[1]_0 ,
    \KR[3].key_host_reg[0][23] ,
    \CD[0].col_reg[3][23] ,
    \CD[2].col_reg[1][23] ,
    \CD[0].col_reg[3][22] ,
    \CD[2].col_reg[1][22] ,
    \CD[0].col_reg[3][21] ,
    \CD[2].col_reg[1][21] ,
    \CD[0].col_reg[3][20] ,
    \CD[2].col_reg[1][20] ,
    \CD[0].col_reg[3][19] ,
    \CD[2].col_reg[1][19] ,
    \CD[0].col_reg[3][18] ,
    \CD[2].col_reg[1][18] ,
    \CD[0].col_reg[3][17] ,
    \CD[2].col_reg[1][17] ,
    \CD[0].col_reg[3][16] ,
    \CD[2].col_reg[1][16] ,
    enable_i,
    \sbox_pp2_reg[18] ,
    \sbox_pp2_reg[23] ,
    \sbox_pp2_reg[22] ,
    \sbox_pp2_reg[19] ,
    \sbox_pp2_reg[20] ,
    \sbox_pp2_reg[17] ,
    \sbox_pp2_reg[23]_0 ,
    key_en,
    \KR[3].key_reg[0][23] ,
    key_sel_mux,
    \KR[3].key_reg[0][23]_0 ,
    \sbox_pp2_reg[21] ,
    \sbox_pp2_reg[16] ,
    \base_new_pp_reg[4]_2 ,
    \base_new_pp_reg[2]_0 ,
    \info_o[23]_INST_0_i_4_0 ,
    \base_new_pp[4]_i_2__0_0 ,
    enc_dec_sbox,
    \info_o[23]_INST_0_i_4_1 ,
    \info_o[23]_INST_0_i_4_2 ,
    \base_new_pp[4]_i_2__0_1 ,
    \CD[1].col[2][23]_i_3 ,
    \CD[1].col[2][23]_i_3_0 ,
    \CD[1].col[2][23]_i_3_1 ,
    \CD[1].col[2][23]_i_3_2 ,
    isomorphism_return179_out_12,
    isomorphism_return114_out_13,
    \base_new_pp_reg[4]_3 ,
    \base_new_pp_reg[3]_0 ,
    clk_i);
  output enable_i_0_sp_1;
  output [7:0]D;
  output \base_new_pp_reg[4]_0 ;
  output [1:0]sbox_out_enc;
  output \base_new_pp_reg[6]_0 ;
  output \base_new_pp_reg[4]_1 ;
  output \base_new_pp_reg[6]_1 ;
  output \base_new_pp_reg[6]_2 ;
  output \base_new_pp_reg[1]_0 ;
  output [7:0]\KR[3].key_host_reg[0][23] ;
  output \CD[0].col_reg[3][23] ;
  output \CD[2].col_reg[1][23] ;
  output \CD[0].col_reg[3][22] ;
  output \CD[2].col_reg[1][22] ;
  output \CD[0].col_reg[3][21] ;
  output \CD[2].col_reg[1][21] ;
  output \CD[0].col_reg[3][20] ;
  output \CD[2].col_reg[1][20] ;
  output \CD[0].col_reg[3][19] ;
  output \CD[2].col_reg[1][19] ;
  output \CD[0].col_reg[3][18] ;
  output \CD[2].col_reg[1][18] ;
  output \CD[0].col_reg[3][17] ;
  output \CD[2].col_reg[1][17] ;
  output \CD[0].col_reg[3][16] ;
  output \CD[2].col_reg[1][16] ;
  input [13:0]enable_i;
  input \sbox_pp2_reg[18] ;
  input \sbox_pp2_reg[23] ;
  input \sbox_pp2_reg[22] ;
  input \sbox_pp2_reg[19] ;
  input \sbox_pp2_reg[20] ;
  input \sbox_pp2_reg[17] ;
  input \sbox_pp2_reg[23]_0 ;
  input [0:0]key_en;
  input [7:0]\KR[3].key_reg[0][23] ;
  input key_sel_mux;
  input [7:0]\KR[3].key_reg[0][23]_0 ;
  input \sbox_pp2_reg[21] ;
  input \sbox_pp2_reg[16] ;
  input \base_new_pp_reg[4]_2 ;
  input [7:0]\base_new_pp_reg[2]_0 ;
  input [7:0]\info_o[23]_INST_0_i_4_0 ;
  input \base_new_pp[4]_i_2__0_0 ;
  input enc_dec_sbox;
  input [7:0]\info_o[23]_INST_0_i_4_1 ;
  input [7:0]\info_o[23]_INST_0_i_4_2 ;
  input \base_new_pp[4]_i_2__0_1 ;
  input [7:0]\CD[1].col[2][23]_i_3 ;
  input \CD[1].col[2][23]_i_3_0 ;
  input [7:0]\CD[1].col[2][23]_i_3_1 ;
  input \CD[1].col[2][23]_i_3_2 ;
  input isomorphism_return179_out_12;
  input isomorphism_return114_out_13;
  input \base_new_pp_reg[4]_3 ;
  input \base_new_pp_reg[3]_0 ;
  input clk_i;

  wire \CD[0].col_reg[3][16] ;
  wire \CD[0].col_reg[3][17] ;
  wire \CD[0].col_reg[3][18] ;
  wire \CD[0].col_reg[3][19] ;
  wire \CD[0].col_reg[3][20] ;
  wire \CD[0].col_reg[3][21] ;
  wire \CD[0].col_reg[3][22] ;
  wire \CD[0].col_reg[3][23] ;
  wire [7:0]\CD[1].col[2][23]_i_3 ;
  wire \CD[1].col[2][23]_i_3_0 ;
  wire [7:0]\CD[1].col[2][23]_i_3_1 ;
  wire \CD[1].col[2][23]_i_3_2 ;
  wire \CD[2].col_reg[1][16] ;
  wire \CD[2].col_reg[1][17] ;
  wire \CD[2].col_reg[1][18] ;
  wire \CD[2].col_reg[1][19] ;
  wire \CD[2].col_reg[1][20] ;
  wire \CD[2].col_reg[1][21] ;
  wire \CD[2].col_reg[1][22] ;
  wire \CD[2].col_reg[1][23] ;
  wire [7:0]D;
  wire [7:0]\KR[3].key_host_reg[0][23] ;
  wire [7:0]\KR[3].key_reg[0][23] ;
  wire [7:0]\KR[3].key_reg[0][23]_0 ;
  wire \base_new_pp[0]_i_1__0_n_0 ;
  wire \base_new_pp[4]_i_1__0_n_0 ;
  wire \base_new_pp[4]_i_2__0_0 ;
  wire \base_new_pp[4]_i_2__0_1 ;
  wire \base_new_pp_reg[1]_0 ;
  wire [7:0]\base_new_pp_reg[2]_0 ;
  wire \base_new_pp_reg[3]_0 ;
  wire \base_new_pp_reg[4]_0 ;
  wire \base_new_pp_reg[4]_1 ;
  wire \base_new_pp_reg[4]_2 ;
  wire \base_new_pp_reg[4]_3 ;
  wire \base_new_pp_reg[6]_0 ;
  wire \base_new_pp_reg[6]_1 ;
  wire \base_new_pp_reg[6]_2 ;
  wire \base_new_pp_reg_n_0_[0] ;
  wire \base_new_pp_reg_n_0_[1] ;
  wire \base_new_pp_reg_n_0_[4] ;
  wire \base_new_pp_reg_n_0_[5] ;
  wire clk_i;
  wire [13:0]enable_i;
  wire enable_i_0_sn_1;
  wire enc_dec_sbox;
  wire [3:0]gf_inv_8_stage1_return;
  wire gf_inv_8_stage1_return1__0;
  wire gf_inv_8_stage1_return2__0;
  wire gf_inv_8_stage1_return349_in;
  wire gf_inv_8_stage1_return540_out;
  wire gf_inv_8_stage1_return542_out;
  wire gf_inv_8_stage1_return546_out;
  wire gf_inv_8_stage1_return547_out;
  wire [1:0]gf_inv_8_stage2_return013_out;
  wire [1:1]gf_inv_8_stage2_return0__3;
  wire [1:0]gf_muls_20_return__1;
  wire [1:0]gf_muls_scl_20_return;
  wire [1:0]gf_muls_scl_2_return;
  wire [1:0]in111_out;
  wire [1:0]in1__0;
  wire [1:0]in2;
  wire [1:0]in21_in;
  wire \info_o[16]_INST_0_i_6_n_0 ;
  wire \info_o[17]_INST_0_i_6_n_0 ;
  wire \info_o[18]_INST_0_i_6_n_0 ;
  wire \info_o[19]_INST_0_i_6_n_0 ;
  wire \info_o[20]_INST_0_i_6_n_0 ;
  wire \info_o[21]_INST_0_i_6_n_0 ;
  wire \info_o[22]_INST_0_i_6_n_0 ;
  wire [7:0]\info_o[23]_INST_0_i_4_0 ;
  wire [7:0]\info_o[23]_INST_0_i_4_1 ;
  wire [7:0]\info_o[23]_INST_0_i_4_2 ;
  wire \info_o[23]_INST_0_i_6_n_0 ;
  wire isomorphism_return076_out;
  wire isomorphism_return114_out_13;
  wire isomorphism_return179_out_12;
  wire isomorphism_return1__0;
  wire isomorphism_return277_out;
  wire [0:0]key_en;
  wire key_sel_mux;
  wire \out_gf_pp[1]_i_3__0_n_0 ;
  wire \out_gf_pp[1]_i_4__0_n_0 ;
  wire \out_gf_pp[2]_i_2__0_n_0 ;
  wire \out_gf_pp[2]_i_6__0_n_0 ;
  wire \out_gf_pp[2]_i_7__0_n_0 ;
  wire \out_gf_pp[3]_i_2__0_n_0 ;
  wire \out_gf_pp[3]_i_5__0_n_0 ;
  wire \out_gf_pp[3]_i_6__0_n_0 ;
  wire \out_gf_pp[3]_i_7__0_n_0 ;
  wire \out_gf_pp_reg_n_0_[0] ;
  wire \out_gf_pp_reg_n_0_[1] ;
  wire \out_gf_pp_reg_n_0_[2] ;
  wire \out_gf_pp_reg_n_0_[3] ;
  wire p_0_in;
  wire p_0_in2_in;
  wire p_0_in9_in;
  wire p_1_in;
  wire p_1_in10_in;
  wire p_1_in17_in;
  wire p_1_in18_in;
  wire p_1_in7_in;
  wire p_72_in;
  wire [16:16]sbox_out_dec;
  wire [1:0]sbox_out_enc;
  wire \sbox_pp2_reg[16] ;
  wire \sbox_pp2_reg[17] ;
  wire \sbox_pp2_reg[18] ;
  wire \sbox_pp2_reg[19] ;
  wire \sbox_pp2_reg[20] ;
  wire \sbox_pp2_reg[21] ;
  wire \sbox_pp2_reg[22] ;
  wire \sbox_pp2_reg[23] ;
  wire \sbox_pp2_reg[23]_0 ;

  assign enable_i_0_sp_1 = enable_i_0_sn_1;
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \KR[2].key[1][16]_i_3 
       (.I0(p_0_in2_in),
        .I1(gf_inv_8_stage2_return013_out[0]),
        .I2(gf_inv_8_stage2_return0__3),
        .O(\base_new_pp_reg[1]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \KR[2].key[1][17]_i_3 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(p_1_in),
        .I2(p_0_in2_in),
        .O(\base_new_pp_reg[4]_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \KR[2].key[1][18]_i_3 
       (.I0(\base_new_pp_reg[6]_2 ),
        .I1(sbox_out_dec),
        .I2(\base_new_pp_reg[4]_1 ),
        .O(sbox_out_enc[0]));
  LUT3 #(
    .INIT(8'h69)) 
    \KR[2].key[1][19]_i_3 
       (.I0(p_0_in2_in),
        .I1(gf_inv_8_stage2_return013_out[0]),
        .I2(\base_new_pp_reg[6]_0 ),
        .O(sbox_out_enc[1]));
  LUT2 #(
    .INIT(4'h9)) 
    \KR[2].key[1][20]_i_3 
       (.I0(\base_new_pp_reg[6]_1 ),
        .I1(p_1_in),
        .O(\base_new_pp_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h96A59955695A66AA)) 
    \KR[2].key[1][21]_i_3 
       (.I0(gf_muls_scl_20_return[0]),
        .I1(\base_new_pp_reg_n_0_[4] ),
        .I2(gf_muls_20_return__1[0]),
        .I3(gf_muls_20_return__1[1]),
        .I4(\base_new_pp_reg_n_0_[5] ),
        .I5(gf_inv_8_stage2_return013_out[0]),
        .O(\base_new_pp_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h609F9F6060606060)) 
    \KR[2].key[1][21]_i_4 
       (.I0(\base_new_pp_reg_n_0_[5] ),
        .I1(in2[1]),
        .I2(in111_out[1]),
        .I3(\base_new_pp_reg_n_0_[4] ),
        .I4(in2[0]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_20_return[0]));
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT4 #(
    .INIT(16'hBE22)) 
    \KR[2].key[1][21]_i_5 
       (.I0(\out_gf_pp_reg_n_0_[2] ),
        .I1(\out_gf_pp_reg_n_0_[0] ),
        .I2(\out_gf_pp_reg_n_0_[1] ),
        .I3(\out_gf_pp_reg_n_0_[3] ),
        .O(gf_muls_20_return__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT4 #(
    .INIT(16'hDD82)) 
    \KR[2].key[1][21]_i_6 
       (.I0(\out_gf_pp_reg_n_0_[3] ),
        .I1(\out_gf_pp_reg_n_0_[1] ),
        .I2(\out_gf_pp_reg_n_0_[0] ),
        .I3(\out_gf_pp_reg_n_0_[2] ),
        .O(gf_muls_20_return__1[1]));
  LUT6 #(
    .INIT(64'hE4281BD71BD7E428)) 
    \KR[2].key[1][22]_i_3 
       (.I0(in2[0]),
        .I1(in1__0[0]),
        .I2(in1__0[1]),
        .I3(in2[1]),
        .I4(gf_muls_scl_20_return[1]),
        .I5(gf_inv_8_stage2_return013_out[1]),
        .O(\base_new_pp_reg[6]_1 ));
  LUT6 #(
    .INIT(64'h1BD7E428E4281BD7)) 
    \KR[2].key[1][23]_i_3 
       (.I0(in2[0]),
        .I1(in1__0[0]),
        .I2(in1__0[1]),
        .I3(in2[1]),
        .I4(gf_muls_scl_20_return[1]),
        .I5(p_1_in),
        .O(\base_new_pp_reg[6]_2 ));
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT4 #(
    .INIT(16'hB2E2)) 
    \KR[2].key[1][23]_i_4 
       (.I0(\out_gf_pp_reg_n_0_[0] ),
        .I1(\out_gf_pp_reg_n_0_[2] ),
        .I2(\out_gf_pp_reg_n_0_[1] ),
        .I3(\out_gf_pp_reg_n_0_[3] ),
        .O(in1__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT4 #(
    .INIT(16'hE4C6)) 
    \KR[2].key[1][23]_i_5 
       (.I0(\out_gf_pp_reg_n_0_[1] ),
        .I1(\out_gf_pp_reg_n_0_[0] ),
        .I2(\out_gf_pp_reg_n_0_[3] ),
        .I3(\out_gf_pp_reg_n_0_[2] ),
        .O(in1__0[1]));
  LUT6 #(
    .INIT(64'h0FF0666669960000)) 
    \KR[2].key[1][23]_i_6 
       (.I0(in2[1]),
        .I1(\base_new_pp_reg_n_0_[5] ),
        .I2(in2[0]),
        .I3(\base_new_pp_reg_n_0_[4] ),
        .I4(in111_out[1]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_20_return[1]));
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT4 #(
    .INIT(16'h23D6)) 
    \KR[2].key[1][23]_i_7 
       (.I0(\out_gf_pp_reg_n_0_[2] ),
        .I1(\out_gf_pp_reg_n_0_[3] ),
        .I2(\out_gf_pp_reg_n_0_[0] ),
        .I3(\out_gf_pp_reg_n_0_[1] ),
        .O(in111_out[1]));
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT4 #(
    .INIT(16'h6DB0)) 
    \KR[2].key[1][23]_i_8 
       (.I0(\out_gf_pp_reg_n_0_[3] ),
        .I1(\out_gf_pp_reg_n_0_[1] ),
        .I2(\out_gf_pp_reg_n_0_[2] ),
        .I3(\out_gf_pp_reg_n_0_[0] ),
        .O(in111_out[0]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][16]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][23] [0]),
        .I2(enable_i[6]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[1]_0 ),
        .I5(\KR[3].key_reg[0][23]_0 [0]),
        .O(\KR[3].key_host_reg[0][23] [0]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][17]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][23] [1]),
        .I2(enable_i[7]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[4]_0 ),
        .I5(\KR[3].key_reg[0][23]_0 [1]),
        .O(\KR[3].key_host_reg[0][23] [1]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][18]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][23] [2]),
        .I2(enable_i[8]),
        .I3(key_sel_mux),
        .I4(sbox_out_enc[0]),
        .I5(\KR[3].key_reg[0][23]_0 [2]),
        .O(\KR[3].key_host_reg[0][23] [2]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][19]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][23] [3]),
        .I2(enable_i[9]),
        .I3(key_sel_mux),
        .I4(sbox_out_enc[1]),
        .I5(\KR[3].key_reg[0][23]_0 [3]),
        .O(\KR[3].key_host_reg[0][23] [3]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][20]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][23] [4]),
        .I2(enable_i[10]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[6]_0 ),
        .I5(\KR[3].key_reg[0][23]_0 [4]),
        .O(\KR[3].key_host_reg[0][23] [4]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][21]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][23] [5]),
        .I2(enable_i[11]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[4]_1 ),
        .I5(\KR[3].key_reg[0][23]_0 [5]),
        .O(\KR[3].key_host_reg[0][23] [5]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][22]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][23] [6]),
        .I2(enable_i[12]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[6]_1 ),
        .I5(\KR[3].key_reg[0][23]_0 [6]),
        .O(\KR[3].key_host_reg[0][23] [6]));
  LUT6 #(
    .INIT(64'hFFE400E400E4FFE4)) 
    \KR[3].key[0][23]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][23] [7]),
        .I2(enable_i[13]),
        .I3(key_sel_mux),
        .I4(\base_new_pp_reg[6]_2 ),
        .I5(\KR[3].key_reg[0][23]_0 [7]),
        .O(\KR[3].key_host_reg[0][23] [7]));
  LUT5 #(
    .INIT(32'h66F0660F)) 
    \base_new_pp[0]_i_1__0 
       (.I0(\CD[0].col_reg[3][18] ),
        .I1(isomorphism_return1__0),
        .I2(\CD[0].col_reg[3][17] ),
        .I3(enc_dec_sbox),
        .I4(isomorphism_return076_out),
        .O(\base_new_pp[0]_i_1__0_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \base_new_pp[0]_i_2__0 
       (.I0(\CD[0].col_reg[3][17] ),
        .I1(\CD[0].col_reg[3][16] ),
        .I2(\CD[0].col_reg[3][22] ),
        .I3(\CD[0].col_reg[3][19] ),
        .O(isomorphism_return1__0));
  LUT4 #(
    .INIT(16'h9669)) 
    \base_new_pp[0]_i_3__0 
       (.I0(\CD[0].col_reg[3][21] ),
        .I1(\CD[0].col_reg[3][16] ),
        .I2(\CD[0].col_reg[3][22] ),
        .I3(\CD[0].col_reg[3][20] ),
        .O(isomorphism_return076_out));
  LUT6 #(
    .INIT(64'hF00F0FF066996699)) 
    \base_new_pp[1]_i_1__0 
       (.I0(\CD[0].col_reg[3][20] ),
        .I1(\CD[0].col_reg[3][19] ),
        .I2(\CD[0].col_reg[3][22] ),
        .I3(\CD[0].col_reg[3][16] ),
        .I4(\CD[0].col_reg[3][21] ),
        .I5(enc_dec_sbox),
        .O(p_0_in));
  LUT5 #(
    .INIT(32'h8BB8B88B)) 
    \base_new_pp[2]_i_1__0 
       (.I0(\CD[0].col_reg[3][16] ),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][18] ),
        .I3(\CD[0].col_reg[3][21] ),
        .I4(\CD[0].col_reg[3][23] ),
        .O(p_0_in9_in));
  LUT6 #(
    .INIT(64'h1DD1E22EE22E1DD1)) 
    \base_new_pp[3]_i_1__0 
       (.I0(\CD[0].col_reg[3][22] ),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][17] ),
        .I3(p_72_in),
        .I4(\CD[0].col_reg[3][23] ),
        .I5(\CD[0].col_reg[3][20] ),
        .O(p_1_in17_in));
  LUT6 #(
    .INIT(64'h011101110111FEEE)) 
    \base_new_pp[3]_i_2__0 
       (.I0(\CD[2].col_reg[1][16] ),
        .I1(\info_o[16]_INST_0_i_6_n_0 ),
        .I2(\base_new_pp_reg[2]_0 [0]),
        .I3(\base_new_pp_reg[4]_2 ),
        .I4(\CD[2].col_reg[1][19] ),
        .I5(\base_new_pp_reg[3]_0 ),
        .O(p_72_in));
  LUT6 #(
    .INIT(64'hF00F66660FF09999)) 
    \base_new_pp[4]_i_1__0 
       (.I0(\CD[0].col_reg[3][19] ),
        .I1(\CD[0].col_reg[3][17] ),
        .I2(\CD[0].col_reg[3][21] ),
        .I3(\CD[0].col_reg[3][23] ),
        .I4(enc_dec_sbox),
        .I5(isomorphism_return277_out),
        .O(\base_new_pp[4]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h011101110111FEEE)) 
    \base_new_pp[4]_i_2__0 
       (.I0(\CD[2].col_reg[1][16] ),
        .I1(\info_o[16]_INST_0_i_6_n_0 ),
        .I2(\base_new_pp_reg[2]_0 [0]),
        .I3(\base_new_pp_reg[4]_2 ),
        .I4(\CD[2].col_reg[1][22] ),
        .I5(\base_new_pp_reg[4]_3 ),
        .O(isomorphism_return277_out));
  LUT6 #(
    .INIT(64'h69966996FF0000FF)) 
    \base_new_pp[5]_i_1__0 
       (.I0(\CD[0].col_reg[3][17] ),
        .I1(\CD[0].col_reg[3][21] ),
        .I2(\CD[0].col_reg[3][16] ),
        .I3(\CD[0].col_reg[3][22] ),
        .I4(\CD[0].col_reg[3][20] ),
        .I5(enc_dec_sbox),
        .O(p_1_in7_in));
  LUT6 #(
    .INIT(64'h3CC3C33CA55A5AA5)) 
    \base_new_pp[6]_i_1__0 
       (.I0(\CD[0].col_reg[3][17] ),
        .I1(\CD[0].col_reg[3][21] ),
        .I2(\CD[0].col_reg[3][16] ),
        .I3(\CD[0].col_reg[3][22] ),
        .I4(\CD[0].col_reg[3][20] ),
        .I5(enc_dec_sbox),
        .O(p_1_in10_in));
  LUT6 #(
    .INIT(64'h3CC36666C33C6666)) 
    \base_new_pp[7]_i_1__0 
       (.I0(\CD[0].col_reg[3][20] ),
        .I1(\CD[0].col_reg[3][23] ),
        .I2(\CD[0].col_reg[3][21] ),
        .I3(\CD[0].col_reg[3][18] ),
        .I4(enc_dec_sbox),
        .I5(isomorphism_return179_out_12),
        .O(p_1_in18_in));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\base_new_pp[0]_i_1__0_n_0 ),
        .Q(\base_new_pp_reg_n_0_[0] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in),
        .Q(\base_new_pp_reg_n_0_[1] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in9_in),
        .Q(in21_in[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in17_in),
        .Q(in21_in[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\base_new_pp[4]_i_1__0_n_0 ),
        .Q(\base_new_pp_reg_n_0_[4] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in7_in),
        .Q(\base_new_pp_reg_n_0_[5] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in10_in),
        .Q(in2[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in18_in),
        .Q(in2[1]),
        .R(1'b0));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[16]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [0]),
        .I2(\info_o[16]_INST_0_i_6_n_0 ),
        .I3(\CD[2].col_reg[1][16] ),
        .O(\CD[0].col_reg[3][16] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[16]_INST_0_i_6 
       (.I0(\info_o[23]_INST_0_i_4_0 [0]),
        .I1(\base_new_pp[4]_i_2__0_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[23]_INST_0_i_4_1 [0]),
        .I4(\info_o[23]_INST_0_i_4_2 [0]),
        .I5(\base_new_pp[4]_i_2__0_1 ),
        .O(\info_o[16]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[16]_INST_0_i_7 
       (.I0(\CD[1].col[2][23]_i_3 [0]),
        .I1(\CD[1].col[2][23]_i_3_0 ),
        .I2(\CD[1].col[2][23]_i_3_1 [0]),
        .I3(\CD[1].col[2][23]_i_3_2 ),
        .O(\CD[2].col_reg[1][16] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[17]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [1]),
        .I2(\info_o[17]_INST_0_i_6_n_0 ),
        .I3(\CD[2].col_reg[1][17] ),
        .O(\CD[0].col_reg[3][17] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[17]_INST_0_i_6 
       (.I0(\info_o[23]_INST_0_i_4_0 [1]),
        .I1(\base_new_pp[4]_i_2__0_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[23]_INST_0_i_4_1 [1]),
        .I4(\info_o[23]_INST_0_i_4_2 [1]),
        .I5(\base_new_pp[4]_i_2__0_1 ),
        .O(\info_o[17]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[17]_INST_0_i_7 
       (.I0(\CD[1].col[2][23]_i_3 [1]),
        .I1(\CD[1].col[2][23]_i_3_0 ),
        .I2(\CD[1].col[2][23]_i_3_1 [1]),
        .I3(\CD[1].col[2][23]_i_3_2 ),
        .O(\CD[2].col_reg[1][17] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[18]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [2]),
        .I2(\info_o[18]_INST_0_i_6_n_0 ),
        .I3(\CD[2].col_reg[1][18] ),
        .O(\CD[0].col_reg[3][18] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[18]_INST_0_i_6 
       (.I0(\info_o[23]_INST_0_i_4_0 [2]),
        .I1(\base_new_pp[4]_i_2__0_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[23]_INST_0_i_4_1 [2]),
        .I4(\info_o[23]_INST_0_i_4_2 [2]),
        .I5(\base_new_pp[4]_i_2__0_1 ),
        .O(\info_o[18]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[18]_INST_0_i_7 
       (.I0(\CD[1].col[2][23]_i_3 [2]),
        .I1(\CD[1].col[2][23]_i_3_0 ),
        .I2(\CD[1].col[2][23]_i_3_1 [2]),
        .I3(\CD[1].col[2][23]_i_3_2 ),
        .O(\CD[2].col_reg[1][18] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[19]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [3]),
        .I2(\info_o[19]_INST_0_i_6_n_0 ),
        .I3(\CD[2].col_reg[1][19] ),
        .O(\CD[0].col_reg[3][19] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[19]_INST_0_i_6 
       (.I0(\info_o[23]_INST_0_i_4_0 [3]),
        .I1(\base_new_pp[4]_i_2__0_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[23]_INST_0_i_4_1 [3]),
        .I4(\info_o[23]_INST_0_i_4_2 [3]),
        .I5(\base_new_pp[4]_i_2__0_1 ),
        .O(\info_o[19]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[19]_INST_0_i_7 
       (.I0(\CD[1].col[2][23]_i_3 [3]),
        .I1(\CD[1].col[2][23]_i_3_0 ),
        .I2(\CD[1].col[2][23]_i_3_1 [3]),
        .I3(\CD[1].col[2][23]_i_3_2 ),
        .O(\CD[2].col_reg[1][19] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[20]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [4]),
        .I2(\info_o[20]_INST_0_i_6_n_0 ),
        .I3(\CD[2].col_reg[1][20] ),
        .O(\CD[0].col_reg[3][20] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[20]_INST_0_i_6 
       (.I0(\info_o[23]_INST_0_i_4_0 [4]),
        .I1(\base_new_pp[4]_i_2__0_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[23]_INST_0_i_4_1 [4]),
        .I4(\info_o[23]_INST_0_i_4_2 [4]),
        .I5(\base_new_pp[4]_i_2__0_1 ),
        .O(\info_o[20]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[20]_INST_0_i_7 
       (.I0(\CD[1].col[2][23]_i_3 [4]),
        .I1(\CD[1].col[2][23]_i_3_0 ),
        .I2(\CD[1].col[2][23]_i_3_1 [4]),
        .I3(\CD[1].col[2][23]_i_3_2 ),
        .O(\CD[2].col_reg[1][20] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[21]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [5]),
        .I2(\info_o[21]_INST_0_i_6_n_0 ),
        .I3(\CD[2].col_reg[1][21] ),
        .O(\CD[0].col_reg[3][21] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[21]_INST_0_i_6 
       (.I0(\info_o[23]_INST_0_i_4_0 [5]),
        .I1(\base_new_pp[4]_i_2__0_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[23]_INST_0_i_4_1 [5]),
        .I4(\info_o[23]_INST_0_i_4_2 [5]),
        .I5(\base_new_pp[4]_i_2__0_1 ),
        .O(\info_o[21]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[21]_INST_0_i_7 
       (.I0(\CD[1].col[2][23]_i_3 [5]),
        .I1(\CD[1].col[2][23]_i_3_0 ),
        .I2(\CD[1].col[2][23]_i_3_1 [5]),
        .I3(\CD[1].col[2][23]_i_3_2 ),
        .O(\CD[2].col_reg[1][21] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[22]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [6]),
        .I2(\info_o[22]_INST_0_i_6_n_0 ),
        .I3(\CD[2].col_reg[1][22] ),
        .O(\CD[0].col_reg[3][22] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[22]_INST_0_i_6 
       (.I0(\info_o[23]_INST_0_i_4_0 [6]),
        .I1(\base_new_pp[4]_i_2__0_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[23]_INST_0_i_4_1 [6]),
        .I4(\info_o[23]_INST_0_i_4_2 [6]),
        .I5(\base_new_pp[4]_i_2__0_1 ),
        .O(\info_o[22]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[22]_INST_0_i_7 
       (.I0(\CD[1].col[2][23]_i_3 [6]),
        .I1(\CD[1].col[2][23]_i_3_0 ),
        .I2(\CD[1].col[2][23]_i_3_1 [6]),
        .I3(\CD[1].col[2][23]_i_3_2 ),
        .O(\CD[2].col_reg[1][22] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[23]_INST_0_i_4 
       (.I0(\base_new_pp_reg[4]_2 ),
        .I1(\base_new_pp_reg[2]_0 [7]),
        .I2(\info_o[23]_INST_0_i_6_n_0 ),
        .I3(\CD[2].col_reg[1][23] ),
        .O(\CD[0].col_reg[3][23] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[23]_INST_0_i_6 
       (.I0(\info_o[23]_INST_0_i_4_0 [7]),
        .I1(\base_new_pp[4]_i_2__0_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[23]_INST_0_i_4_1 [7]),
        .I4(\info_o[23]_INST_0_i_4_2 [7]),
        .I5(\base_new_pp[4]_i_2__0_1 ),
        .O(\info_o[23]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[23]_INST_0_i_7 
       (.I0(\CD[1].col[2][23]_i_3 [7]),
        .I1(\CD[1].col[2][23]_i_3_0 ),
        .I2(\CD[1].col[2][23]_i_3_1 [7]),
        .I3(\CD[1].col[2][23]_i_3_2 ),
        .O(\CD[2].col_reg[1][23] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF7FFFF)) 
    \info_o[31]_INST_0_i_7 
       (.I0(enable_i[0]),
        .I1(enable_i[5]),
        .I2(enable_i[4]),
        .I3(enable_i[3]),
        .I4(enable_i[1]),
        .I5(enable_i[2]),
        .O(enable_i_0_sn_1));
  LUT6 #(
    .INIT(64'hA9A69A955659656A)) 
    \out_gf_pp[0]_i_1__0 
       (.I0(gf_inv_8_stage1_return2__0),
        .I1(p_1_in7_in),
        .I2(p_0_in),
        .I3(\base_new_pp[4]_i_1__0_n_0 ),
        .I4(\base_new_pp[0]_i_1__0_n_0 ),
        .I5(gf_inv_8_stage1_return1__0),
        .O(gf_inv_8_stage1_return[0]));
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT4 #(
    .INIT(16'hF99F)) 
    \out_gf_pp[0]_i_2__0 
       (.I0(p_1_in18_in),
        .I1(p_1_in7_in),
        .I2(p_1_in17_in),
        .I3(p_0_in),
        .O(gf_inv_8_stage1_return2__0));
  LUT6 #(
    .INIT(64'h9999969699666996)) 
    \out_gf_pp[1]_i_1__0 
       (.I0(gf_inv_8_stage1_return1__0),
        .I1(gf_inv_8_stage1_return349_in),
        .I2(\out_gf_pp[1]_i_3__0_n_0 ),
        .I3(\out_gf_pp[3]_i_5__0_n_0 ),
        .I4(\out_gf_pp[3]_i_6__0_n_0 ),
        .I5(\out_gf_pp[1]_i_4__0_n_0 ),
        .O(gf_inv_8_stage1_return[1]));
  LUT6 #(
    .INIT(64'hF5C5FFCFFFCFFACA)) 
    \out_gf_pp[1]_i_2__0 
       (.I0(\CD[0].col_reg[3][22] ),
        .I1(\CD[0].col_reg[3][17] ),
        .I2(enc_dec_sbox),
        .I3(isomorphism_return114_out_13),
        .I4(p_72_in),
        .I5(\CD[0].col_reg[3][20] ),
        .O(gf_inv_8_stage1_return349_in));
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[1]_i_3__0 
       (.I0(\base_new_pp[4]_i_1__0_n_0 ),
        .I1(p_1_in7_in),
        .O(\out_gf_pp[1]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[1]_i_4__0 
       (.I0(p_1_in18_in),
        .I1(p_1_in10_in),
        .O(\out_gf_pp[1]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h6A6A6A959595956A)) 
    \out_gf_pp[2]_i_1__0 
       (.I0(\out_gf_pp[2]_i_2__0_n_0 ),
        .I1(p_1_in10_in),
        .I2(p_0_in9_in),
        .I3(gf_inv_8_stage1_return542_out),
        .I4(gf_inv_8_stage1_return540_out),
        .I5(gf_inv_8_stage1_return1__0),
        .O(gf_inv_8_stage1_return[2]));
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT4 #(
    .INIT(16'hF99F)) 
    \out_gf_pp[2]_i_2__0 
       (.I0(p_0_in9_in),
        .I1(p_1_in17_in),
        .I2(p_1_in10_in),
        .I3(p_1_in18_in),
        .O(\out_gf_pp[2]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[2]_i_3__0 
       (.I0(p_1_in7_in),
        .I1(p_1_in18_in),
        .O(gf_inv_8_stage1_return542_out));
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[2]_i_4__0 
       (.I0(p_0_in),
        .I1(p_1_in17_in),
        .O(gf_inv_8_stage1_return540_out));
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT5 #(
    .INIT(32'hF9F9F99F)) 
    \out_gf_pp[2]_i_5__0 
       (.I0(p_1_in10_in),
        .I1(\base_new_pp[4]_i_1__0_n_0 ),
        .I2(p_0_in9_in),
        .I3(\out_gf_pp[2]_i_6__0_n_0 ),
        .I4(\out_gf_pp[2]_i_7__0_n_0 ),
        .O(gf_inv_8_stage1_return1__0));
  LUT6 #(
    .INIT(64'h9669000069960000)) 
    \out_gf_pp[2]_i_6__0 
       (.I0(\CD[0].col_reg[3][17] ),
        .I1(\CD[0].col_reg[3][16] ),
        .I2(\CD[0].col_reg[3][22] ),
        .I3(\CD[0].col_reg[3][19] ),
        .I4(enc_dec_sbox),
        .I5(\CD[0].col_reg[3][18] ),
        .O(\out_gf_pp[2]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000966900006996)) 
    \out_gf_pp[2]_i_7__0 
       (.I0(\CD[0].col_reg[3][21] ),
        .I1(\CD[0].col_reg[3][16] ),
        .I2(\CD[0].col_reg[3][22] ),
        .I3(\CD[0].col_reg[3][20] ),
        .I4(enc_dec_sbox),
        .I5(\CD[0].col_reg[3][17] ),
        .O(\out_gf_pp[2]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h5656565656A9A956)) 
    \out_gf_pp[3]_i_1__0 
       (.I0(\out_gf_pp[3]_i_2__0_n_0 ),
        .I1(gf_inv_8_stage1_return547_out),
        .I2(gf_inv_8_stage1_return546_out),
        .I3(\out_gf_pp[3]_i_5__0_n_0 ),
        .I4(\out_gf_pp[3]_i_6__0_n_0 ),
        .I5(\out_gf_pp[3]_i_7__0_n_0 ),
        .O(gf_inv_8_stage1_return[3]));
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT4 #(
    .INIT(16'hA6C0)) 
    \out_gf_pp[3]_i_2__0 
       (.I0(p_1_in18_in),
        .I1(p_1_in10_in),
        .I2(p_1_in17_in),
        .I3(p_0_in9_in),
        .O(\out_gf_pp[3]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[3]_i_3__0 
       (.I0(\base_new_pp[4]_i_1__0_n_0 ),
        .I1(p_1_in10_in),
        .O(gf_inv_8_stage1_return547_out));
  LUT6 #(
    .INIT(64'hDE1212DE21EDED21)) 
    \out_gf_pp[3]_i_4__0 
       (.I0(isomorphism_return076_out),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][17] ),
        .I3(isomorphism_return1__0),
        .I4(\CD[0].col_reg[3][18] ),
        .I5(p_0_in9_in),
        .O(gf_inv_8_stage1_return546_out));
  LUT6 #(
    .INIT(64'hDE1212DE21EDED21)) 
    \out_gf_pp[3]_i_5__0 
       (.I0(isomorphism_return076_out),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][17] ),
        .I3(isomorphism_return1__0),
        .I4(\CD[0].col_reg[3][18] ),
        .I5(p_0_in),
        .O(\out_gf_pp[3]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[3]_i_6__0 
       (.I0(p_1_in17_in),
        .I1(p_0_in9_in),
        .O(\out_gf_pp[3]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \out_gf_pp[3]_i_7__0 
       (.I0(p_1_in10_in),
        .I1(p_1_in18_in),
        .I2(p_1_in7_in),
        .I3(\base_new_pp[4]_i_1__0_n_0 ),
        .O(\out_gf_pp[3]_i_7__0_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[0]),
        .Q(\out_gf_pp_reg_n_0_[0] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[1]),
        .Q(\out_gf_pp_reg_n_0_[1] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[2]),
        .Q(\out_gf_pp_reg_n_0_[2] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[3]),
        .Q(\out_gf_pp_reg_n_0_[3] ),
        .R(1'b0));
  LUT4 #(
    .INIT(16'h0F66)) 
    \sbox_pp2[16]_i_1 
       (.I0(sbox_out_dec),
        .I1(\sbox_pp2_reg[16] ),
        .I2(\base_new_pp_reg[1]_0 ),
        .I3(\sbox_pp2_reg[23] ),
        .O(D[0]));
  LUT5 #(
    .INIT(32'h00FF9696)) 
    \sbox_pp2[17]_i_1 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(p_1_in),
        .I2(\sbox_pp2_reg[17] ),
        .I3(\base_new_pp_reg[4]_0 ),
        .I4(\sbox_pp2_reg[23] ),
        .O(D[1]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[17]_i_2 
       (.I0(\base_new_pp_reg_n_0_[0] ),
        .I1(gf_muls_20_return__1[0]),
        .I2(gf_muls_20_return__1[1]),
        .I3(\base_new_pp_reg_n_0_[1] ),
        .I4(gf_muls_scl_2_return[1]),
        .O(p_1_in));
  LUT5 #(
    .INIT(32'hFF960096)) 
    \sbox_pp2[18]_i_1 
       (.I0(\base_new_pp_reg[4]_0 ),
        .I1(gf_inv_8_stage2_return013_out[1]),
        .I2(\sbox_pp2_reg[18] ),
        .I3(\sbox_pp2_reg[23] ),
        .I4(sbox_out_enc[0]),
        .O(D[2]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[18]_i_2 
       (.I0(in21_in[0]),
        .I1(in1__0[0]),
        .I2(in1__0[1]),
        .I3(in21_in[1]),
        .I4(gf_muls_scl_2_return[1]),
        .O(gf_inv_8_stage2_return013_out[1]));
  LUT6 #(
    .INIT(64'h0FF0666669960000)) 
    \sbox_pp2[18]_i_3 
       (.I0(in21_in[1]),
        .I1(\base_new_pp_reg_n_0_[1] ),
        .I2(in21_in[0]),
        .I3(\base_new_pp_reg_n_0_[0] ),
        .I4(in111_out[1]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_2_return[1]));
  LUT6 #(
    .INIT(64'hFFFF966900009669)) 
    \sbox_pp2[19]_i_1 
       (.I0(\base_new_pp_reg[6]_2 ),
        .I1(sbox_out_dec),
        .I2(\base_new_pp_reg[1]_0 ),
        .I3(\sbox_pp2_reg[19] ),
        .I4(\sbox_pp2_reg[23] ),
        .I5(sbox_out_enc[1]),
        .O(D[3]));
  LUT5 #(
    .INIT(32'h00FF9696)) 
    \sbox_pp2[20]_i_1 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(gf_inv_8_stage2_return013_out[0]),
        .I2(\sbox_pp2_reg[20] ),
        .I3(\base_new_pp_reg[6]_0 ),
        .I4(\sbox_pp2_reg[23] ),
        .O(D[4]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[20]_i_2 
       (.I0(in21_in[1]),
        .I1(in1__0[1]),
        .I2(in1__0[0]),
        .I3(in21_in[0]),
        .I4(gf_muls_scl_2_return[0]),
        .O(gf_inv_8_stage2_return013_out[0]));
  LUT5 #(
    .INIT(32'h00FF9669)) 
    \sbox_pp2[21]_i_1 
       (.I0(\base_new_pp_reg[6]_0 ),
        .I1(sbox_out_dec),
        .I2(\sbox_pp2_reg[21] ),
        .I3(\base_new_pp_reg[4]_1 ),
        .I4(\sbox_pp2_reg[23] ),
        .O(D[5]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[21]_i_2 
       (.I0(in2[1]),
        .I1(in1__0[1]),
        .I2(in1__0[0]),
        .I3(in2[0]),
        .I4(gf_muls_scl_20_return[0]),
        .O(sbox_out_dec));
  LUT6 #(
    .INIT(64'h0000FFFF96699669)) 
    \sbox_pp2[22]_i_1 
       (.I0(\base_new_pp_reg[6]_0 ),
        .I1(\base_new_pp_reg[4]_1 ),
        .I2(gf_inv_8_stage2_return0__3),
        .I3(\sbox_pp2_reg[22] ),
        .I4(\base_new_pp_reg[6]_1 ),
        .I5(\sbox_pp2_reg[23] ),
        .O(D[6]));
  LUT5 #(
    .INIT(32'h00FF9696)) 
    \sbox_pp2[23]_i_1 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(p_0_in2_in),
        .I2(\sbox_pp2_reg[23]_0 ),
        .I3(\base_new_pp_reg[6]_2 ),
        .I4(\sbox_pp2_reg[23] ),
        .O(D[7]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[23]_i_2 
       (.I0(\base_new_pp_reg_n_0_[4] ),
        .I1(gf_muls_20_return__1[0]),
        .I2(gf_muls_20_return__1[1]),
        .I3(\base_new_pp_reg_n_0_[5] ),
        .I4(gf_muls_scl_20_return[1]),
        .O(gf_inv_8_stage2_return0__3));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[23]_i_3 
       (.I0(\base_new_pp_reg_n_0_[1] ),
        .I1(gf_muls_20_return__1[1]),
        .I2(gf_muls_20_return__1[0]),
        .I3(\base_new_pp_reg_n_0_[0] ),
        .I4(gf_muls_scl_2_return[0]),
        .O(p_0_in2_in));
  LUT6 #(
    .INIT(64'h609F9F6060606060)) 
    \sbox_pp2[23]_i_4 
       (.I0(\base_new_pp_reg_n_0_[1] ),
        .I1(in21_in[1]),
        .I2(in111_out[1]),
        .I3(\base_new_pp_reg_n_0_[0] ),
        .I4(in21_in[0]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_2_return[0]));
endmodule

(* ORIG_REF_NAME = "sBox_8" *) 
module switch_elements_sBox_8_3
   (\round_pp1_reg[0] ,
    \round_pp1_reg[3] ,
    \round_pp1_reg[3]_0 ,
    \round_pp1_reg[0]_0 ,
    \round_pp1_reg[3]_1 ,
    D,
    \round_pp1_reg[0]_1 ,
    \KR[3].key_host_reg[0][31] ,
    g_func,
    \CD[0].col_reg[3][31] ,
    \CD[2].col_reg[1][31] ,
    \CD[0].col_reg[3][30] ,
    \CD[2].col_reg[1][30] ,
    \CD[0].col_reg[3][29] ,
    \CD[2].col_reg[1][29] ,
    \CD[0].col_reg[3][28] ,
    \CD[2].col_reg[1][28] ,
    \CD[0].col_reg[3][27] ,
    \CD[2].col_reg[1][27] ,
    \CD[0].col_reg[3][26] ,
    \CD[2].col_reg[1][26] ,
    \CD[0].col_reg[3][25] ,
    \CD[2].col_reg[1][25] ,
    \CD[0].col_reg[3][24] ,
    \CD[2].col_reg[1][24] ,
    Q,
    enc_dec_sbox,
    \sbox_pp2_reg[30] ,
    \sbox_pp2_reg[31] ,
    \sbox_pp2_reg[26] ,
    \sbox_pp2_reg[28] ,
    \sbox_pp2_reg[27] ,
    \sbox_pp2_reg[24] ,
    \sbox_pp2_reg[25] ,
    \sbox_pp2_reg[31]_0 ,
    key_en,
    \KR[3].key_reg[0][31] ,
    enable_i,
    key_sel_mux,
    \KR[3].key_reg[0][31]_0 ,
    \sbox_pp2_reg[29] ,
    \base_new_pp_reg[4]_0 ,
    \base_new_pp_reg[2]_0 ,
    \info_o[31]_INST_0_i_9_0 ,
    \base_new_pp[4]_i_2_0 ,
    \info_o[31]_INST_0_i_9_1 ,
    \info_o[31]_INST_0_i_9_2 ,
    \base_new_pp[4]_i_2_1 ,
    \CD[0].col[3][31]_i_14 ,
    \CD[0].col[3][31]_i_14_0 ,
    \CD[0].col[3][31]_i_14_1 ,
    \CD[0].col[3][31]_i_14_2 ,
    rc,
    isomorphism_return179_out,
    isomorphism_return114_out,
    \base_new_pp_reg[4]_1 ,
    \base_new_pp_reg[3]_0 ,
    clk_i);
  output \round_pp1_reg[0] ;
  output \round_pp1_reg[3] ;
  output \round_pp1_reg[3]_0 ;
  output \round_pp1_reg[0]_0 ;
  output \round_pp1_reg[3]_1 ;
  output [7:0]D;
  output \round_pp1_reg[0]_1 ;
  output [7:0]\KR[3].key_host_reg[0][31] ;
  output [1:0]g_func;
  output \CD[0].col_reg[3][31] ;
  output \CD[2].col_reg[1][31] ;
  output \CD[0].col_reg[3][30] ;
  output \CD[2].col_reg[1][30] ;
  output \CD[0].col_reg[3][29] ;
  output \CD[2].col_reg[1][29] ;
  output \CD[0].col_reg[3][28] ;
  output \CD[2].col_reg[1][28] ;
  output \CD[0].col_reg[3][27] ;
  output \CD[2].col_reg[1][27] ;
  output \CD[0].col_reg[3][26] ;
  output \CD[2].col_reg[1][26] ;
  output \CD[0].col_reg[3][25] ;
  output \CD[2].col_reg[1][25] ;
  output \CD[0].col_reg[3][24] ;
  output \CD[2].col_reg[1][24] ;
  input [3:0]Q;
  input enc_dec_sbox;
  input \sbox_pp2_reg[30] ;
  input \sbox_pp2_reg[31] ;
  input \sbox_pp2_reg[26] ;
  input \sbox_pp2_reg[28] ;
  input \sbox_pp2_reg[27] ;
  input \sbox_pp2_reg[24] ;
  input \sbox_pp2_reg[25] ;
  input \sbox_pp2_reg[31]_0 ;
  input [0:0]key_en;
  input [7:0]\KR[3].key_reg[0][31] ;
  input [7:0]enable_i;
  input key_sel_mux;
  input [7:0]\KR[3].key_reg[0][31]_0 ;
  input \sbox_pp2_reg[29] ;
  input \base_new_pp_reg[4]_0 ;
  input [7:0]\base_new_pp_reg[2]_0 ;
  input [7:0]\info_o[31]_INST_0_i_9_0 ;
  input \base_new_pp[4]_i_2_0 ;
  input [7:0]\info_o[31]_INST_0_i_9_1 ;
  input [7:0]\info_o[31]_INST_0_i_9_2 ;
  input \base_new_pp[4]_i_2_1 ;
  input [7:0]\CD[0].col[3][31]_i_14 ;
  input \CD[0].col[3][31]_i_14_0 ;
  input [7:0]\CD[0].col[3][31]_i_14_1 ;
  input \CD[0].col[3][31]_i_14_2 ;
  input [1:0]rc;
  input isomorphism_return179_out;
  input isomorphism_return114_out;
  input \base_new_pp_reg[4]_1 ;
  input \base_new_pp_reg[3]_0 ;
  input clk_i;

  wire [7:0]\CD[0].col[3][31]_i_14 ;
  wire \CD[0].col[3][31]_i_14_0 ;
  wire [7:0]\CD[0].col[3][31]_i_14_1 ;
  wire \CD[0].col[3][31]_i_14_2 ;
  wire \CD[0].col_reg[3][24] ;
  wire \CD[0].col_reg[3][25] ;
  wire \CD[0].col_reg[3][26] ;
  wire \CD[0].col_reg[3][27] ;
  wire \CD[0].col_reg[3][28] ;
  wire \CD[0].col_reg[3][29] ;
  wire \CD[0].col_reg[3][30] ;
  wire \CD[0].col_reg[3][31] ;
  wire \CD[2].col_reg[1][24] ;
  wire \CD[2].col_reg[1][25] ;
  wire \CD[2].col_reg[1][26] ;
  wire \CD[2].col_reg[1][27] ;
  wire \CD[2].col_reg[1][28] ;
  wire \CD[2].col_reg[1][29] ;
  wire \CD[2].col_reg[1][30] ;
  wire \CD[2].col_reg[1][31] ;
  wire [7:0]D;
  wire [7:0]\KR[3].key_host_reg[0][31] ;
  wire [7:0]\KR[3].key_reg[0][31] ;
  wire [7:0]\KR[3].key_reg[0][31]_0 ;
  wire [3:0]Q;
  wire \base_new_pp[0]_i_1_n_0 ;
  wire \base_new_pp[4]_i_1_n_0 ;
  wire \base_new_pp[4]_i_2_0 ;
  wire \base_new_pp[4]_i_2_1 ;
  wire [7:0]\base_new_pp_reg[2]_0 ;
  wire \base_new_pp_reg[3]_0 ;
  wire \base_new_pp_reg[4]_0 ;
  wire \base_new_pp_reg[4]_1 ;
  wire \base_new_pp_reg_n_0_[0] ;
  wire \base_new_pp_reg_n_0_[1] ;
  wire \base_new_pp_reg_n_0_[4] ;
  wire \base_new_pp_reg_n_0_[5] ;
  wire clk_i;
  wire [7:0]enable_i;
  wire enc_dec_sbox;
  wire [1:0]g_func;
  wire [3:0]gf_inv_8_stage1_return;
  wire gf_inv_8_stage1_return1__0;
  wire gf_inv_8_stage1_return2__0;
  wire gf_inv_8_stage1_return349_in;
  wire gf_inv_8_stage1_return540_out;
  wire gf_inv_8_stage1_return542_out;
  wire gf_inv_8_stage1_return546_out;
  wire gf_inv_8_stage1_return547_out;
  wire [1:0]gf_inv_8_stage2_return013_out;
  wire [1:1]gf_inv_8_stage2_return0__3;
  wire [1:0]gf_muls_20_return__1;
  wire [1:0]gf_muls_scl_20_return;
  wire [1:0]gf_muls_scl_2_return;
  wire [1:0]in111_out;
  wire [1:0]in1__0;
  wire [1:0]in2;
  wire [1:0]in21_in;
  wire \info_o[24]_INST_0_i_9_n_0 ;
  wire \info_o[25]_INST_0_i_9_n_0 ;
  wire \info_o[26]_INST_0_i_9_n_0 ;
  wire \info_o[27]_INST_0_i_9_n_0 ;
  wire \info_o[28]_INST_0_i_11_n_0 ;
  wire \info_o[29]_INST_0_i_11_n_0 ;
  wire \info_o[30]_INST_0_i_11_n_0 ;
  wire \info_o[31]_INST_0_i_20_n_0 ;
  wire [7:0]\info_o[31]_INST_0_i_9_0 ;
  wire [7:0]\info_o[31]_INST_0_i_9_1 ;
  wire [7:0]\info_o[31]_INST_0_i_9_2 ;
  wire isomorphism_inv_return033_out;
  wire isomorphism_inv_return03_out;
  wire isomorphism_inv_return05_out;
  wire isomorphism_return076_out;
  wire isomorphism_return114_out;
  wire isomorphism_return179_out;
  wire isomorphism_return1__0;
  wire isomorphism_return277_out;
  wire [0:0]key_en;
  wire key_sel_mux;
  wire \out_gf_pp[1]_i_3_n_0 ;
  wire \out_gf_pp[1]_i_4_n_0 ;
  wire \out_gf_pp[2]_i_2_n_0 ;
  wire \out_gf_pp[2]_i_6_n_0 ;
  wire \out_gf_pp[2]_i_7_n_0 ;
  wire \out_gf_pp[3]_i_2_n_0 ;
  wire \out_gf_pp[3]_i_5_n_0 ;
  wire \out_gf_pp[3]_i_6_n_0 ;
  wire \out_gf_pp[3]_i_7_n_0 ;
  wire \out_gf_pp_reg_n_0_[0] ;
  wire \out_gf_pp_reg_n_0_[1] ;
  wire \out_gf_pp_reg_n_0_[2] ;
  wire \out_gf_pp_reg_n_0_[3] ;
  wire p_0_in;
  wire p_0_in2_in;
  wire p_0_in9_in;
  wire p_16_in;
  wire p_1_in;
  wire p_1_in10_in;
  wire p_1_in17_in;
  wire p_1_in18_in;
  wire p_1_in7_in;
  wire p_72_in;
  wire p_92_in;
  wire p_93_in;
  wire p_95_in;
  wire [1:0]rc;
  wire \round_pp1_reg[0] ;
  wire \round_pp1_reg[0]_0 ;
  wire \round_pp1_reg[0]_1 ;
  wire \round_pp1_reg[3] ;
  wire \round_pp1_reg[3]_0 ;
  wire \round_pp1_reg[3]_1 ;
  wire [24:24]sbox_out_dec;
  wire \sbox_pp2_reg[24] ;
  wire \sbox_pp2_reg[25] ;
  wire \sbox_pp2_reg[26] ;
  wire \sbox_pp2_reg[27] ;
  wire \sbox_pp2_reg[28] ;
  wire \sbox_pp2_reg[29] ;
  wire \sbox_pp2_reg[30] ;
  wire \sbox_pp2_reg[31] ;
  wire \sbox_pp2_reg[31]_0 ;

  LUT6 #(
    .INIT(64'h9999999699999969)) 
    \KR[2].key[1][24]_i_3 
       (.I0(p_95_in),
        .I1(gf_inv_8_stage2_return0__3),
        .I2(Q[0]),
        .I3(Q[2]),
        .I4(Q[1]),
        .I5(enc_dec_sbox),
        .O(\round_pp1_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h03020103FCFDFEFC)) 
    \KR[2].key[1][25]_i_3 
       (.I0(Q[3]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(Q[0]),
        .I4(enc_dec_sbox),
        .I5(p_16_in),
        .O(\round_pp1_reg[3]_1 ));
  LUT3 #(
    .INIT(8'h69)) 
    \KR[2].key[1][26]_i_3 
       (.I0(rc[0]),
        .I1(p_93_in),
        .I2(p_92_in),
        .O(g_func[0]));
  LUT3 #(
    .INIT(8'h69)) 
    \KR[2].key[1][27]_i_3 
       (.I0(rc[1]),
        .I1(p_95_in),
        .I2(isomorphism_inv_return03_out),
        .O(g_func[1]));
  LUT6 #(
    .INIT(64'h02121101FDEDEEFE)) 
    \KR[2].key[1][28]_i_3 
       (.I0(Q[3]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(Q[0]),
        .I4(enc_dec_sbox),
        .I5(isomorphism_inv_return03_out),
        .O(\round_pp1_reg[3] ));
  LUT6 #(
    .INIT(64'h02080005FDF7FFFA)) 
    \KR[2].key[1][29]_i_3 
       (.I0(Q[0]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[3]),
        .I4(enc_dec_sbox),
        .I5(p_93_in),
        .O(\round_pp1_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h10000200EFFFFDFF)) 
    \KR[2].key[1][30]_i_3 
       (.I0(Q[0]),
        .I1(Q[3]),
        .I2(Q[2]),
        .I3(Q[1]),
        .I4(enc_dec_sbox),
        .I5(isomorphism_inv_return033_out),
        .O(\round_pp1_reg[0] ));
  LUT6 #(
    .INIT(64'h40000100BFFFFEFF)) 
    \KR[2].key[1][31]_i_4 
       (.I0(Q[3]),
        .I1(Q[0]),
        .I2(Q[2]),
        .I3(Q[1]),
        .I4(enc_dec_sbox),
        .I5(isomorphism_inv_return05_out),
        .O(\round_pp1_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][24]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][31] [0]),
        .I2(enable_i[0]),
        .I3(key_sel_mux),
        .I4(\round_pp1_reg[0]_1 ),
        .I5(\KR[3].key_reg[0][31]_0 [0]),
        .O(\KR[3].key_host_reg[0][31] [0]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][25]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][31] [1]),
        .I2(enable_i[1]),
        .I3(key_sel_mux),
        .I4(\round_pp1_reg[3]_1 ),
        .I5(\KR[3].key_reg[0][31]_0 [1]),
        .O(\KR[3].key_host_reg[0][31] [1]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][26]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][31] [2]),
        .I2(enable_i[2]),
        .I3(key_sel_mux),
        .I4(g_func[0]),
        .I5(\KR[3].key_reg[0][31]_0 [2]),
        .O(\KR[3].key_host_reg[0][31] [2]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][27]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][31] [3]),
        .I2(enable_i[3]),
        .I3(key_sel_mux),
        .I4(g_func[1]),
        .I5(\KR[3].key_reg[0][31]_0 [3]),
        .O(\KR[3].key_host_reg[0][31] [3]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][28]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][31] [4]),
        .I2(enable_i[4]),
        .I3(key_sel_mux),
        .I4(\round_pp1_reg[3] ),
        .I5(\KR[3].key_reg[0][31]_0 [4]),
        .O(\KR[3].key_host_reg[0][31] [4]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][29]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][31] [5]),
        .I2(enable_i[5]),
        .I3(key_sel_mux),
        .I4(\round_pp1_reg[0]_0 ),
        .I5(\KR[3].key_reg[0][31]_0 [5]),
        .O(\KR[3].key_host_reg[0][31] [5]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][30]_i_1 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][31] [6]),
        .I2(enable_i[6]),
        .I3(key_sel_mux),
        .I4(\round_pp1_reg[0] ),
        .I5(\KR[3].key_reg[0][31]_0 [6]),
        .O(\KR[3].key_host_reg[0][31] [6]));
  LUT6 #(
    .INIT(64'h00E4FFE4FFE400E4)) 
    \KR[3].key[0][31]_i_2 
       (.I0(key_en),
        .I1(\KR[3].key_reg[0][31] [7]),
        .I2(enable_i[7]),
        .I3(key_sel_mux),
        .I4(\round_pp1_reg[3]_0 ),
        .I5(\KR[3].key_reg[0][31]_0 [7]),
        .O(\KR[3].key_host_reg[0][31] [7]));
  LUT5 #(
    .INIT(32'h66F0660F)) 
    \base_new_pp[0]_i_1 
       (.I0(\CD[0].col_reg[3][26] ),
        .I1(isomorphism_return1__0),
        .I2(\CD[0].col_reg[3][25] ),
        .I3(enc_dec_sbox),
        .I4(isomorphism_return076_out),
        .O(\base_new_pp[0]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h6996)) 
    \base_new_pp[0]_i_2 
       (.I0(\CD[0].col_reg[3][25] ),
        .I1(\CD[0].col_reg[3][24] ),
        .I2(\CD[0].col_reg[3][30] ),
        .I3(\CD[0].col_reg[3][27] ),
        .O(isomorphism_return1__0));
  LUT4 #(
    .INIT(16'h9669)) 
    \base_new_pp[0]_i_3 
       (.I0(\CD[0].col_reg[3][29] ),
        .I1(\CD[0].col_reg[3][24] ),
        .I2(\CD[0].col_reg[3][30] ),
        .I3(\CD[0].col_reg[3][28] ),
        .O(isomorphism_return076_out));
  LUT6 #(
    .INIT(64'hF00F0FF066996699)) 
    \base_new_pp[1]_i_1 
       (.I0(\CD[0].col_reg[3][28] ),
        .I1(\CD[0].col_reg[3][27] ),
        .I2(\CD[0].col_reg[3][30] ),
        .I3(\CD[0].col_reg[3][24] ),
        .I4(\CD[0].col_reg[3][29] ),
        .I5(enc_dec_sbox),
        .O(p_0_in));
  LUT5 #(
    .INIT(32'h8BB8B88B)) 
    \base_new_pp[2]_i_1 
       (.I0(\CD[0].col_reg[3][24] ),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][26] ),
        .I3(\CD[0].col_reg[3][29] ),
        .I4(\CD[0].col_reg[3][31] ),
        .O(p_0_in9_in));
  LUT6 #(
    .INIT(64'h1DD1E22EE22E1DD1)) 
    \base_new_pp[3]_i_1 
       (.I0(\CD[0].col_reg[3][30] ),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][25] ),
        .I3(p_72_in),
        .I4(\CD[0].col_reg[3][31] ),
        .I5(\CD[0].col_reg[3][28] ),
        .O(p_1_in17_in));
  LUT6 #(
    .INIT(64'h011101110111FEEE)) 
    \base_new_pp[3]_i_2 
       (.I0(\CD[2].col_reg[1][24] ),
        .I1(\info_o[24]_INST_0_i_9_n_0 ),
        .I2(\base_new_pp_reg[2]_0 [0]),
        .I3(\base_new_pp_reg[4]_0 ),
        .I4(\CD[2].col_reg[1][27] ),
        .I5(\base_new_pp_reg[3]_0 ),
        .O(p_72_in));
  LUT6 #(
    .INIT(64'hF00F66660FF09999)) 
    \base_new_pp[4]_i_1 
       (.I0(\CD[0].col_reg[3][27] ),
        .I1(\CD[0].col_reg[3][25] ),
        .I2(\CD[0].col_reg[3][29] ),
        .I3(\CD[0].col_reg[3][31] ),
        .I4(enc_dec_sbox),
        .I5(isomorphism_return277_out),
        .O(\base_new_pp[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h011101110111FEEE)) 
    \base_new_pp[4]_i_2 
       (.I0(\CD[2].col_reg[1][24] ),
        .I1(\info_o[24]_INST_0_i_9_n_0 ),
        .I2(\base_new_pp_reg[2]_0 [0]),
        .I3(\base_new_pp_reg[4]_0 ),
        .I4(\CD[2].col_reg[1][30] ),
        .I5(\base_new_pp_reg[4]_1 ),
        .O(isomorphism_return277_out));
  LUT6 #(
    .INIT(64'h69966996FF0000FF)) 
    \base_new_pp[5]_i_1 
       (.I0(\CD[0].col_reg[3][25] ),
        .I1(\CD[0].col_reg[3][29] ),
        .I2(\CD[0].col_reg[3][24] ),
        .I3(\CD[0].col_reg[3][30] ),
        .I4(\CD[0].col_reg[3][28] ),
        .I5(enc_dec_sbox),
        .O(p_1_in7_in));
  LUT6 #(
    .INIT(64'h3CC3C33CA55A5AA5)) 
    \base_new_pp[6]_i_1 
       (.I0(\CD[0].col_reg[3][25] ),
        .I1(\CD[0].col_reg[3][29] ),
        .I2(\CD[0].col_reg[3][24] ),
        .I3(\CD[0].col_reg[3][30] ),
        .I4(\CD[0].col_reg[3][28] ),
        .I5(enc_dec_sbox),
        .O(p_1_in10_in));
  LUT6 #(
    .INIT(64'h3CC36666C33C6666)) 
    \base_new_pp[7]_i_1 
       (.I0(\CD[0].col_reg[3][28] ),
        .I1(\CD[0].col_reg[3][31] ),
        .I2(\CD[0].col_reg[3][29] ),
        .I3(\CD[0].col_reg[3][26] ),
        .I4(enc_dec_sbox),
        .I5(isomorphism_return179_out),
        .O(p_1_in18_in));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\base_new_pp[0]_i_1_n_0 ),
        .Q(\base_new_pp_reg_n_0_[0] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in),
        .Q(\base_new_pp_reg_n_0_[1] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_0_in9_in),
        .Q(in21_in[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in17_in),
        .Q(in21_in[1]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[4] 
       (.C(clk_i),
        .CE(1'b1),
        .D(\base_new_pp[4]_i_1_n_0 ),
        .Q(\base_new_pp_reg_n_0_[4] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[5] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in7_in),
        .Q(\base_new_pp_reg_n_0_[5] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[6] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in10_in),
        .Q(in2[0]),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \base_new_pp_reg[7] 
       (.C(clk_i),
        .CE(1'b1),
        .D(p_1_in18_in),
        .Q(in2[1]),
        .R(1'b0));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[24]_INST_0_i_10 
       (.I0(\CD[0].col[3][31]_i_14 [0]),
        .I1(\CD[0].col[3][31]_i_14_0 ),
        .I2(\CD[0].col[3][31]_i_14_1 [0]),
        .I3(\CD[0].col[3][31]_i_14_2 ),
        .O(\CD[2].col_reg[1][24] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[24]_INST_0_i_5 
       (.I0(\base_new_pp_reg[4]_0 ),
        .I1(\base_new_pp_reg[2]_0 [0]),
        .I2(\info_o[24]_INST_0_i_9_n_0 ),
        .I3(\CD[2].col_reg[1][24] ),
        .O(\CD[0].col_reg[3][24] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[24]_INST_0_i_9 
       (.I0(\info_o[31]_INST_0_i_9_0 [0]),
        .I1(\base_new_pp[4]_i_2_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_9_1 [0]),
        .I4(\info_o[31]_INST_0_i_9_2 [0]),
        .I5(\base_new_pp[4]_i_2_1 ),
        .O(\info_o[24]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[25]_INST_0_i_10 
       (.I0(\CD[0].col[3][31]_i_14 [1]),
        .I1(\CD[0].col[3][31]_i_14_0 ),
        .I2(\CD[0].col[3][31]_i_14_1 [1]),
        .I3(\CD[0].col[3][31]_i_14_2 ),
        .O(\CD[2].col_reg[1][25] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[25]_INST_0_i_5 
       (.I0(\base_new_pp_reg[4]_0 ),
        .I1(\base_new_pp_reg[2]_0 [1]),
        .I2(\info_o[25]_INST_0_i_9_n_0 ),
        .I3(\CD[2].col_reg[1][25] ),
        .O(\CD[0].col_reg[3][25] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[25]_INST_0_i_9 
       (.I0(\info_o[31]_INST_0_i_9_0 [1]),
        .I1(\base_new_pp[4]_i_2_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_9_1 [1]),
        .I4(\info_o[31]_INST_0_i_9_2 [1]),
        .I5(\base_new_pp[4]_i_2_1 ),
        .O(\info_o[25]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[26]_INST_0_i_10 
       (.I0(\CD[0].col[3][31]_i_14 [2]),
        .I1(\CD[0].col[3][31]_i_14_0 ),
        .I2(\CD[0].col[3][31]_i_14_1 [2]),
        .I3(\CD[0].col[3][31]_i_14_2 ),
        .O(\CD[2].col_reg[1][26] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[26]_INST_0_i_5 
       (.I0(\base_new_pp_reg[4]_0 ),
        .I1(\base_new_pp_reg[2]_0 [2]),
        .I2(\info_o[26]_INST_0_i_9_n_0 ),
        .I3(\CD[2].col_reg[1][26] ),
        .O(\CD[0].col_reg[3][26] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[26]_INST_0_i_9 
       (.I0(\info_o[31]_INST_0_i_9_0 [2]),
        .I1(\base_new_pp[4]_i_2_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_9_1 [2]),
        .I4(\info_o[31]_INST_0_i_9_2 [2]),
        .I5(\base_new_pp[4]_i_2_1 ),
        .O(\info_o[26]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[27]_INST_0_i_10 
       (.I0(\CD[0].col[3][31]_i_14 [3]),
        .I1(\CD[0].col[3][31]_i_14_0 ),
        .I2(\CD[0].col[3][31]_i_14_1 [3]),
        .I3(\CD[0].col[3][31]_i_14_2 ),
        .O(\CD[2].col_reg[1][27] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[27]_INST_0_i_5 
       (.I0(\base_new_pp_reg[4]_0 ),
        .I1(\base_new_pp_reg[2]_0 [3]),
        .I2(\info_o[27]_INST_0_i_9_n_0 ),
        .I3(\CD[2].col_reg[1][27] ),
        .O(\CD[0].col_reg[3][27] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[27]_INST_0_i_9 
       (.I0(\info_o[31]_INST_0_i_9_0 [3]),
        .I1(\base_new_pp[4]_i_2_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_9_1 [3]),
        .I4(\info_o[31]_INST_0_i_9_2 [3]),
        .I5(\base_new_pp[4]_i_2_1 ),
        .O(\info_o[27]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[28]_INST_0_i_11 
       (.I0(\info_o[31]_INST_0_i_9_0 [4]),
        .I1(\base_new_pp[4]_i_2_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_9_1 [4]),
        .I4(\info_o[31]_INST_0_i_9_2 [4]),
        .I5(\base_new_pp[4]_i_2_1 ),
        .O(\info_o[28]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[28]_INST_0_i_12 
       (.I0(\CD[0].col[3][31]_i_14 [4]),
        .I1(\CD[0].col[3][31]_i_14_0 ),
        .I2(\CD[0].col[3][31]_i_14_1 [4]),
        .I3(\CD[0].col[3][31]_i_14_2 ),
        .O(\CD[2].col_reg[1][28] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[28]_INST_0_i_5 
       (.I0(\base_new_pp_reg[4]_0 ),
        .I1(\base_new_pp_reg[2]_0 [4]),
        .I2(\info_o[28]_INST_0_i_11_n_0 ),
        .I3(\CD[2].col_reg[1][28] ),
        .O(\CD[0].col_reg[3][28] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[29]_INST_0_i_11 
       (.I0(\info_o[31]_INST_0_i_9_0 [5]),
        .I1(\base_new_pp[4]_i_2_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_9_1 [5]),
        .I4(\info_o[31]_INST_0_i_9_2 [5]),
        .I5(\base_new_pp[4]_i_2_1 ),
        .O(\info_o[29]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[29]_INST_0_i_12 
       (.I0(\CD[0].col[3][31]_i_14 [5]),
        .I1(\CD[0].col[3][31]_i_14_0 ),
        .I2(\CD[0].col[3][31]_i_14_1 [5]),
        .I3(\CD[0].col[3][31]_i_14_2 ),
        .O(\CD[2].col_reg[1][29] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[29]_INST_0_i_5 
       (.I0(\base_new_pp_reg[4]_0 ),
        .I1(\base_new_pp_reg[2]_0 [5]),
        .I2(\info_o[29]_INST_0_i_11_n_0 ),
        .I3(\CD[2].col_reg[1][29] ),
        .O(\CD[0].col_reg[3][29] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[30]_INST_0_i_11 
       (.I0(\info_o[31]_INST_0_i_9_0 [6]),
        .I1(\base_new_pp[4]_i_2_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_9_1 [6]),
        .I4(\info_o[31]_INST_0_i_9_2 [6]),
        .I5(\base_new_pp[4]_i_2_1 ),
        .O(\info_o[30]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[30]_INST_0_i_12 
       (.I0(\CD[0].col[3][31]_i_14 [6]),
        .I1(\CD[0].col[3][31]_i_14_0 ),
        .I2(\CD[0].col[3][31]_i_14_1 [6]),
        .I3(\CD[0].col[3][31]_i_14_2 ),
        .O(\CD[2].col_reg[1][30] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[30]_INST_0_i_5 
       (.I0(\base_new_pp_reg[4]_0 ),
        .I1(\base_new_pp_reg[2]_0 [6]),
        .I2(\info_o[30]_INST_0_i_11_n_0 ),
        .I3(\CD[2].col_reg[1][30] ),
        .O(\CD[0].col_reg[3][30] ));
  LUT6 #(
    .INIT(64'hF8FF8F8888888888)) 
    \info_o[31]_INST_0_i_20 
       (.I0(\info_o[31]_INST_0_i_9_0 [7]),
        .I1(\base_new_pp[4]_i_2_0 ),
        .I2(enc_dec_sbox),
        .I3(\info_o[31]_INST_0_i_9_1 [7]),
        .I4(\info_o[31]_INST_0_i_9_2 [7]),
        .I5(\base_new_pp[4]_i_2_1 ),
        .O(\info_o[31]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \info_o[31]_INST_0_i_21 
       (.I0(\CD[0].col[3][31]_i_14 [7]),
        .I1(\CD[0].col[3][31]_i_14_0 ),
        .I2(\CD[0].col[3][31]_i_14_1 [7]),
        .I3(\CD[0].col[3][31]_i_14_2 ),
        .O(\CD[2].col_reg[1][31] ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \info_o[31]_INST_0_i_9 
       (.I0(\base_new_pp_reg[4]_0 ),
        .I1(\base_new_pp_reg[2]_0 [7]),
        .I2(\info_o[31]_INST_0_i_20_n_0 ),
        .I3(\CD[2].col_reg[1][31] ),
        .O(\CD[0].col_reg[3][31] ));
  LUT6 #(
    .INIT(64'hA9A69A955659656A)) 
    \out_gf_pp[0]_i_1 
       (.I0(gf_inv_8_stage1_return2__0),
        .I1(p_1_in7_in),
        .I2(p_0_in),
        .I3(\base_new_pp[4]_i_1_n_0 ),
        .I4(\base_new_pp[0]_i_1_n_0 ),
        .I5(gf_inv_8_stage1_return1__0),
        .O(gf_inv_8_stage1_return[0]));
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT4 #(
    .INIT(16'hF99F)) 
    \out_gf_pp[0]_i_2 
       (.I0(p_1_in18_in),
        .I1(p_1_in7_in),
        .I2(p_1_in17_in),
        .I3(p_0_in),
        .O(gf_inv_8_stage1_return2__0));
  LUT6 #(
    .INIT(64'h9999969699666996)) 
    \out_gf_pp[1]_i_1 
       (.I0(gf_inv_8_stage1_return1__0),
        .I1(gf_inv_8_stage1_return349_in),
        .I2(\out_gf_pp[1]_i_3_n_0 ),
        .I3(\out_gf_pp[3]_i_5_n_0 ),
        .I4(\out_gf_pp[3]_i_6_n_0 ),
        .I5(\out_gf_pp[1]_i_4_n_0 ),
        .O(gf_inv_8_stage1_return[1]));
  LUT6 #(
    .INIT(64'hF5C5FFCFFFCFFACA)) 
    \out_gf_pp[1]_i_2 
       (.I0(\CD[0].col_reg[3][30] ),
        .I1(\CD[0].col_reg[3][25] ),
        .I2(enc_dec_sbox),
        .I3(isomorphism_return114_out),
        .I4(p_72_in),
        .I5(\CD[0].col_reg[3][28] ),
        .O(gf_inv_8_stage1_return349_in));
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[1]_i_3 
       (.I0(\base_new_pp[4]_i_1_n_0 ),
        .I1(p_1_in7_in),
        .O(\out_gf_pp[1]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[1]_i_4 
       (.I0(p_1_in18_in),
        .I1(p_1_in10_in),
        .O(\out_gf_pp[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h6A6A6A959595956A)) 
    \out_gf_pp[2]_i_1 
       (.I0(\out_gf_pp[2]_i_2_n_0 ),
        .I1(p_1_in10_in),
        .I2(p_0_in9_in),
        .I3(gf_inv_8_stage1_return542_out),
        .I4(gf_inv_8_stage1_return540_out),
        .I5(gf_inv_8_stage1_return1__0),
        .O(gf_inv_8_stage1_return[2]));
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT4 #(
    .INIT(16'hF99F)) 
    \out_gf_pp[2]_i_2 
       (.I0(p_0_in9_in),
        .I1(p_1_in17_in),
        .I2(p_1_in10_in),
        .I3(p_1_in18_in),
        .O(\out_gf_pp[2]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[2]_i_3 
       (.I0(p_1_in7_in),
        .I1(p_1_in18_in),
        .O(gf_inv_8_stage1_return542_out));
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[2]_i_4 
       (.I0(p_0_in),
        .I1(p_1_in17_in),
        .O(gf_inv_8_stage1_return540_out));
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT5 #(
    .INIT(32'hF9F9F99F)) 
    \out_gf_pp[2]_i_5 
       (.I0(p_1_in10_in),
        .I1(\base_new_pp[4]_i_1_n_0 ),
        .I2(p_0_in9_in),
        .I3(\out_gf_pp[2]_i_6_n_0 ),
        .I4(\out_gf_pp[2]_i_7_n_0 ),
        .O(gf_inv_8_stage1_return1__0));
  LUT6 #(
    .INIT(64'h9669000069960000)) 
    \out_gf_pp[2]_i_6 
       (.I0(\CD[0].col_reg[3][25] ),
        .I1(\CD[0].col_reg[3][24] ),
        .I2(\CD[0].col_reg[3][30] ),
        .I3(\CD[0].col_reg[3][27] ),
        .I4(enc_dec_sbox),
        .I5(\CD[0].col_reg[3][26] ),
        .O(\out_gf_pp[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000966900006996)) 
    \out_gf_pp[2]_i_7 
       (.I0(\CD[0].col_reg[3][29] ),
        .I1(\CD[0].col_reg[3][24] ),
        .I2(\CD[0].col_reg[3][30] ),
        .I3(\CD[0].col_reg[3][28] ),
        .I4(enc_dec_sbox),
        .I5(\CD[0].col_reg[3][25] ),
        .O(\out_gf_pp[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h5656565656A9A956)) 
    \out_gf_pp[3]_i_1 
       (.I0(\out_gf_pp[3]_i_2_n_0 ),
        .I1(gf_inv_8_stage1_return547_out),
        .I2(gf_inv_8_stage1_return546_out),
        .I3(\out_gf_pp[3]_i_5_n_0 ),
        .I4(\out_gf_pp[3]_i_6_n_0 ),
        .I5(\out_gf_pp[3]_i_7_n_0 ),
        .O(gf_inv_8_stage1_return[3]));
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT4 #(
    .INIT(16'hA6C0)) 
    \out_gf_pp[3]_i_2 
       (.I0(p_1_in18_in),
        .I1(p_1_in10_in),
        .I2(p_1_in17_in),
        .I3(p_0_in9_in),
        .O(\out_gf_pp[3]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[3]_i_3 
       (.I0(\base_new_pp[4]_i_1_n_0 ),
        .I1(p_1_in10_in),
        .O(gf_inv_8_stage1_return547_out));
  LUT6 #(
    .INIT(64'hDE1212DE21EDED21)) 
    \out_gf_pp[3]_i_4 
       (.I0(isomorphism_return076_out),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][25] ),
        .I3(isomorphism_return1__0),
        .I4(\CD[0].col_reg[3][26] ),
        .I5(p_0_in9_in),
        .O(gf_inv_8_stage1_return546_out));
  LUT6 #(
    .INIT(64'hDE1212DE21EDED21)) 
    \out_gf_pp[3]_i_5 
       (.I0(isomorphism_return076_out),
        .I1(enc_dec_sbox),
        .I2(\CD[0].col_reg[3][25] ),
        .I3(isomorphism_return1__0),
        .I4(\CD[0].col_reg[3][26] ),
        .I5(p_0_in),
        .O(\out_gf_pp[3]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_gf_pp[3]_i_6 
       (.I0(p_1_in17_in),
        .I1(p_0_in9_in),
        .O(\out_gf_pp[3]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \out_gf_pp[3]_i_7 
       (.I0(p_1_in10_in),
        .I1(p_1_in18_in),
        .I2(p_1_in7_in),
        .I3(\base_new_pp[4]_i_1_n_0 ),
        .O(\out_gf_pp[3]_i_7_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[0] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[0]),
        .Q(\out_gf_pp_reg_n_0_[0] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[1] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[1]),
        .Q(\out_gf_pp_reg_n_0_[1] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[2] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[2]),
        .Q(\out_gf_pp_reg_n_0_[2] ),
        .R(1'b0));
  FDRE #(
    .INIT(1'b0)) 
    \out_gf_pp_reg[3] 
       (.C(clk_i),
        .CE(1'b1),
        .D(gf_inv_8_stage1_return[3]),
        .Q(\out_gf_pp_reg_n_0_[3] ),
        .R(1'b0));
  LUT5 #(
    .INIT(32'h99990FF0)) 
    \sbox_pp2[24]_i_1 
       (.I0(p_95_in),
        .I1(gf_inv_8_stage2_return0__3),
        .I2(sbox_out_dec),
        .I3(\sbox_pp2_reg[24] ),
        .I4(\sbox_pp2_reg[31] ),
        .O(D[0]));
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT5 #(
    .INIT(32'h66999696)) 
    \sbox_pp2[25]_i_1 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(p_1_in),
        .I2(\sbox_pp2_reg[25] ),
        .I3(p_0_in2_in),
        .I4(\sbox_pp2_reg[31] ),
        .O(D[1]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[25]_i_2 
       (.I0(\base_new_pp_reg_n_0_[0] ),
        .I1(gf_muls_20_return__1[0]),
        .I2(gf_muls_20_return__1[1]),
        .I3(\base_new_pp_reg_n_0_[1] ),
        .I4(gf_muls_scl_2_return[1]),
        .O(p_1_in));
  LUT6 #(
    .INIT(64'h99999999F00F0FF0)) 
    \sbox_pp2[26]_i_1 
       (.I0(p_92_in),
        .I1(p_93_in),
        .I2(p_16_in),
        .I3(gf_inv_8_stage2_return013_out[1]),
        .I4(\sbox_pp2_reg[26] ),
        .I5(\sbox_pp2_reg[31] ),
        .O(D[2]));
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \sbox_pp2[26]_i_2 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(p_1_in),
        .I2(p_0_in2_in),
        .O(p_16_in));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[26]_i_3 
       (.I0(in21_in[0]),
        .I1(in1__0[0]),
        .I2(in1__0[1]),
        .I3(in21_in[1]),
        .I4(gf_muls_scl_2_return[1]),
        .O(gf_inv_8_stage2_return013_out[1]));
  LUT6 #(
    .INIT(64'h0FF0666669960000)) 
    \sbox_pp2[26]_i_4 
       (.I0(in21_in[1]),
        .I1(\base_new_pp_reg_n_0_[1] ),
        .I2(in21_in[0]),
        .I3(\base_new_pp_reg_n_0_[0] ),
        .I4(in111_out[1]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_2_return[1]));
  LUT6 #(
    .INIT(64'hAA55AA5596966969)) 
    \sbox_pp2[27]_i_1 
       (.I0(p_95_in),
        .I1(gf_inv_8_stage2_return0__3),
        .I2(p_92_in),
        .I3(isomorphism_inv_return03_out),
        .I4(\sbox_pp2_reg[27] ),
        .I5(\sbox_pp2_reg[31] ),
        .O(D[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \sbox_pp2[27]_i_2 
       (.I0(p_0_in2_in),
        .I1(gf_inv_8_stage2_return013_out[0]),
        .O(p_95_in));
  LUT2 #(
    .INIT(4'h6)) 
    \sbox_pp2[27]_i_3 
       (.I0(isomorphism_inv_return05_out),
        .I1(sbox_out_dec),
        .O(p_92_in));
  LUT5 #(
    .INIT(32'h00FF9696)) 
    \sbox_pp2[28]_i_1 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(gf_inv_8_stage2_return013_out[0]),
        .I2(\sbox_pp2_reg[28] ),
        .I3(isomorphism_inv_return03_out),
        .I4(\sbox_pp2_reg[31] ),
        .O(D[4]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[28]_i_2 
       (.I0(in21_in[1]),
        .I1(in1__0[1]),
        .I2(in1__0[0]),
        .I3(in21_in[0]),
        .I4(gf_muls_scl_2_return[0]),
        .O(gf_inv_8_stage2_return013_out[0]));
  LUT5 #(
    .INIT(32'h00FF9669)) 
    \sbox_pp2[29]_i_1 
       (.I0(isomorphism_inv_return03_out),
        .I1(sbox_out_dec),
        .I2(\sbox_pp2_reg[29] ),
        .I3(p_93_in),
        .I4(\sbox_pp2_reg[31] ),
        .O(D[5]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[29]_i_2 
       (.I0(in2[1]),
        .I1(in1__0[1]),
        .I2(in1__0[0]),
        .I3(in2[0]),
        .I4(gf_muls_scl_20_return[0]),
        .O(sbox_out_dec));
  LUT6 #(
    .INIT(64'h0000FFFF96699669)) 
    \sbox_pp2[30]_i_1 
       (.I0(isomorphism_inv_return03_out),
        .I1(p_93_in),
        .I2(gf_inv_8_stage2_return0__3),
        .I3(\sbox_pp2_reg[30] ),
        .I4(isomorphism_inv_return033_out),
        .I5(\sbox_pp2_reg[31] ),
        .O(D[6]));
  LUT2 #(
    .INIT(4'h9)) 
    \sbox_pp2[30]_i_2 
       (.I0(isomorphism_inv_return033_out),
        .I1(p_1_in),
        .O(isomorphism_inv_return03_out));
  LUT6 #(
    .INIT(64'h96A59955695A66AA)) 
    \sbox_pp2[30]_i_3 
       (.I0(gf_muls_scl_20_return[0]),
        .I1(\base_new_pp_reg_n_0_[4] ),
        .I2(gf_muls_20_return__1[0]),
        .I3(gf_muls_20_return__1[1]),
        .I4(\base_new_pp_reg_n_0_[5] ),
        .I5(gf_inv_8_stage2_return013_out[0]),
        .O(p_93_in));
  LUT6 #(
    .INIT(64'hE4281BD71BD7E428)) 
    \sbox_pp2[30]_i_4 
       (.I0(in2[0]),
        .I1(in1__0[0]),
        .I2(in1__0[1]),
        .I3(in2[1]),
        .I4(gf_muls_scl_20_return[1]),
        .I5(gf_inv_8_stage2_return013_out[1]),
        .O(isomorphism_inv_return033_out));
  LUT6 #(
    .INIT(64'h609F9F6060606060)) 
    \sbox_pp2[30]_i_5 
       (.I0(\base_new_pp_reg_n_0_[5] ),
        .I1(in2[1]),
        .I2(in111_out[1]),
        .I3(\base_new_pp_reg_n_0_[4] ),
        .I4(in2[0]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_20_return[0]));
  LUT5 #(
    .INIT(32'h00FF9696)) 
    \sbox_pp2[31]_i_1 
       (.I0(gf_inv_8_stage2_return0__3),
        .I1(p_0_in2_in),
        .I2(\sbox_pp2_reg[31]_0 ),
        .I3(isomorphism_inv_return05_out),
        .I4(\sbox_pp2_reg[31] ),
        .O(D[7]));
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT4 #(
    .INIT(16'hB2E2)) 
    \sbox_pp2[31]_i_10 
       (.I0(\out_gf_pp_reg_n_0_[0] ),
        .I1(\out_gf_pp_reg_n_0_[2] ),
        .I2(\out_gf_pp_reg_n_0_[1] ),
        .I3(\out_gf_pp_reg_n_0_[3] ),
        .O(in1__0[0]));
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT4 #(
    .INIT(16'hE4C6)) 
    \sbox_pp2[31]_i_11 
       (.I0(\out_gf_pp_reg_n_0_[1] ),
        .I1(\out_gf_pp_reg_n_0_[0] ),
        .I2(\out_gf_pp_reg_n_0_[3] ),
        .I3(\out_gf_pp_reg_n_0_[2] ),
        .O(in1__0[1]));
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT4 #(
    .INIT(16'h23D6)) 
    \sbox_pp2[31]_i_12 
       (.I0(\out_gf_pp_reg_n_0_[2] ),
        .I1(\out_gf_pp_reg_n_0_[3] ),
        .I2(\out_gf_pp_reg_n_0_[0] ),
        .I3(\out_gf_pp_reg_n_0_[1] ),
        .O(in111_out[1]));
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT4 #(
    .INIT(16'h6DB0)) 
    \sbox_pp2[31]_i_13 
       (.I0(\out_gf_pp_reg_n_0_[3] ),
        .I1(\out_gf_pp_reg_n_0_[1] ),
        .I2(\out_gf_pp_reg_n_0_[2] ),
        .I3(\out_gf_pp_reg_n_0_[0] ),
        .O(in111_out[0]));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[31]_i_2 
       (.I0(\base_new_pp_reg_n_0_[4] ),
        .I1(gf_muls_20_return__1[0]),
        .I2(gf_muls_20_return__1[1]),
        .I3(\base_new_pp_reg_n_0_[5] ),
        .I4(gf_muls_scl_20_return[1]),
        .O(gf_inv_8_stage2_return0__3));
  LUT5 #(
    .INIT(32'h1BD7E428)) 
    \sbox_pp2[31]_i_3 
       (.I0(\base_new_pp_reg_n_0_[1] ),
        .I1(gf_muls_20_return__1[1]),
        .I2(gf_muls_20_return__1[0]),
        .I3(\base_new_pp_reg_n_0_[0] ),
        .I4(gf_muls_scl_2_return[0]),
        .O(p_0_in2_in));
  LUT6 #(
    .INIT(64'h1BD7E428E4281BD7)) 
    \sbox_pp2[31]_i_4 
       (.I0(in2[0]),
        .I1(in1__0[0]),
        .I2(in1__0[1]),
        .I3(in2[1]),
        .I4(gf_muls_scl_20_return[1]),
        .I5(p_1_in),
        .O(isomorphism_inv_return05_out));
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT4 #(
    .INIT(16'hBE22)) 
    \sbox_pp2[31]_i_6 
       (.I0(\out_gf_pp_reg_n_0_[2] ),
        .I1(\out_gf_pp_reg_n_0_[0] ),
        .I2(\out_gf_pp_reg_n_0_[1] ),
        .I3(\out_gf_pp_reg_n_0_[3] ),
        .O(gf_muls_20_return__1[0]));
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT4 #(
    .INIT(16'hDD82)) 
    \sbox_pp2[31]_i_7 
       (.I0(\out_gf_pp_reg_n_0_[3] ),
        .I1(\out_gf_pp_reg_n_0_[1] ),
        .I2(\out_gf_pp_reg_n_0_[0] ),
        .I3(\out_gf_pp_reg_n_0_[2] ),
        .O(gf_muls_20_return__1[1]));
  LUT6 #(
    .INIT(64'h0FF0666669960000)) 
    \sbox_pp2[31]_i_8 
       (.I0(in2[1]),
        .I1(\base_new_pp_reg_n_0_[5] ),
        .I2(in2[0]),
        .I3(\base_new_pp_reg_n_0_[4] ),
        .I4(in111_out[1]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_20_return[1]));
  LUT6 #(
    .INIT(64'h609F9F6060606060)) 
    \sbox_pp2[31]_i_9 
       (.I0(\base_new_pp_reg_n_0_[1] ),
        .I1(in21_in[1]),
        .I2(in111_out[1]),
        .I3(\base_new_pp_reg_n_0_[0] ),
        .I4(in21_in[0]),
        .I5(in111_out[0]),
        .O(gf_muls_scl_2_return[0]));
endmodule
`ifndef GLBL
`define GLBL
`timescale  1 ps / 1 ps

module glbl ();

    parameter ROC_WIDTH = 100000;
    parameter TOC_WIDTH = 0;

//--------   STARTUP Globals --------------
    wire GSR;
    wire GTS;
    wire GWE;
    wire PRLD;
    tri1 p_up_tmp;
    tri (weak1, strong0) PLL_LOCKG = p_up_tmp;

    wire PROGB_GLBL;
    wire CCLKO_GLBL;
    wire FCSBO_GLBL;
    wire [3:0] DO_GLBL;
    wire [3:0] DI_GLBL;
   
    reg GSR_int;
    reg GTS_int;
    reg PRLD_int;

//--------   JTAG Globals --------------
    wire JTAG_TDO_GLBL;
    wire JTAG_TCK_GLBL;
    wire JTAG_TDI_GLBL;
    wire JTAG_TMS_GLBL;
    wire JTAG_TRST_GLBL;

    reg JTAG_CAPTURE_GLBL;
    reg JTAG_RESET_GLBL;
    reg JTAG_SHIFT_GLBL;
    reg JTAG_UPDATE_GLBL;
    reg JTAG_RUNTEST_GLBL;

    reg JTAG_SEL1_GLBL = 0;
    reg JTAG_SEL2_GLBL = 0 ;
    reg JTAG_SEL3_GLBL = 0;
    reg JTAG_SEL4_GLBL = 0;

    reg JTAG_USER_TDO1_GLBL = 1'bz;
    reg JTAG_USER_TDO2_GLBL = 1'bz;
    reg JTAG_USER_TDO3_GLBL = 1'bz;
    reg JTAG_USER_TDO4_GLBL = 1'bz;

    assign (strong1, weak0) GSR = GSR_int;
    assign (strong1, weak0) GTS = GTS_int;
    assign (weak1, weak0) PRLD = PRLD_int;

    initial begin
	GSR_int = 1'b1;
	PRLD_int = 1'b1;
	#(ROC_WIDTH)
	GSR_int = 1'b0;
	PRLD_int = 1'b0;
    end

    initial begin
	GTS_int = 1'b1;
	#(TOC_WIDTH)
	GTS_int = 1'b0;
    end

endmodule
`endif
