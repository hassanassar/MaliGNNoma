`timescale 1 ps / 1 ps
`define XIL_TIMING

(* dont_touch = "true" *) 
(* NotValidForBitStream *)
module switch_elements
   (enable_i,
    clk_i,
    rst_i,
    info_o);
  input [31:0]enable_i;
  input clk_i;
  input rst_i;
  output [31:0]info_o;

  wire [31:0]enable_i;
  wire [31:0]info_o;

  (* BOX_TYPE = "black_box" *) 
  (* DONT_TOUCH *) 
  switch_elements_muxer__1 \activity_blocks[0].switch 
       (.enable_i(enable_i[0]),
        .info_o(info_o[0]));
  (* BOX_TYPE = "black_box" *) 
  (* DONT_TOUCH *) 
  switch_elements_muxer__2 \activity_blocks[1].switch 
       (.enable_i(enable_i[1]),
        .info_o(info_o[1]));
  (* BOX_TYPE = "black_box" *) 
  (* DONT_TOUCH *) 
  switch_elements_muxer__3 \activity_blocks[2].switch 
       (.enable_i(enable_i[2]),
        .info_o(info_o[2]));
  (* BOX_TYPE = "black_box" *) 
  (* DONT_TOUCH *) 
  switch_elements_muxer__4 \activity_blocks[3].switch 
       (.enable_i(enable_i[3]),
        .info_o(info_o[3]));
  (* BOX_TYPE = "black_box" *) 
  (* DONT_TOUCH *) 
  switch_elements_muxer__5 \activity_blocks[4].switch 
       (.enable_i(enable_i[4]),
        .info_o(info_o[4]));
  (* BOX_TYPE = "black_box" *) 
  (* DONT_TOUCH *) 
  switch_elements_muxer__6 \activity_blocks[5].switch 
       (.enable_i(enable_i[5]),
        .info_o(info_o[5]));
  (* BOX_TYPE = "black_box" *) 
  (* DONT_TOUCH *) 
  switch_elements_muxer__7 \activity_blocks[6].switch 
       (.enable_i(enable_i[6]),
        .info_o(info_o[6]));
  (* BOX_TYPE = "black_box" *) 
  (* DONT_TOUCH *) 
  switch_elements_muxer \activity_blocks[7].switch 
       (.enable_i(enable_i[7]),
        .info_o(info_o[7]));
endmodule

(* ORIG_REF_NAME = "muxer" *) (* box_type = "black_box" *) (* dont_touch = "true" *) 
module switch_elements_muxer
   (enable_i,
    info_o);
  input enable_i;
  output info_o;

  wire enable_i;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf7;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf8;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf9;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [1802:0]self_sf7;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf8;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf9;

  assign info_o = info_sf7[1];
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[0]),
        .S(info_sf7[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1000].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1000]),
        .S(self_sf7[1000]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1001].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1001]),
        .S(self_sf7[1001]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1002].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1002]),
        .S(self_sf7[1002]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1003].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1003]),
        .S(self_sf7[1003]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1004].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1004]),
        .S(self_sf7[1004]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1005].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1005]),
        .S(self_sf7[1005]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1006].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1006]),
        .S(self_sf7[1006]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1007].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1007]),
        .S(self_sf7[1007]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1008].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1008]),
        .S(self_sf7[1008]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1009].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1009]),
        .S(self_sf7[1009]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[100]),
        .S(self_sf7[100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1010].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1010]),
        .S(self_sf7[1010]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1011].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1011]),
        .S(self_sf7[1011]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1012].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1012]),
        .S(self_sf7[1012]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1013].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1013]),
        .S(self_sf7[1013]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1014].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1014]),
        .S(self_sf7[1014]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1015].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1015]),
        .S(self_sf7[1015]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1016].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1016]),
        .S(self_sf7[1016]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1017].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1017]),
        .S(self_sf7[1017]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1018].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1018]),
        .S(self_sf7[1018]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1019].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1019]),
        .S(self_sf7[1019]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[101]),
        .S(self_sf7[101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1020].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1020]),
        .S(self_sf7[1020]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1021].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1021]),
        .S(self_sf7[1021]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1022].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1022]),
        .S(self_sf7[1022]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1023].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1023]),
        .S(self_sf7[1023]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1024].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1024]),
        .S(self_sf7[1024]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1025].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1025]),
        .S(self_sf7[1025]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1026].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1026]),
        .S(self_sf7[1026]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1027].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1027]),
        .S(self_sf7[1027]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1028].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1028]),
        .S(self_sf7[1028]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1029].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1029]),
        .S(self_sf7[1029]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[102]),
        .S(self_sf7[102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1030].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1030]),
        .S(self_sf7[1030]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1031].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1031]),
        .S(self_sf7[1031]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1032].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1032]),
        .S(self_sf7[1032]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1033].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1033]),
        .S(self_sf7[1033]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1034].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1034]),
        .S(self_sf7[1034]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1035].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1035]),
        .S(self_sf7[1035]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1036].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1036]),
        .S(self_sf7[1036]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1037].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1037]),
        .S(self_sf7[1037]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1038].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1038]),
        .S(self_sf7[1038]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1039].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1039]),
        .S(self_sf7[1039]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[103]),
        .S(self_sf7[103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1040].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1040]),
        .S(self_sf7[1040]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1041].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1041]),
        .S(self_sf7[1041]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1042].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1042]),
        .S(self_sf7[1042]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1043].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1043]),
        .S(self_sf7[1043]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1044].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1044]),
        .S(self_sf7[1044]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1045].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1045]),
        .S(self_sf7[1045]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1046].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1046]),
        .S(self_sf7[1046]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1047].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1047]),
        .S(self_sf7[1047]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1048].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1048]),
        .S(self_sf7[1048]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1049].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1049]),
        .S(self_sf7[1049]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[104]),
        .S(self_sf7[104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1050].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1050]),
        .S(self_sf7[1050]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1051].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1051]),
        .S(self_sf7[1051]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1052].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1052]),
        .S(self_sf7[1052]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1053].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1053]),
        .S(self_sf7[1053]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1054].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1054]),
        .S(self_sf7[1054]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1055].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1055]),
        .S(self_sf7[1055]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1056].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1056]),
        .S(self_sf7[1056]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1057].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1057]),
        .S(self_sf7[1057]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1058].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1058]),
        .S(self_sf7[1058]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1059].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1059]),
        .S(self_sf7[1059]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[105]),
        .S(self_sf7[105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1060].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1060]),
        .S(self_sf7[1060]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1061].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1061]),
        .S(self_sf7[1061]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1062].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1062]),
        .S(self_sf7[1062]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1063].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1063]),
        .S(self_sf7[1063]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1064].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1064]),
        .S(self_sf7[1064]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1065].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1065]),
        .S(self_sf7[1065]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1066].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1066]),
        .S(self_sf7[1066]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1067].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1067]),
        .S(self_sf7[1067]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1068].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1068]),
        .S(self_sf7[1068]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1069].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1069]),
        .S(self_sf7[1069]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[106]),
        .S(self_sf7[106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1070].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1070]),
        .S(self_sf7[1070]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1071].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1071]),
        .S(self_sf7[1071]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1072].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1072]),
        .S(self_sf7[1072]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1073].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1073]),
        .S(self_sf7[1073]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1074].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1074]),
        .S(self_sf7[1074]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1075].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1075]),
        .S(self_sf7[1075]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1076].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1076]),
        .S(self_sf7[1076]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1077].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1077]),
        .S(self_sf7[1077]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1078].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1078]),
        .S(self_sf7[1078]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1079].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1079]),
        .S(self_sf7[1079]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[107]),
        .S(self_sf7[107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1080].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1080]),
        .S(self_sf7[1080]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1081].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1081]),
        .S(self_sf7[1081]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1082].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1082]),
        .S(self_sf7[1082]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1083].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1083]),
        .S(self_sf7[1083]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1084].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1084]),
        .S(self_sf7[1084]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1085].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1085]),
        .S(self_sf7[1085]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1086].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1086]),
        .S(self_sf7[1086]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1087].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1087]),
        .S(self_sf7[1087]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1088].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1088]),
        .S(self_sf7[1088]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1089].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1089]),
        .S(self_sf7[1089]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[108]),
        .S(self_sf7[108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1090].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1090]),
        .S(self_sf7[1090]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1091].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1091]),
        .S(self_sf7[1091]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1092].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1092]),
        .S(self_sf7[1092]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1093].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1093]),
        .S(self_sf7[1093]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1094].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1094]),
        .S(self_sf7[1094]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1095].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1095]),
        .S(self_sf7[1095]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1096].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1096]),
        .S(self_sf7[1096]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1097].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1097]),
        .S(self_sf7[1097]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1098].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1098]),
        .S(self_sf7[1098]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1099].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1099]),
        .S(self_sf7[1099]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[109]),
        .S(self_sf7[109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[10].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[10]),
        .S(self_sf7[10]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1100]),
        .S(self_sf7[1100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1101]),
        .S(self_sf7[1101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1102]),
        .S(self_sf7[1102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1103]),
        .S(self_sf7[1103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1104]),
        .S(self_sf7[1104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1105]),
        .S(self_sf7[1105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1106]),
        .S(self_sf7[1106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1107]),
        .S(self_sf7[1107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1108]),
        .S(self_sf7[1108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1109]),
        .S(self_sf7[1109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[110]),
        .S(self_sf7[110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1110]),
        .S(self_sf7[1110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1111]),
        .S(self_sf7[1111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1112]),
        .S(self_sf7[1112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1113]),
        .S(self_sf7[1113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1114]),
        .S(self_sf7[1114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1115]),
        .S(self_sf7[1115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1116]),
        .S(self_sf7[1116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1117]),
        .S(self_sf7[1117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1118]),
        .S(self_sf7[1118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1119]),
        .S(self_sf7[1119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[111]),
        .S(self_sf7[111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1120]),
        .S(self_sf7[1120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1121]),
        .S(self_sf7[1121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1122]),
        .S(self_sf7[1122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1123]),
        .S(self_sf7[1123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1124]),
        .S(self_sf7[1124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1125]),
        .S(self_sf7[1125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1126]),
        .S(self_sf7[1126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1127]),
        .S(self_sf7[1127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1128]),
        .S(self_sf7[1128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1129]),
        .S(self_sf7[1129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[112]),
        .S(self_sf7[112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1130]),
        .S(self_sf7[1130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1131]),
        .S(self_sf7[1131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1132]),
        .S(self_sf7[1132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1133]),
        .S(self_sf7[1133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1134]),
        .S(self_sf7[1134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1135]),
        .S(self_sf7[1135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1136]),
        .S(self_sf7[1136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1137]),
        .S(self_sf7[1137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1138]),
        .S(self_sf7[1138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1139]),
        .S(self_sf7[1139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[113]),
        .S(self_sf7[113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1140]),
        .S(self_sf7[1140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1141]),
        .S(self_sf7[1141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1142]),
        .S(self_sf7[1142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1143]),
        .S(self_sf7[1143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1144]),
        .S(self_sf7[1144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1145]),
        .S(self_sf7[1145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1146]),
        .S(self_sf7[1146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1147]),
        .S(self_sf7[1147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1148]),
        .S(self_sf7[1148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1149]),
        .S(self_sf7[1149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[114]),
        .S(self_sf7[114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1150]),
        .S(self_sf7[1150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1151]),
        .S(self_sf7[1151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1152]),
        .S(self_sf7[1152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1153]),
        .S(self_sf7[1153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1154]),
        .S(self_sf7[1154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1155]),
        .S(self_sf7[1155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1156]),
        .S(self_sf7[1156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1157]),
        .S(self_sf7[1157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1158]),
        .S(self_sf7[1158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1159]),
        .S(self_sf7[1159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[115]),
        .S(self_sf7[115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1160]),
        .S(self_sf7[1160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1161]),
        .S(self_sf7[1161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1162]),
        .S(self_sf7[1162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1163]),
        .S(self_sf7[1163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1164]),
        .S(self_sf7[1164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1165]),
        .S(self_sf7[1165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1166]),
        .S(self_sf7[1166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1167]),
        .S(self_sf7[1167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1168]),
        .S(self_sf7[1168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1169]),
        .S(self_sf7[1169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[116]),
        .S(self_sf7[116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1170]),
        .S(self_sf7[1170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1171]),
        .S(self_sf7[1171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1172]),
        .S(self_sf7[1172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1173]),
        .S(self_sf7[1173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1174]),
        .S(self_sf7[1174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1175]),
        .S(self_sf7[1175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1176]),
        .S(self_sf7[1176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1177]),
        .S(self_sf7[1177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1178]),
        .S(self_sf7[1178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1179]),
        .S(self_sf7[1179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[117]),
        .S(self_sf7[117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1180]),
        .S(self_sf7[1180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1181]),
        .S(self_sf7[1181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1182]),
        .S(self_sf7[1182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1183]),
        .S(self_sf7[1183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1184]),
        .S(self_sf7[1184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1185]),
        .S(self_sf7[1185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1186]),
        .S(self_sf7[1186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1187]),
        .S(self_sf7[1187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1188]),
        .S(self_sf7[1188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1189]),
        .S(self_sf7[1189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[118]),
        .S(self_sf7[118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1190]),
        .S(self_sf7[1190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1191]),
        .S(self_sf7[1191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1192]),
        .S(self_sf7[1192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1193]),
        .S(self_sf7[1193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1194]),
        .S(self_sf7[1194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1195]),
        .S(self_sf7[1195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1196]),
        .S(self_sf7[1196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1197]),
        .S(self_sf7[1197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1198]),
        .S(self_sf7[1198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1199]),
        .S(self_sf7[1199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[119]),
        .S(self_sf7[119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[11].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[11]),
        .S(self_sf7[11]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1200]),
        .S(self_sf7[1200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1201]),
        .S(self_sf7[1201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1202]),
        .S(self_sf7[1202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1203]),
        .S(self_sf7[1203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1204]),
        .S(self_sf7[1204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1205]),
        .S(self_sf7[1205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1206]),
        .S(self_sf7[1206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1207]),
        .S(self_sf7[1207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1208]),
        .S(self_sf7[1208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1209]),
        .S(self_sf7[1209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[120]),
        .S(self_sf7[120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1210]),
        .S(self_sf7[1210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1211]),
        .S(self_sf7[1211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1212]),
        .S(self_sf7[1212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1213]),
        .S(self_sf7[1213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1214]),
        .S(self_sf7[1214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1215]),
        .S(self_sf7[1215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1216]),
        .S(self_sf7[1216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1217]),
        .S(self_sf7[1217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1218]),
        .S(self_sf7[1218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1219]),
        .S(self_sf7[1219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[121]),
        .S(self_sf7[121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1220]),
        .S(self_sf7[1220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1221]),
        .S(self_sf7[1221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1222]),
        .S(self_sf7[1222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1223]),
        .S(self_sf7[1223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1224]),
        .S(self_sf7[1224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1225]),
        .S(self_sf7[1225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1226]),
        .S(self_sf7[1226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1227]),
        .S(self_sf7[1227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1228]),
        .S(self_sf7[1228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1229]),
        .S(self_sf7[1229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[122]),
        .S(self_sf7[122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1230]),
        .S(self_sf7[1230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1231]),
        .S(self_sf7[1231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1232]),
        .S(self_sf7[1232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1233]),
        .S(self_sf7[1233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1234]),
        .S(self_sf7[1234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1235]),
        .S(self_sf7[1235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1236]),
        .S(self_sf7[1236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1237]),
        .S(self_sf7[1237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1238]),
        .S(self_sf7[1238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1239]),
        .S(self_sf7[1239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[123]),
        .S(self_sf7[123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1240]),
        .S(self_sf7[1240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1241]),
        .S(self_sf7[1241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1242]),
        .S(self_sf7[1242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1243]),
        .S(self_sf7[1243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1244]),
        .S(self_sf7[1244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1245]),
        .S(self_sf7[1245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1246]),
        .S(self_sf7[1246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1247]),
        .S(self_sf7[1247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1248]),
        .S(self_sf7[1248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1249]),
        .S(self_sf7[1249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[124]),
        .S(self_sf7[124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1250]),
        .S(self_sf7[1250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1251]),
        .S(self_sf7[1251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1252]),
        .S(self_sf7[1252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1253]),
        .S(self_sf7[1253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1254]),
        .S(self_sf7[1254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1255]),
        .S(self_sf7[1255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1256]),
        .S(self_sf7[1256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1257]),
        .S(self_sf7[1257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1258]),
        .S(self_sf7[1258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1259]),
        .S(self_sf7[1259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[125]),
        .S(self_sf7[125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1260]),
        .S(self_sf7[1260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1261]),
        .S(self_sf7[1261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1262]),
        .S(self_sf7[1262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1263]),
        .S(self_sf7[1263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1264]),
        .S(self_sf7[1264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1265]),
        .S(self_sf7[1265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1266]),
        .S(self_sf7[1266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1267]),
        .S(self_sf7[1267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1268]),
        .S(self_sf7[1268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1269]),
        .S(self_sf7[1269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[126]),
        .S(self_sf7[126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1270]),
        .S(self_sf7[1270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1271]),
        .S(self_sf7[1271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1272]),
        .S(self_sf7[1272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1273]),
        .S(self_sf7[1273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1274]),
        .S(self_sf7[1274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1275]),
        .S(self_sf7[1275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1276]),
        .S(self_sf7[1276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1277]),
        .S(self_sf7[1277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1278]),
        .S(self_sf7[1278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1279]),
        .S(self_sf7[1279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[127]),
        .S(self_sf7[127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1280]),
        .S(self_sf7[1280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1281]),
        .S(self_sf7[1281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1282]),
        .S(self_sf7[1282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1283]),
        .S(self_sf7[1283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1284]),
        .S(self_sf7[1284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1285]),
        .S(self_sf7[1285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1286]),
        .S(self_sf7[1286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1287]),
        .S(self_sf7[1287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1288]),
        .S(self_sf7[1288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1289]),
        .S(self_sf7[1289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[128]),
        .S(self_sf7[128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1290]),
        .S(self_sf7[1290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1291]),
        .S(self_sf7[1291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1292]),
        .S(self_sf7[1292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1293]),
        .S(self_sf7[1293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1294]),
        .S(self_sf7[1294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1295]),
        .S(self_sf7[1295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1296]),
        .S(self_sf7[1296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1297]),
        .S(self_sf7[1297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1298]),
        .S(self_sf7[1298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1299]),
        .S(self_sf7[1299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[129]),
        .S(self_sf7[129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[12].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[12]),
        .S(self_sf7[12]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1300]),
        .S(self_sf7[1300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1301]),
        .S(self_sf7[1301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1302]),
        .S(self_sf7[1302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1303]),
        .S(self_sf7[1303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1304]),
        .S(self_sf7[1304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1305]),
        .S(self_sf7[1305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1306]),
        .S(self_sf7[1306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1307]),
        .S(self_sf7[1307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1308]),
        .S(self_sf7[1308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1309]),
        .S(self_sf7[1309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[130]),
        .S(self_sf7[130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1310]),
        .S(self_sf7[1310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1311]),
        .S(self_sf7[1311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1312]),
        .S(self_sf7[1312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1313]),
        .S(self_sf7[1313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1314]),
        .S(self_sf7[1314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1315]),
        .S(self_sf7[1315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1316]),
        .S(self_sf7[1316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1317]),
        .S(self_sf7[1317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1318]),
        .S(self_sf7[1318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1319]),
        .S(self_sf7[1319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[131]),
        .S(self_sf7[131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1320]),
        .S(self_sf7[1320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1321]),
        .S(self_sf7[1321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1322]),
        .S(self_sf7[1322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1323]),
        .S(self_sf7[1323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1324]),
        .S(self_sf7[1324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1325]),
        .S(self_sf7[1325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1326]),
        .S(self_sf7[1326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1327]),
        .S(self_sf7[1327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1328]),
        .S(self_sf7[1328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1329]),
        .S(self_sf7[1329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[132]),
        .S(self_sf7[132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1330]),
        .S(self_sf7[1330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1331]),
        .S(self_sf7[1331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1332]),
        .S(self_sf7[1332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1333]),
        .S(self_sf7[1333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1334]),
        .S(self_sf7[1334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1335]),
        .S(self_sf7[1335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1336]),
        .S(self_sf7[1336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1337]),
        .S(self_sf7[1337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1338]),
        .S(self_sf7[1338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1339]),
        .S(self_sf7[1339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[133]),
        .S(self_sf7[133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1340]),
        .S(self_sf7[1340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1341]),
        .S(self_sf7[1341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1342]),
        .S(self_sf7[1342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1343]),
        .S(self_sf7[1343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1344]),
        .S(self_sf7[1344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1345]),
        .S(self_sf7[1345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1346]),
        .S(self_sf7[1346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1347]),
        .S(self_sf7[1347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1348]),
        .S(self_sf7[1348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1349]),
        .S(self_sf7[1349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[134]),
        .S(self_sf7[134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1350]),
        .S(self_sf7[1350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1351]),
        .S(self_sf7[1351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1352]),
        .S(self_sf7[1352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1353]),
        .S(self_sf7[1353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1354]),
        .S(self_sf7[1354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1355]),
        .S(self_sf7[1355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1356]),
        .S(self_sf7[1356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1357]),
        .S(self_sf7[1357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1358]),
        .S(self_sf7[1358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1359]),
        .S(self_sf7[1359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[135]),
        .S(self_sf7[135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1360]),
        .S(self_sf7[1360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1361]),
        .S(self_sf7[1361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1362]),
        .S(self_sf7[1362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1363]),
        .S(self_sf7[1363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1364]),
        .S(self_sf7[1364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1365]),
        .S(self_sf7[1365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1366]),
        .S(self_sf7[1366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1367]),
        .S(self_sf7[1367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1368]),
        .S(self_sf7[1368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1369]),
        .S(self_sf7[1369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[136]),
        .S(self_sf7[136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1370]),
        .S(self_sf7[1370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1371]),
        .S(self_sf7[1371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1372]),
        .S(self_sf7[1372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1373]),
        .S(self_sf7[1373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1374]),
        .S(self_sf7[1374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1375]),
        .S(self_sf7[1375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1376]),
        .S(self_sf7[1376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1377]),
        .S(self_sf7[1377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1378]),
        .S(self_sf7[1378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1379]),
        .S(self_sf7[1379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[137]),
        .S(self_sf7[137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1380]),
        .S(self_sf7[1380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1381]),
        .S(self_sf7[1381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1382]),
        .S(self_sf7[1382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1383]),
        .S(self_sf7[1383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1384]),
        .S(self_sf7[1384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1385]),
        .S(self_sf7[1385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1386]),
        .S(self_sf7[1386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1387]),
        .S(self_sf7[1387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1388]),
        .S(self_sf7[1388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1389]),
        .S(self_sf7[1389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[138]),
        .S(self_sf7[138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1390]),
        .S(self_sf7[1390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1391]),
        .S(self_sf7[1391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1392]),
        .S(self_sf7[1392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1393]),
        .S(self_sf7[1393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1394]),
        .S(self_sf7[1394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1395]),
        .S(self_sf7[1395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1396]),
        .S(self_sf7[1396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1397]),
        .S(self_sf7[1397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1398]),
        .S(self_sf7[1398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1399]),
        .S(self_sf7[1399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[139]),
        .S(self_sf7[139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[13].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[13]),
        .S(self_sf7[13]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1400]),
        .S(self_sf7[1400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1401]),
        .S(self_sf7[1401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1402]),
        .S(self_sf7[1402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1403]),
        .S(self_sf7[1403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1404]),
        .S(self_sf7[1404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1405]),
        .S(self_sf7[1405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1406]),
        .S(self_sf7[1406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1407]),
        .S(self_sf7[1407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1408]),
        .S(self_sf7[1408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1409]),
        .S(self_sf7[1409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[140]),
        .S(self_sf7[140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1410]),
        .S(self_sf7[1410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1411]),
        .S(self_sf7[1411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1412]),
        .S(self_sf7[1412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1413]),
        .S(self_sf7[1413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1414]),
        .S(self_sf7[1414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1415]),
        .S(self_sf7[1415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1416]),
        .S(self_sf7[1416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1417]),
        .S(self_sf7[1417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1418]),
        .S(self_sf7[1418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1419]),
        .S(self_sf7[1419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[141]),
        .S(self_sf7[141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1420]),
        .S(self_sf7[1420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1421]),
        .S(self_sf7[1421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1422]),
        .S(self_sf7[1422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1423]),
        .S(self_sf7[1423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1424]),
        .S(self_sf7[1424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1425]),
        .S(self_sf7[1425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1426]),
        .S(self_sf7[1426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1427]),
        .S(self_sf7[1427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1428]),
        .S(self_sf7[1428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1429]),
        .S(self_sf7[1429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[142]),
        .S(self_sf7[142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1430]),
        .S(self_sf7[1430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1431]),
        .S(self_sf7[1431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1432]),
        .S(self_sf7[1432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1433]),
        .S(self_sf7[1433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1434]),
        .S(self_sf7[1434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1435]),
        .S(self_sf7[1435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1436]),
        .S(self_sf7[1436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1437]),
        .S(self_sf7[1437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1438]),
        .S(self_sf7[1438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1439]),
        .S(self_sf7[1439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[143]),
        .S(self_sf7[143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1440]),
        .S(self_sf7[1440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1441]),
        .S(self_sf7[1441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1442]),
        .S(self_sf7[1442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1443]),
        .S(self_sf7[1443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1444]),
        .S(self_sf7[1444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1445]),
        .S(self_sf7[1445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1446]),
        .S(self_sf7[1446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1447]),
        .S(self_sf7[1447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1448]),
        .S(self_sf7[1448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1449]),
        .S(self_sf7[1449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[144]),
        .S(self_sf7[144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1450]),
        .S(self_sf7[1450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1451]),
        .S(self_sf7[1451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1452]),
        .S(self_sf7[1452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1453]),
        .S(self_sf7[1453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1454]),
        .S(self_sf7[1454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1455]),
        .S(self_sf7[1455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1456]),
        .S(self_sf7[1456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1457]),
        .S(self_sf7[1457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1458]),
        .S(self_sf7[1458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1459]),
        .S(self_sf7[1459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[145]),
        .S(self_sf7[145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1460]),
        .S(self_sf7[1460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1461]),
        .S(self_sf7[1461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1462]),
        .S(self_sf7[1462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1463]),
        .S(self_sf7[1463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1464]),
        .S(self_sf7[1464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1465]),
        .S(self_sf7[1465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1466]),
        .S(self_sf7[1466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1467]),
        .S(self_sf7[1467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1468]),
        .S(self_sf7[1468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1469]),
        .S(self_sf7[1469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[146]),
        .S(self_sf7[146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1470]),
        .S(self_sf7[1470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1471]),
        .S(self_sf7[1471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1472]),
        .S(self_sf7[1472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1473]),
        .S(self_sf7[1473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1474]),
        .S(self_sf7[1474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1475]),
        .S(self_sf7[1475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1476]),
        .S(self_sf7[1476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1477]),
        .S(self_sf7[1477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1478]),
        .S(self_sf7[1478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1479]),
        .S(self_sf7[1479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[147]),
        .S(self_sf7[147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1480]),
        .S(self_sf7[1480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1481]),
        .S(self_sf7[1481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1482]),
        .S(self_sf7[1482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1483]),
        .S(self_sf7[1483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1484]),
        .S(self_sf7[1484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1485]),
        .S(self_sf7[1485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1486]),
        .S(self_sf7[1486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1487]),
        .S(self_sf7[1487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1488]),
        .S(self_sf7[1488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1489]),
        .S(self_sf7[1489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[148]),
        .S(self_sf7[148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1490]),
        .S(self_sf7[1490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1491]),
        .S(self_sf7[1491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1492]),
        .S(self_sf7[1492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1493]),
        .S(self_sf7[1493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1494]),
        .S(self_sf7[1494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1495]),
        .S(self_sf7[1495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1496]),
        .S(self_sf7[1496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1497]),
        .S(self_sf7[1497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1498]),
        .S(self_sf7[1498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1499]),
        .S(self_sf7[1499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[149]),
        .S(self_sf7[149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[14].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[14]),
        .S(self_sf7[14]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1500]),
        .S(self_sf7[1500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1501]),
        .S(self_sf7[1501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1502]),
        .S(self_sf7[1502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1503]),
        .S(self_sf7[1503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1504]),
        .S(self_sf7[1504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1505]),
        .S(self_sf7[1505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1506]),
        .S(self_sf7[1506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1507]),
        .S(self_sf7[1507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1508]),
        .S(self_sf7[1508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1509]),
        .S(self_sf7[1509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[150]),
        .S(self_sf7[150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1510]),
        .S(self_sf7[1510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1511]),
        .S(self_sf7[1511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1512]),
        .S(self_sf7[1512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1513]),
        .S(self_sf7[1513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1514]),
        .S(self_sf7[1514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1515]),
        .S(self_sf7[1515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1516]),
        .S(self_sf7[1516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1517]),
        .S(self_sf7[1517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1518]),
        .S(self_sf7[1518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1519]),
        .S(self_sf7[1519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[151]),
        .S(self_sf7[151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1520]),
        .S(self_sf7[1520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1521]),
        .S(self_sf7[1521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1522]),
        .S(self_sf7[1522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1523]),
        .S(self_sf7[1523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1524]),
        .S(self_sf7[1524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1525]),
        .S(self_sf7[1525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1526]),
        .S(self_sf7[1526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1527]),
        .S(self_sf7[1527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1528]),
        .S(self_sf7[1528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1529]),
        .S(self_sf7[1529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[152]),
        .S(self_sf7[152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1530]),
        .S(self_sf7[1530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1531]),
        .S(self_sf7[1531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1532]),
        .S(self_sf7[1532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1533]),
        .S(self_sf7[1533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1534]),
        .S(self_sf7[1534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1535]),
        .S(self_sf7[1535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1536]),
        .S(self_sf7[1536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1537]),
        .S(self_sf7[1537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1538]),
        .S(self_sf7[1538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1539]),
        .S(self_sf7[1539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[153]),
        .S(self_sf7[153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1540]),
        .S(self_sf7[1540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1541]),
        .S(self_sf7[1541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1542]),
        .S(self_sf7[1542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1543]),
        .S(self_sf7[1543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1544]),
        .S(self_sf7[1544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1545]),
        .S(self_sf7[1545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1546]),
        .S(self_sf7[1546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1547]),
        .S(self_sf7[1547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1548]),
        .S(self_sf7[1548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1549]),
        .S(self_sf7[1549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[154]),
        .S(self_sf7[154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1550]),
        .S(self_sf7[1550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1551]),
        .S(self_sf7[1551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1552]),
        .S(self_sf7[1552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1553]),
        .S(self_sf7[1553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1554]),
        .S(self_sf7[1554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1555]),
        .S(self_sf7[1555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1556]),
        .S(self_sf7[1556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1557]),
        .S(self_sf7[1557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1558]),
        .S(self_sf7[1558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1559]),
        .S(self_sf7[1559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[155]),
        .S(self_sf7[155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1560]),
        .S(self_sf7[1560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1561]),
        .S(self_sf7[1561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1562]),
        .S(self_sf7[1562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1563]),
        .S(self_sf7[1563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1564]),
        .S(self_sf7[1564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1565]),
        .S(self_sf7[1565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1566]),
        .S(self_sf7[1566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1567]),
        .S(self_sf7[1567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1568]),
        .S(self_sf7[1568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1569]),
        .S(self_sf7[1569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[156]),
        .S(self_sf7[156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1570]),
        .S(self_sf7[1570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1571]),
        .S(self_sf7[1571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1572]),
        .S(self_sf7[1572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1573]),
        .S(self_sf7[1573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1574]),
        .S(self_sf7[1574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1575]),
        .S(self_sf7[1575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1576]),
        .S(self_sf7[1576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1577]),
        .S(self_sf7[1577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1578]),
        .S(self_sf7[1578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1579]),
        .S(self_sf7[1579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[157]),
        .S(self_sf7[157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1580]),
        .S(self_sf7[1580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1581]),
        .S(self_sf7[1581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1582]),
        .S(self_sf7[1582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1583]),
        .S(self_sf7[1583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1584]),
        .S(self_sf7[1584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1585]),
        .S(self_sf7[1585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1586]),
        .S(self_sf7[1586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1587]),
        .S(self_sf7[1587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1588]),
        .S(self_sf7[1588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1589]),
        .S(self_sf7[1589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[158]),
        .S(self_sf7[158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1590]),
        .S(self_sf7[1590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1591]),
        .S(self_sf7[1591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1592]),
        .S(self_sf7[1592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1593]),
        .S(self_sf7[1593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1594]),
        .S(self_sf7[1594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1595]),
        .S(self_sf7[1595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1596]),
        .S(self_sf7[1596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1597]),
        .S(self_sf7[1597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1598]),
        .S(self_sf7[1598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1599]),
        .S(self_sf7[1599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[159]),
        .S(self_sf7[159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[15].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[15]),
        .S(self_sf7[15]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1600]),
        .S(self_sf7[1600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1601]),
        .S(self_sf7[1601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1602]),
        .S(self_sf7[1602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1603]),
        .S(self_sf7[1603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1604]),
        .S(self_sf7[1604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1605]),
        .S(self_sf7[1605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1606]),
        .S(self_sf7[1606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1607]),
        .S(self_sf7[1607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1608]),
        .S(self_sf7[1608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1609]),
        .S(self_sf7[1609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[160]),
        .S(self_sf7[160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1610]),
        .S(self_sf7[1610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1611]),
        .S(self_sf7[1611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1612]),
        .S(self_sf7[1612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1613]),
        .S(self_sf7[1613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1614]),
        .S(self_sf7[1614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1615]),
        .S(self_sf7[1615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1616]),
        .S(self_sf7[1616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1617]),
        .S(self_sf7[1617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1618]),
        .S(self_sf7[1618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1619]),
        .S(self_sf7[1619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[161]),
        .S(self_sf7[161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1620]),
        .S(self_sf7[1620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1621]),
        .S(self_sf7[1621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1622]),
        .S(self_sf7[1622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1623]),
        .S(self_sf7[1623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1624]),
        .S(self_sf7[1624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1625]),
        .S(self_sf7[1625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1626]),
        .S(self_sf7[1626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1627]),
        .S(self_sf7[1627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1628]),
        .S(self_sf7[1628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1629]),
        .S(self_sf7[1629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[162]),
        .S(self_sf7[162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1630]),
        .S(self_sf7[1630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1631]),
        .S(self_sf7[1631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1632]),
        .S(self_sf7[1632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1633]),
        .S(self_sf7[1633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1634]),
        .S(self_sf7[1634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1635]),
        .S(self_sf7[1635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1636]),
        .S(self_sf7[1636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1637]),
        .S(self_sf7[1637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1638]),
        .S(self_sf7[1638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1639]),
        .S(self_sf7[1639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[163]),
        .S(self_sf7[163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1640]),
        .S(self_sf7[1640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1641]),
        .S(self_sf7[1641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1642]),
        .S(self_sf7[1642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1643]),
        .S(self_sf7[1643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1644]),
        .S(self_sf7[1644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1645]),
        .S(self_sf7[1645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1646]),
        .S(self_sf7[1646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1647]),
        .S(self_sf7[1647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1648]),
        .S(self_sf7[1648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1649]),
        .S(self_sf7[1649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[164]),
        .S(self_sf7[164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1650]),
        .S(self_sf7[1650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1651]),
        .S(self_sf7[1651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1652]),
        .S(self_sf7[1652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1653]),
        .S(self_sf7[1653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1654]),
        .S(self_sf7[1654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1655]),
        .S(self_sf7[1655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1656]),
        .S(self_sf7[1656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1657]),
        .S(self_sf7[1657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1658]),
        .S(self_sf7[1658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1659]),
        .S(self_sf7[1659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[165]),
        .S(self_sf7[165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1660]),
        .S(self_sf7[1660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1661]),
        .S(self_sf7[1661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1662]),
        .S(self_sf7[1662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1663]),
        .S(self_sf7[1663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1664]),
        .S(self_sf7[1664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1665]),
        .S(self_sf7[1665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1666]),
        .S(self_sf7[1666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1667]),
        .S(self_sf7[1667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1668]),
        .S(self_sf7[1668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1669]),
        .S(self_sf7[1669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[166]),
        .S(self_sf7[166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1670]),
        .S(self_sf7[1670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1671]),
        .S(self_sf7[1671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1672]),
        .S(self_sf7[1672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1673]),
        .S(self_sf7[1673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1674]),
        .S(self_sf7[1674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1675]),
        .S(self_sf7[1675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1676]),
        .S(self_sf7[1676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1677]),
        .S(self_sf7[1677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1678]),
        .S(self_sf7[1678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1679]),
        .S(self_sf7[1679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[167]),
        .S(self_sf7[167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1680]),
        .S(self_sf7[1680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1681]),
        .S(self_sf7[1681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1682]),
        .S(self_sf7[1682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1683]),
        .S(self_sf7[1683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1684]),
        .S(self_sf7[1684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1685]),
        .S(self_sf7[1685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1686]),
        .S(self_sf7[1686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1687]),
        .S(self_sf7[1687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1688]),
        .S(self_sf7[1688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1689]),
        .S(self_sf7[1689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[168]),
        .S(self_sf7[168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1690]),
        .S(self_sf7[1690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1691]),
        .S(self_sf7[1691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1692]),
        .S(self_sf7[1692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1693]),
        .S(self_sf7[1693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1694]),
        .S(self_sf7[1694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1695]),
        .S(self_sf7[1695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1696]),
        .S(self_sf7[1696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1697]),
        .S(self_sf7[1697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1698]),
        .S(self_sf7[1698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1699]),
        .S(self_sf7[1699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[169]),
        .S(self_sf7[169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[16].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[16]),
        .S(self_sf7[16]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1700]),
        .S(self_sf7[1700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1701]),
        .S(self_sf7[1701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1702]),
        .S(self_sf7[1702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1703]),
        .S(self_sf7[1703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1704]),
        .S(self_sf7[1704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1705]),
        .S(self_sf7[1705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1706]),
        .S(self_sf7[1706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1707]),
        .S(self_sf7[1707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1708]),
        .S(self_sf7[1708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1709]),
        .S(self_sf7[1709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[170]),
        .S(self_sf7[170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1710]),
        .S(self_sf7[1710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1711]),
        .S(self_sf7[1711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1712]),
        .S(self_sf7[1712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1713]),
        .S(self_sf7[1713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1714]),
        .S(self_sf7[1714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1715]),
        .S(self_sf7[1715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1716]),
        .S(self_sf7[1716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1717]),
        .S(self_sf7[1717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1718]),
        .S(self_sf7[1718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1719]),
        .S(self_sf7[1719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[171]),
        .S(self_sf7[171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1720]),
        .S(self_sf7[1720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1721]),
        .S(self_sf7[1721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1722]),
        .S(self_sf7[1722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1723]),
        .S(self_sf7[1723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1724]),
        .S(self_sf7[1724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1725]),
        .S(self_sf7[1725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1726]),
        .S(self_sf7[1726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1727]),
        .S(self_sf7[1727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1728]),
        .S(self_sf7[1728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1729]),
        .S(self_sf7[1729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[172]),
        .S(self_sf7[172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1730]),
        .S(self_sf7[1730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1731]),
        .S(self_sf7[1731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1732]),
        .S(self_sf7[1732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1733]),
        .S(self_sf7[1733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1734]),
        .S(self_sf7[1734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1735]),
        .S(self_sf7[1735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1736]),
        .S(self_sf7[1736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1737]),
        .S(self_sf7[1737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1738]),
        .S(self_sf7[1738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1739]),
        .S(self_sf7[1739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[173]),
        .S(self_sf7[173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1740]),
        .S(self_sf7[1740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1741]),
        .S(self_sf7[1741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1742]),
        .S(self_sf7[1742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1743]),
        .S(self_sf7[1743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1744]),
        .S(self_sf7[1744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1745]),
        .S(self_sf7[1745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1746]),
        .S(self_sf7[1746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1747]),
        .S(self_sf7[1747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1748]),
        .S(self_sf7[1748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1749]),
        .S(self_sf7[1749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[174]),
        .S(self_sf7[174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1750]),
        .S(self_sf7[1750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1751]),
        .S(self_sf7[1751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1752]),
        .S(self_sf7[1752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1753]),
        .S(self_sf7[1753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1754]),
        .S(self_sf7[1754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1755]),
        .S(self_sf7[1755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1756]),
        .S(self_sf7[1756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1757]),
        .S(self_sf7[1757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1758]),
        .S(self_sf7[1758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1759]),
        .S(self_sf7[1759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[175]),
        .S(self_sf7[175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1760]),
        .S(self_sf7[1760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1761]),
        .S(self_sf7[1761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1762]),
        .S(self_sf7[1762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1763]),
        .S(self_sf7[1763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1764]),
        .S(self_sf7[1764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1765]),
        .S(self_sf7[1765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1766]),
        .S(self_sf7[1766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1767]),
        .S(self_sf7[1767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1768]),
        .S(self_sf7[1768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1769]),
        .S(self_sf7[1769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[176]),
        .S(self_sf7[176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1770]),
        .S(self_sf7[1770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1771]),
        .S(self_sf7[1771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1772]),
        .S(self_sf7[1772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1773]),
        .S(self_sf7[1773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1774]),
        .S(self_sf7[1774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1775]),
        .S(self_sf7[1775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1776]),
        .S(self_sf7[1776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1777]),
        .S(self_sf7[1777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1778]),
        .S(self_sf7[1778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1779]),
        .S(self_sf7[1779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[177]),
        .S(self_sf7[177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1780]),
        .S(self_sf7[1780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1781]),
        .S(self_sf7[1781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1782]),
        .S(self_sf7[1782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1783]),
        .S(self_sf7[1783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1784]),
        .S(self_sf7[1784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1785]),
        .S(self_sf7[1785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1786]),
        .S(self_sf7[1786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1787]),
        .S(self_sf7[1787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1788]),
        .S(self_sf7[1788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1789]),
        .S(self_sf7[1789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[178]),
        .S(self_sf7[178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1790]),
        .S(self_sf7[1790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1791]),
        .S(self_sf7[1791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1792]),
        .S(self_sf7[1792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1793]),
        .S(self_sf7[1793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1794]),
        .S(self_sf7[1794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1795]),
        .S(self_sf7[1795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1796]),
        .S(self_sf7[1796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1797]),
        .S(self_sf7[1797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1798]),
        .S(self_sf7[1798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1799]),
        .S(self_sf7[1799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[179]),
        .S(self_sf7[179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[17].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[17]),
        .S(self_sf7[17]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[180]),
        .S(self_sf7[180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[181]),
        .S(self_sf7[181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[182]),
        .S(self_sf7[182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[183]),
        .S(self_sf7[183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[184]),
        .S(self_sf7[184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[185]),
        .S(self_sf7[185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[186]),
        .S(self_sf7[186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[187]),
        .S(self_sf7[187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[188]),
        .S(self_sf7[188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[189]),
        .S(self_sf7[189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[18].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[18]),
        .S(self_sf7[18]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[190]),
        .S(self_sf7[190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[191]),
        .S(self_sf7[191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[192]),
        .S(self_sf7[192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[193]),
        .S(self_sf7[193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[194]),
        .S(self_sf7[194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[195]),
        .S(self_sf7[195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[196]),
        .S(self_sf7[196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[197]),
        .S(self_sf7[197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[198]),
        .S(self_sf7[198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[199]),
        .S(self_sf7[199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[19].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[19]),
        .S(self_sf7[19]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1]),
        .S(info_sf7[1]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[200]),
        .S(self_sf7[200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[201]),
        .S(self_sf7[201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[202]),
        .S(self_sf7[202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[203]),
        .S(self_sf7[203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[204]),
        .S(self_sf7[204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[205]),
        .S(self_sf7[205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[206]),
        .S(self_sf7[206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[207]),
        .S(self_sf7[207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[208]),
        .S(self_sf7[208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[209]),
        .S(self_sf7[209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[20].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[20]),
        .S(self_sf7[20]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[210]),
        .S(self_sf7[210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[211]),
        .S(self_sf7[211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[212]),
        .S(self_sf7[212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[213]),
        .S(self_sf7[213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[214]),
        .S(self_sf7[214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[215]),
        .S(self_sf7[215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[216]),
        .S(self_sf7[216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[217]),
        .S(self_sf7[217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[218]),
        .S(self_sf7[218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[219]),
        .S(self_sf7[219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[21].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[21]),
        .S(self_sf7[21]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[220]),
        .S(self_sf7[220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[221]),
        .S(self_sf7[221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[222]),
        .S(self_sf7[222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[223]),
        .S(self_sf7[223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[224]),
        .S(self_sf7[224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[225]),
        .S(self_sf7[225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[226]),
        .S(self_sf7[226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[227]),
        .S(self_sf7[227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[228]),
        .S(self_sf7[228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[229]),
        .S(self_sf7[229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[22].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[22]),
        .S(self_sf7[22]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[230]),
        .S(self_sf7[230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[231]),
        .S(self_sf7[231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[232]),
        .S(self_sf7[232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[233]),
        .S(self_sf7[233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[234]),
        .S(self_sf7[234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[235]),
        .S(self_sf7[235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[236]),
        .S(self_sf7[236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[237]),
        .S(self_sf7[237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[238]),
        .S(self_sf7[238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[239]),
        .S(self_sf7[239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[23].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[23]),
        .S(self_sf7[23]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[240]),
        .S(self_sf7[240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[241]),
        .S(self_sf7[241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[242]),
        .S(self_sf7[242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[243]),
        .S(self_sf7[243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[244]),
        .S(self_sf7[244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[245]),
        .S(self_sf7[245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[246]),
        .S(self_sf7[246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[247]),
        .S(self_sf7[247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[248]),
        .S(self_sf7[248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[249]),
        .S(self_sf7[249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[24].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[24]),
        .S(self_sf7[24]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[250]),
        .S(self_sf7[250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[251]),
        .S(self_sf7[251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[252]),
        .S(self_sf7[252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[253]),
        .S(self_sf7[253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[254]),
        .S(self_sf7[254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[255]),
        .S(self_sf7[255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[256]),
        .S(self_sf7[256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[257]),
        .S(self_sf7[257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[258]),
        .S(self_sf7[258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[259]),
        .S(self_sf7[259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[25].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[25]),
        .S(self_sf7[25]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[260]),
        .S(self_sf7[260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[261]),
        .S(self_sf7[261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[262]),
        .S(self_sf7[262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[263]),
        .S(self_sf7[263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[264]),
        .S(self_sf7[264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[265]),
        .S(self_sf7[265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[266]),
        .S(self_sf7[266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[267]),
        .S(self_sf7[267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[268]),
        .S(self_sf7[268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[269]),
        .S(self_sf7[269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[26].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[26]),
        .S(self_sf7[26]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[270]),
        .S(self_sf7[270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[271]),
        .S(self_sf7[271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[272]),
        .S(self_sf7[272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[273]),
        .S(self_sf7[273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[274]),
        .S(self_sf7[274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[275]),
        .S(self_sf7[275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[276]),
        .S(self_sf7[276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[277]),
        .S(self_sf7[277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[278]),
        .S(self_sf7[278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[279]),
        .S(self_sf7[279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[27].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[27]),
        .S(self_sf7[27]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[280]),
        .S(self_sf7[280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[281]),
        .S(self_sf7[281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[282]),
        .S(self_sf7[282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[283]),
        .S(self_sf7[283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[284]),
        .S(self_sf7[284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[285]),
        .S(self_sf7[285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[286]),
        .S(self_sf7[286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[287]),
        .S(self_sf7[287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[288]),
        .S(self_sf7[288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[289]),
        .S(self_sf7[289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[28].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[28]),
        .S(self_sf7[28]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[290]),
        .S(self_sf7[290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[291]),
        .S(self_sf7[291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[292]),
        .S(self_sf7[292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[293]),
        .S(self_sf7[293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[294]),
        .S(self_sf7[294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[295]),
        .S(self_sf7[295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[296]),
        .S(self_sf7[296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[297]),
        .S(self_sf7[297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[298]),
        .S(self_sf7[298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[299]),
        .S(self_sf7[299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[29].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[29]),
        .S(self_sf7[29]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[2].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[2]),
        .S(info_sf7[2]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[300]),
        .S(self_sf7[300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[301]),
        .S(self_sf7[301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[302]),
        .S(self_sf7[302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[303]),
        .S(self_sf7[303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[304]),
        .S(self_sf7[304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[305]),
        .S(self_sf7[305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[306]),
        .S(self_sf7[306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[307]),
        .S(self_sf7[307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[308]),
        .S(self_sf7[308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[309]),
        .S(self_sf7[309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[30].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[30]),
        .S(self_sf7[30]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[310]),
        .S(self_sf7[310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[311]),
        .S(self_sf7[311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[312]),
        .S(self_sf7[312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[313]),
        .S(self_sf7[313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[314]),
        .S(self_sf7[314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[315]),
        .S(self_sf7[315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[316]),
        .S(self_sf7[316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[317]),
        .S(self_sf7[317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[318]),
        .S(self_sf7[318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[319]),
        .S(self_sf7[319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[31].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[31]),
        .S(self_sf7[31]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[320]),
        .S(self_sf7[320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[321]),
        .S(self_sf7[321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[322]),
        .S(self_sf7[322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[323]),
        .S(self_sf7[323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[324]),
        .S(self_sf7[324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[325]),
        .S(self_sf7[325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[326]),
        .S(self_sf7[326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[327]),
        .S(self_sf7[327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[328]),
        .S(self_sf7[328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[329]),
        .S(self_sf7[329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[32].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[32]),
        .S(self_sf7[32]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[330]),
        .S(self_sf7[330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[331]),
        .S(self_sf7[331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[332]),
        .S(self_sf7[332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[333]),
        .S(self_sf7[333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[334]),
        .S(self_sf7[334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[335]),
        .S(self_sf7[335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[336]),
        .S(self_sf7[336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[337]),
        .S(self_sf7[337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[338]),
        .S(self_sf7[338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[339]),
        .S(self_sf7[339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[33].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[33]),
        .S(self_sf7[33]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[340]),
        .S(self_sf7[340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[341]),
        .S(self_sf7[341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[342]),
        .S(self_sf7[342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[343]),
        .S(self_sf7[343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[344]),
        .S(self_sf7[344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[345]),
        .S(self_sf7[345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[346]),
        .S(self_sf7[346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[347]),
        .S(self_sf7[347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[348]),
        .S(self_sf7[348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[349]),
        .S(self_sf7[349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[34].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[34]),
        .S(self_sf7[34]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[350]),
        .S(self_sf7[350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[351]),
        .S(self_sf7[351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[352]),
        .S(self_sf7[352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[353]),
        .S(self_sf7[353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[354]),
        .S(self_sf7[354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[355]),
        .S(self_sf7[355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[356]),
        .S(self_sf7[356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[357]),
        .S(self_sf7[357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[358]),
        .S(self_sf7[358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[359]),
        .S(self_sf7[359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[35].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[35]),
        .S(self_sf7[35]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[360]),
        .S(self_sf7[360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[361]),
        .S(self_sf7[361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[362]),
        .S(self_sf7[362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[363]),
        .S(self_sf7[363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[364]),
        .S(self_sf7[364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[365]),
        .S(self_sf7[365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[366]),
        .S(self_sf7[366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[367]),
        .S(self_sf7[367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[368]),
        .S(self_sf7[368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[369]),
        .S(self_sf7[369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[36].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[36]),
        .S(self_sf7[36]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[370]),
        .S(self_sf7[370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[371]),
        .S(self_sf7[371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[372]),
        .S(self_sf7[372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[373]),
        .S(self_sf7[373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[374]),
        .S(self_sf7[374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[375]),
        .S(self_sf7[375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[376]),
        .S(self_sf7[376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[377]),
        .S(self_sf7[377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[378]),
        .S(self_sf7[378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[379]),
        .S(self_sf7[379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[37].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[37]),
        .S(self_sf7[37]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[380]),
        .S(self_sf7[380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[381]),
        .S(self_sf7[381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[382]),
        .S(self_sf7[382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[383]),
        .S(self_sf7[383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[384]),
        .S(self_sf7[384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[385]),
        .S(self_sf7[385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[386]),
        .S(self_sf7[386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[387]),
        .S(self_sf7[387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[388]),
        .S(self_sf7[388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[389]),
        .S(self_sf7[389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[38].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[38]),
        .S(self_sf7[38]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[390]),
        .S(self_sf7[390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[391]),
        .S(self_sf7[391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[392]),
        .S(self_sf7[392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[393]),
        .S(self_sf7[393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[394]),
        .S(self_sf7[394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[395]),
        .S(self_sf7[395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[396]),
        .S(self_sf7[396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[397]),
        .S(self_sf7[397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[398]),
        .S(self_sf7[398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[399]),
        .S(self_sf7[399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[39].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[39]),
        .S(self_sf7[39]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[3].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[3]),
        .S(info_sf7[3]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[400]),
        .S(self_sf7[400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[401]),
        .S(self_sf7[401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[402]),
        .S(self_sf7[402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[403]),
        .S(self_sf7[403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[404]),
        .S(self_sf7[404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[405]),
        .S(self_sf7[405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[406]),
        .S(self_sf7[406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[407]),
        .S(self_sf7[407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[408]),
        .S(self_sf7[408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[409]),
        .S(self_sf7[409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[40].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[40]),
        .S(self_sf7[40]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[410]),
        .S(self_sf7[410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[411]),
        .S(self_sf7[411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[412]),
        .S(self_sf7[412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[413]),
        .S(self_sf7[413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[414]),
        .S(self_sf7[414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[415]),
        .S(self_sf7[415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[416]),
        .S(self_sf7[416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[417]),
        .S(self_sf7[417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[418]),
        .S(self_sf7[418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[419]),
        .S(self_sf7[419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[41].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[41]),
        .S(self_sf7[41]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[420]),
        .S(self_sf7[420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[421]),
        .S(self_sf7[421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[422]),
        .S(self_sf7[422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[423]),
        .S(self_sf7[423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[424]),
        .S(self_sf7[424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[425]),
        .S(self_sf7[425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[426]),
        .S(self_sf7[426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[427]),
        .S(self_sf7[427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[428]),
        .S(self_sf7[428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[429]),
        .S(self_sf7[429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[42].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[42]),
        .S(self_sf7[42]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[430]),
        .S(self_sf7[430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[431]),
        .S(self_sf7[431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[432]),
        .S(self_sf7[432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[433]),
        .S(self_sf7[433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[434]),
        .S(self_sf7[434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[435]),
        .S(self_sf7[435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[436]),
        .S(self_sf7[436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[437]),
        .S(self_sf7[437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[438]),
        .S(self_sf7[438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[439]),
        .S(self_sf7[439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[43].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[43]),
        .S(self_sf7[43]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[440]),
        .S(self_sf7[440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[441]),
        .S(self_sf7[441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[442]),
        .S(self_sf7[442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[443]),
        .S(self_sf7[443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[444]),
        .S(self_sf7[444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[445]),
        .S(self_sf7[445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[446]),
        .S(self_sf7[446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[447]),
        .S(self_sf7[447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[448]),
        .S(self_sf7[448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[449]),
        .S(self_sf7[449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[44].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[44]),
        .S(self_sf7[44]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[450]),
        .S(self_sf7[450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[451]),
        .S(self_sf7[451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[452]),
        .S(self_sf7[452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[453]),
        .S(self_sf7[453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[454]),
        .S(self_sf7[454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[455]),
        .S(self_sf7[455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[456]),
        .S(self_sf7[456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[457]),
        .S(self_sf7[457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[458]),
        .S(self_sf7[458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[459]),
        .S(self_sf7[459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[45].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[45]),
        .S(self_sf7[45]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[460]),
        .S(self_sf7[460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[461]),
        .S(self_sf7[461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[462]),
        .S(self_sf7[462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[463]),
        .S(self_sf7[463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[464]),
        .S(self_sf7[464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[465]),
        .S(self_sf7[465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[466]),
        .S(self_sf7[466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[467]),
        .S(self_sf7[467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[468]),
        .S(self_sf7[468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[469]),
        .S(self_sf7[469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[46].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[46]),
        .S(self_sf7[46]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[470]),
        .S(self_sf7[470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[471]),
        .S(self_sf7[471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[472]),
        .S(self_sf7[472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[473]),
        .S(self_sf7[473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[474]),
        .S(self_sf7[474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[475]),
        .S(self_sf7[475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[476]),
        .S(self_sf7[476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[477]),
        .S(self_sf7[477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[478]),
        .S(self_sf7[478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[479]),
        .S(self_sf7[479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[47].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[47]),
        .S(self_sf7[47]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[480]),
        .S(self_sf7[480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[481]),
        .S(self_sf7[481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[482]),
        .S(self_sf7[482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[483]),
        .S(self_sf7[483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[484]),
        .S(self_sf7[484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[485]),
        .S(self_sf7[485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[486]),
        .S(self_sf7[486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[487]),
        .S(self_sf7[487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[488]),
        .S(self_sf7[488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[489]),
        .S(self_sf7[489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[48].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[48]),
        .S(self_sf7[48]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[490]),
        .S(self_sf7[490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[491]),
        .S(self_sf7[491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[492]),
        .S(self_sf7[492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[493]),
        .S(self_sf7[493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[494]),
        .S(self_sf7[494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[495]),
        .S(self_sf7[495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[496]),
        .S(self_sf7[496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[497]),
        .S(self_sf7[497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[498]),
        .S(self_sf7[498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[499]),
        .S(self_sf7[499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[49].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[49]),
        .S(self_sf7[49]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[4].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[4]),
        .S(info_sf7[4]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[500]),
        .S(self_sf7[500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[501]),
        .S(self_sf7[501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[502]),
        .S(self_sf7[502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[503]),
        .S(self_sf7[503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[504]),
        .S(self_sf7[504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[505]),
        .S(self_sf7[505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[506]),
        .S(self_sf7[506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[507]),
        .S(self_sf7[507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[508]),
        .S(self_sf7[508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[509]),
        .S(self_sf7[509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[50].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[50]),
        .S(self_sf7[50]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[510]),
        .S(self_sf7[510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[511]),
        .S(self_sf7[511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[512]),
        .S(self_sf7[512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[513]),
        .S(self_sf7[513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[514]),
        .S(self_sf7[514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[515]),
        .S(self_sf7[515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[516]),
        .S(self_sf7[516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[517]),
        .S(self_sf7[517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[518]),
        .S(self_sf7[518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[519]),
        .S(self_sf7[519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[51].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[51]),
        .S(self_sf7[51]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[520]),
        .S(self_sf7[520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[521]),
        .S(self_sf7[521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[522]),
        .S(self_sf7[522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[523]),
        .S(self_sf7[523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[524]),
        .S(self_sf7[524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[525]),
        .S(self_sf7[525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[526]),
        .S(self_sf7[526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[527]),
        .S(self_sf7[527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[528]),
        .S(self_sf7[528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[529]),
        .S(self_sf7[529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[52].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[52]),
        .S(self_sf7[52]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[530]),
        .S(self_sf7[530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[531]),
        .S(self_sf7[531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[532]),
        .S(self_sf7[532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[533]),
        .S(self_sf7[533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[534]),
        .S(self_sf7[534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[535]),
        .S(self_sf7[535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[536]),
        .S(self_sf7[536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[537]),
        .S(self_sf7[537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[538]),
        .S(self_sf7[538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[539]),
        .S(self_sf7[539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[53].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[53]),
        .S(self_sf7[53]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[540]),
        .S(self_sf7[540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[541]),
        .S(self_sf7[541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[542]),
        .S(self_sf7[542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[543]),
        .S(self_sf7[543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[544]),
        .S(self_sf7[544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[545]),
        .S(self_sf7[545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[546]),
        .S(self_sf7[546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[547]),
        .S(self_sf7[547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[548]),
        .S(self_sf7[548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[549]),
        .S(self_sf7[549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[54].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[54]),
        .S(self_sf7[54]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[550]),
        .S(self_sf7[550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[551]),
        .S(self_sf7[551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[552]),
        .S(self_sf7[552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[553]),
        .S(self_sf7[553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[554]),
        .S(self_sf7[554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[555]),
        .S(self_sf7[555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[556]),
        .S(self_sf7[556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[557]),
        .S(self_sf7[557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[558]),
        .S(self_sf7[558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[559]),
        .S(self_sf7[559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[55].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[55]),
        .S(self_sf7[55]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[560]),
        .S(self_sf7[560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[561]),
        .S(self_sf7[561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[562]),
        .S(self_sf7[562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[563]),
        .S(self_sf7[563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[564]),
        .S(self_sf7[564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[565]),
        .S(self_sf7[565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[566]),
        .S(self_sf7[566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[567]),
        .S(self_sf7[567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[568]),
        .S(self_sf7[568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[569]),
        .S(self_sf7[569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[56].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[56]),
        .S(self_sf7[56]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[570]),
        .S(self_sf7[570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[571]),
        .S(self_sf7[571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[572]),
        .S(self_sf7[572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[573]),
        .S(self_sf7[573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[574]),
        .S(self_sf7[574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[575]),
        .S(self_sf7[575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[576]),
        .S(self_sf7[576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[577]),
        .S(self_sf7[577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[578]),
        .S(self_sf7[578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[579]),
        .S(self_sf7[579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[57].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[57]),
        .S(self_sf7[57]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[580]),
        .S(self_sf7[580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[581]),
        .S(self_sf7[581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[582]),
        .S(self_sf7[582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[583]),
        .S(self_sf7[583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[584]),
        .S(self_sf7[584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[585]),
        .S(self_sf7[585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[586]),
        .S(self_sf7[586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[587]),
        .S(self_sf7[587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[588]),
        .S(self_sf7[588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[589]),
        .S(self_sf7[589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[58].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[58]),
        .S(self_sf7[58]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[590]),
        .S(self_sf7[590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[591]),
        .S(self_sf7[591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[592]),
        .S(self_sf7[592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[593]),
        .S(self_sf7[593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[594]),
        .S(self_sf7[594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[595]),
        .S(self_sf7[595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[596]),
        .S(self_sf7[596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[597]),
        .S(self_sf7[597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[598]),
        .S(self_sf7[598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[599]),
        .S(self_sf7[599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[59].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[59]),
        .S(self_sf7[59]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[5].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[5]),
        .S(info_sf7[5]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[600]),
        .S(self_sf7[600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[601]),
        .S(self_sf7[601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[602]),
        .S(self_sf7[602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[603]),
        .S(self_sf7[603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[604]),
        .S(self_sf7[604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[605]),
        .S(self_sf7[605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[606]),
        .S(self_sf7[606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[607]),
        .S(self_sf7[607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[608]),
        .S(self_sf7[608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[609]),
        .S(self_sf7[609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[60].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[60]),
        .S(self_sf7[60]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[610]),
        .S(self_sf7[610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[611]),
        .S(self_sf7[611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[612]),
        .S(self_sf7[612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[613]),
        .S(self_sf7[613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[614]),
        .S(self_sf7[614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[615]),
        .S(self_sf7[615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[616]),
        .S(self_sf7[616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[617]),
        .S(self_sf7[617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[618]),
        .S(self_sf7[618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[619]),
        .S(self_sf7[619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[61].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[61]),
        .S(self_sf7[61]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[620]),
        .S(self_sf7[620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[621]),
        .S(self_sf7[621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[622]),
        .S(self_sf7[622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[623]),
        .S(self_sf7[623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[624]),
        .S(self_sf7[624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[625]),
        .S(self_sf7[625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[626]),
        .S(self_sf7[626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[627]),
        .S(self_sf7[627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[628]),
        .S(self_sf7[628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[629]),
        .S(self_sf7[629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[62].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[62]),
        .S(self_sf7[62]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[630]),
        .S(self_sf7[630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[631]),
        .S(self_sf7[631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[632]),
        .S(self_sf7[632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[633]),
        .S(self_sf7[633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[634]),
        .S(self_sf7[634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[635]),
        .S(self_sf7[635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[636]),
        .S(self_sf7[636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[637]),
        .S(self_sf7[637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[638]),
        .S(self_sf7[638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[639]),
        .S(self_sf7[639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[63].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[63]),
        .S(self_sf7[63]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[640]),
        .S(self_sf7[640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[641]),
        .S(self_sf7[641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[642]),
        .S(self_sf7[642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[643]),
        .S(self_sf7[643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[644]),
        .S(self_sf7[644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[645]),
        .S(self_sf7[645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[646]),
        .S(self_sf7[646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[647]),
        .S(self_sf7[647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[648]),
        .S(self_sf7[648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[649]),
        .S(self_sf7[649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[64].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[64]),
        .S(self_sf7[64]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[650]),
        .S(self_sf7[650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[651]),
        .S(self_sf7[651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[652]),
        .S(self_sf7[652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[653]),
        .S(self_sf7[653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[654]),
        .S(self_sf7[654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[655]),
        .S(self_sf7[655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[656]),
        .S(self_sf7[656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[657]),
        .S(self_sf7[657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[658]),
        .S(self_sf7[658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[659]),
        .S(self_sf7[659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[65].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[65]),
        .S(self_sf7[65]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[660]),
        .S(self_sf7[660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[661]),
        .S(self_sf7[661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[662]),
        .S(self_sf7[662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[663]),
        .S(self_sf7[663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[664]),
        .S(self_sf7[664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[665]),
        .S(self_sf7[665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[666]),
        .S(self_sf7[666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[667]),
        .S(self_sf7[667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[668]),
        .S(self_sf7[668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[669]),
        .S(self_sf7[669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[66].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[66]),
        .S(self_sf7[66]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[670]),
        .S(self_sf7[670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[671]),
        .S(self_sf7[671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[672]),
        .S(self_sf7[672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[673]),
        .S(self_sf7[673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[674]),
        .S(self_sf7[674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[675]),
        .S(self_sf7[675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[676]),
        .S(self_sf7[676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[677]),
        .S(self_sf7[677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[678]),
        .S(self_sf7[678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[679]),
        .S(self_sf7[679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[67].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[67]),
        .S(self_sf7[67]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[680]),
        .S(self_sf7[680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[681]),
        .S(self_sf7[681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[682]),
        .S(self_sf7[682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[683]),
        .S(self_sf7[683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[684]),
        .S(self_sf7[684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[685]),
        .S(self_sf7[685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[686]),
        .S(self_sf7[686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[687]),
        .S(self_sf7[687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[688]),
        .S(self_sf7[688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[689]),
        .S(self_sf7[689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[68].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[68]),
        .S(self_sf7[68]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[690]),
        .S(self_sf7[690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[691]),
        .S(self_sf7[691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[692]),
        .S(self_sf7[692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[693]),
        .S(self_sf7[693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[694]),
        .S(self_sf7[694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[695]),
        .S(self_sf7[695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[696]),
        .S(self_sf7[696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[697]),
        .S(self_sf7[697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[698]),
        .S(self_sf7[698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[699]),
        .S(self_sf7[699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[69].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[69]),
        .S(self_sf7[69]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[6].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[6]),
        .S(info_sf7[6]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[700]),
        .S(self_sf7[700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[701]),
        .S(self_sf7[701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[702]),
        .S(self_sf7[702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[703]),
        .S(self_sf7[703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[704]),
        .S(self_sf7[704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[705]),
        .S(self_sf7[705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[706]),
        .S(self_sf7[706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[707]),
        .S(self_sf7[707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[708]),
        .S(self_sf7[708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[709]),
        .S(self_sf7[709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[70].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[70]),
        .S(self_sf7[70]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[710]),
        .S(self_sf7[710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[711]),
        .S(self_sf7[711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[712]),
        .S(self_sf7[712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[713]),
        .S(self_sf7[713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[714]),
        .S(self_sf7[714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[715]),
        .S(self_sf7[715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[716]),
        .S(self_sf7[716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[717]),
        .S(self_sf7[717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[718]),
        .S(self_sf7[718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[719]),
        .S(self_sf7[719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[71].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[71]),
        .S(self_sf7[71]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[720]),
        .S(self_sf7[720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[721]),
        .S(self_sf7[721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[722]),
        .S(self_sf7[722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[723]),
        .S(self_sf7[723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[724]),
        .S(self_sf7[724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[725]),
        .S(self_sf7[725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[726]),
        .S(self_sf7[726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[727]),
        .S(self_sf7[727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[728]),
        .S(self_sf7[728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[729]),
        .S(self_sf7[729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[72].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[72]),
        .S(self_sf7[72]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[730]),
        .S(self_sf7[730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[731]),
        .S(self_sf7[731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[732]),
        .S(self_sf7[732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[733]),
        .S(self_sf7[733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[734]),
        .S(self_sf7[734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[735]),
        .S(self_sf7[735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[736]),
        .S(self_sf7[736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[737]),
        .S(self_sf7[737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[738]),
        .S(self_sf7[738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[739]),
        .S(self_sf7[739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[73].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[73]),
        .S(self_sf7[73]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[740]),
        .S(self_sf7[740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[741]),
        .S(self_sf7[741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[742]),
        .S(self_sf7[742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[743]),
        .S(self_sf7[743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[744]),
        .S(self_sf7[744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[745]),
        .S(self_sf7[745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[746]),
        .S(self_sf7[746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[747]),
        .S(self_sf7[747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[748]),
        .S(self_sf7[748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[749]),
        .S(self_sf7[749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[74].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[74]),
        .S(self_sf7[74]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[750]),
        .S(self_sf7[750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[751]),
        .S(self_sf7[751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[752]),
        .S(self_sf7[752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[753]),
        .S(self_sf7[753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[754]),
        .S(self_sf7[754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[755]),
        .S(self_sf7[755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[756]),
        .S(self_sf7[756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[757]),
        .S(self_sf7[757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[758]),
        .S(self_sf7[758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[759]),
        .S(self_sf7[759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[75].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[75]),
        .S(self_sf7[75]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[760]),
        .S(self_sf7[760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[761]),
        .S(self_sf7[761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[762]),
        .S(self_sf7[762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[763]),
        .S(self_sf7[763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[764]),
        .S(self_sf7[764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[765]),
        .S(self_sf7[765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[766]),
        .S(self_sf7[766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[767]),
        .S(self_sf7[767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[768]),
        .S(self_sf7[768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[769]),
        .S(self_sf7[769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[76].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[76]),
        .S(self_sf7[76]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[770]),
        .S(self_sf7[770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[771]),
        .S(self_sf7[771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[772]),
        .S(self_sf7[772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[773]),
        .S(self_sf7[773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[774]),
        .S(self_sf7[774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[775]),
        .S(self_sf7[775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[776]),
        .S(self_sf7[776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[777]),
        .S(self_sf7[777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[778]),
        .S(self_sf7[778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[779]),
        .S(self_sf7[779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[77].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[77]),
        .S(self_sf7[77]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[780]),
        .S(self_sf7[780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[781]),
        .S(self_sf7[781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[782]),
        .S(self_sf7[782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[783]),
        .S(self_sf7[783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[784]),
        .S(self_sf7[784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[785]),
        .S(self_sf7[785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[786]),
        .S(self_sf7[786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[787]),
        .S(self_sf7[787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[788]),
        .S(self_sf7[788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[789]),
        .S(self_sf7[789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[78].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[78]),
        .S(self_sf7[78]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[790]),
        .S(self_sf7[790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[791]),
        .S(self_sf7[791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[792]),
        .S(self_sf7[792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[793]),
        .S(self_sf7[793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[794]),
        .S(self_sf7[794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[795]),
        .S(self_sf7[795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[796]),
        .S(self_sf7[796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[797]),
        .S(self_sf7[797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[798]),
        .S(self_sf7[798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[799]),
        .S(self_sf7[799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[79].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[79]),
        .S(self_sf7[79]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[7].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[7]),
        .S(info_sf7[7]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[800].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[800]),
        .S(self_sf7[800]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[801].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[801]),
        .S(self_sf7[801]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[802].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[802]),
        .S(self_sf7[802]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[803].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[803]),
        .S(self_sf7[803]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[804].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[804]),
        .S(self_sf7[804]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[805].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[805]),
        .S(self_sf7[805]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[806].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[806]),
        .S(self_sf7[806]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[807].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[807]),
        .S(self_sf7[807]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[808].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[808]),
        .S(self_sf7[808]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[809].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[809]),
        .S(self_sf7[809]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[80].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[80]),
        .S(self_sf7[80]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[810].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[810]),
        .S(self_sf7[810]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[811].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[811]),
        .S(self_sf7[811]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[812].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[812]),
        .S(self_sf7[812]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[813].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[813]),
        .S(self_sf7[813]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[814].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[814]),
        .S(self_sf7[814]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[815].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[815]),
        .S(self_sf7[815]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[816].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[816]),
        .S(self_sf7[816]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[817].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[817]),
        .S(self_sf7[817]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[818].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[818]),
        .S(self_sf7[818]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[819].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[819]),
        .S(self_sf7[819]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[81].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[81]),
        .S(self_sf7[81]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[820].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[820]),
        .S(self_sf7[820]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[821].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[821]),
        .S(self_sf7[821]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[822].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[822]),
        .S(self_sf7[822]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[823].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[823]),
        .S(self_sf7[823]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[824].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[824]),
        .S(self_sf7[824]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[825].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[825]),
        .S(self_sf7[825]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[826].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[826]),
        .S(self_sf7[826]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[827].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[827]),
        .S(self_sf7[827]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[828].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[828]),
        .S(self_sf7[828]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[829].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[829]),
        .S(self_sf7[829]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[82].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[82]),
        .S(self_sf7[82]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[830].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[830]),
        .S(self_sf7[830]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[831].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[831]),
        .S(self_sf7[831]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[832].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[832]),
        .S(self_sf7[832]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[833].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[833]),
        .S(self_sf7[833]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[834].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[834]),
        .S(self_sf7[834]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[835].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[835]),
        .S(self_sf7[835]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[836].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[836]),
        .S(self_sf7[836]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[837].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[837]),
        .S(self_sf7[837]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[838].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[838]),
        .S(self_sf7[838]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[839].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[839]),
        .S(self_sf7[839]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[83].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[83]),
        .S(self_sf7[83]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[840].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[840]),
        .S(self_sf7[840]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[841].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[841]),
        .S(self_sf7[841]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[842].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[842]),
        .S(self_sf7[842]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[843].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[843]),
        .S(self_sf7[843]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[844].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[844]),
        .S(self_sf7[844]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[845].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[845]),
        .S(self_sf7[845]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[846].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[846]),
        .S(self_sf7[846]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[847].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[847]),
        .S(self_sf7[847]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[848].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[848]),
        .S(self_sf7[848]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[849].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[849]),
        .S(self_sf7[849]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[84].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[84]),
        .S(self_sf7[84]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[850].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[850]),
        .S(self_sf7[850]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[851].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[851]),
        .S(self_sf7[851]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[852].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[852]),
        .S(self_sf7[852]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[853].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[853]),
        .S(self_sf7[853]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[854].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[854]),
        .S(self_sf7[854]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[855].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[855]),
        .S(self_sf7[855]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[856].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[856]),
        .S(self_sf7[856]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[857].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[857]),
        .S(self_sf7[857]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[858].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[858]),
        .S(self_sf7[858]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[859].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[859]),
        .S(self_sf7[859]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[85].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[85]),
        .S(self_sf7[85]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[860].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[860]),
        .S(self_sf7[860]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[861].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[861]),
        .S(self_sf7[861]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[862].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[862]),
        .S(self_sf7[862]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[863].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[863]),
        .S(self_sf7[863]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[864].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[864]),
        .S(self_sf7[864]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[865].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[865]),
        .S(self_sf7[865]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[866].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[866]),
        .S(self_sf7[866]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[867].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[867]),
        .S(self_sf7[867]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[868].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[868]),
        .S(self_sf7[868]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[869].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[869]),
        .S(self_sf7[869]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[86].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[86]),
        .S(self_sf7[86]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[870].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[870]),
        .S(self_sf7[870]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[871].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[871]),
        .S(self_sf7[871]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[872].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[872]),
        .S(self_sf7[872]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[873].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[873]),
        .S(self_sf7[873]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[874].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[874]),
        .S(self_sf7[874]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[875].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[875]),
        .S(self_sf7[875]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[876].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[876]),
        .S(self_sf7[876]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[877].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[877]),
        .S(self_sf7[877]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[878].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[878]),
        .S(self_sf7[878]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[879].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[879]),
        .S(self_sf7[879]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[87].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[87]),
        .S(self_sf7[87]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[880].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[880]),
        .S(self_sf7[880]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[881].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[881]),
        .S(self_sf7[881]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[882].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[882]),
        .S(self_sf7[882]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[883].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[883]),
        .S(self_sf7[883]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[884].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[884]),
        .S(self_sf7[884]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[885].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[885]),
        .S(self_sf7[885]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[886].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[886]),
        .S(self_sf7[886]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[887].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[887]),
        .S(self_sf7[887]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[888].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[888]),
        .S(self_sf7[888]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[889].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[889]),
        .S(self_sf7[889]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[88].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[88]),
        .S(self_sf7[88]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[890].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[890]),
        .S(self_sf7[890]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[891].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[891]),
        .S(self_sf7[891]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[892].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[892]),
        .S(self_sf7[892]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[893].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[893]),
        .S(self_sf7[893]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[894].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[894]),
        .S(self_sf7[894]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[895].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[895]),
        .S(self_sf7[895]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[896].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[896]),
        .S(self_sf7[896]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[897].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[897]),
        .S(self_sf7[897]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[898].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[898]),
        .S(self_sf7[898]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[899].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[899]),
        .S(self_sf7[899]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[89].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[89]),
        .S(self_sf7[89]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[8].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[8]),
        .S(self_sf7[8]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[900].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[900]),
        .S(self_sf7[900]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[901].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[901]),
        .S(self_sf7[901]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[902].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[902]),
        .S(self_sf7[902]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[903].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[903]),
        .S(self_sf7[903]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[904].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[904]),
        .S(self_sf7[904]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[905].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[905]),
        .S(self_sf7[905]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[906].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[906]),
        .S(self_sf7[906]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[907].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[907]),
        .S(self_sf7[907]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[908].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[908]),
        .S(self_sf7[908]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[909].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[909]),
        .S(self_sf7[909]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[90].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[90]),
        .S(self_sf7[90]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[910].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[910]),
        .S(self_sf7[910]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[911].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[911]),
        .S(self_sf7[911]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[912].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[912]),
        .S(self_sf7[912]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[913].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[913]),
        .S(self_sf7[913]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[914].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[914]),
        .S(self_sf7[914]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[915].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[915]),
        .S(self_sf7[915]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[916].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[916]),
        .S(self_sf7[916]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[917].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[917]),
        .S(self_sf7[917]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[918].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[918]),
        .S(self_sf7[918]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[919].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[919]),
        .S(self_sf7[919]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[91].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[91]),
        .S(self_sf7[91]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[920].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[920]),
        .S(self_sf7[920]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[921].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[921]),
        .S(self_sf7[921]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[922].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[922]),
        .S(self_sf7[922]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[923].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[923]),
        .S(self_sf7[923]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[924].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[924]),
        .S(self_sf7[924]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[925].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[925]),
        .S(self_sf7[925]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[926].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[926]),
        .S(self_sf7[926]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[927].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[927]),
        .S(self_sf7[927]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[928].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[928]),
        .S(self_sf7[928]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[929].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[929]),
        .S(self_sf7[929]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[92].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[92]),
        .S(self_sf7[92]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[930].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[930]),
        .S(self_sf7[930]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[931].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[931]),
        .S(self_sf7[931]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[932].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[932]),
        .S(self_sf7[932]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[933].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[933]),
        .S(self_sf7[933]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[934].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[934]),
        .S(self_sf7[934]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[935].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[935]),
        .S(self_sf7[935]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[936].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[936]),
        .S(self_sf7[936]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[937].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[937]),
        .S(self_sf7[937]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[938].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[938]),
        .S(self_sf7[938]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[939].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[939]),
        .S(self_sf7[939]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[93].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[93]),
        .S(self_sf7[93]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[940].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[940]),
        .S(self_sf7[940]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[941].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[941]),
        .S(self_sf7[941]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[942].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[942]),
        .S(self_sf7[942]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[943].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[943]),
        .S(self_sf7[943]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[944].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[944]),
        .S(self_sf7[944]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[945].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[945]),
        .S(self_sf7[945]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[946].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[946]),
        .S(self_sf7[946]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[947].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[947]),
        .S(self_sf7[947]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[948].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[948]),
        .S(self_sf7[948]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[949].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[949]),
        .S(self_sf7[949]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[94].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[94]),
        .S(self_sf7[94]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[950].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[950]),
        .S(self_sf7[950]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[951].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[951]),
        .S(self_sf7[951]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[952].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[952]),
        .S(self_sf7[952]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[953].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[953]),
        .S(self_sf7[953]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[954].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[954]),
        .S(self_sf7[954]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[955].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[955]),
        .S(self_sf7[955]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[956].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[956]),
        .S(self_sf7[956]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[957].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[957]),
        .S(self_sf7[957]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[958].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[958]),
        .S(self_sf7[958]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[959].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[959]),
        .S(self_sf7[959]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[95].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[95]),
        .S(self_sf7[95]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[960].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[960]),
        .S(self_sf7[960]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[961].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[961]),
        .S(self_sf7[961]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[962].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[962]),
        .S(self_sf7[962]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[963].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[963]),
        .S(self_sf7[963]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[964].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[964]),
        .S(self_sf7[964]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[965].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[965]),
        .S(self_sf7[965]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[966].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[966]),
        .S(self_sf7[966]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[967].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[967]),
        .S(self_sf7[967]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[968].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[968]),
        .S(self_sf7[968]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[969].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[969]),
        .S(self_sf7[969]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[96].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[96]),
        .S(self_sf7[96]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[970].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[970]),
        .S(self_sf7[970]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[971].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[971]),
        .S(self_sf7[971]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[972].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[972]),
        .S(self_sf7[972]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[973].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[973]),
        .S(self_sf7[973]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[974].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[974]),
        .S(self_sf7[974]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[975].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[975]),
        .S(self_sf7[975]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[976].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[976]),
        .S(self_sf7[976]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[977].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[977]),
        .S(self_sf7[977]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[978].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[978]),
        .S(self_sf7[978]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[979].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[979]),
        .S(self_sf7[979]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[97].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[97]),
        .S(self_sf7[97]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[980].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[980]),
        .S(self_sf7[980]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[981].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[981]),
        .S(self_sf7[981]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[982].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[982]),
        .S(self_sf7[982]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[983].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[983]),
        .S(self_sf7[983]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[984].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[984]),
        .S(self_sf7[984]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[985].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[985]),
        .S(self_sf7[985]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[986].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[986]),
        .S(self_sf7[986]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[987].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[987]),
        .S(self_sf7[987]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[988].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[988]),
        .S(self_sf7[988]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[989].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[989]),
        .S(self_sf7[989]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[98].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[98]),
        .S(self_sf7[98]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[990].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[990]),
        .S(self_sf7[990]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[991].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[991]),
        .S(self_sf7[991]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[992].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[992]),
        .S(self_sf7[992]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[993].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[993]),
        .S(self_sf7[993]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[994].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[994]),
        .S(self_sf7[994]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[995].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[995]),
        .S(self_sf7[995]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[996].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[996]),
        .S(self_sf7[996]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[997].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[997]),
        .S(self_sf7[997]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[998].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[998]),
        .S(self_sf7[998]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[999].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[999]),
        .S(self_sf7[999]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[99].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[99]),
        .S(self_sf7[99]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[9].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[9]),
        .S(self_sf7[9]));
  (* BOX_TYPE = "black_box" *) 
  MUXF8 \activity_ROsf8[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf8[0]),
        .S(self_sf8[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF9 \activity_ROsf9[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf9[0]),
        .S(self_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_0
       (.I0(1'b0),
        .O(self_sf7[1802]));
  LUT1 #(
    .INIT(2'h2)) 
    i_1
       (.I0(1'b0),
        .O(self_sf7[1801]));
  LUT1 #(
    .INIT(2'h2)) 
    i_10
       (.I0(1'b0),
        .O(info_sf8[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_11
       (.I0(1'b0),
        .O(info_sf8[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_12
       (.I0(1'b0),
        .O(info_sf8[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_13
       (.I0(1'b0),
        .O(info_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_14
       (.I0(1'b0),
        .O(info_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_15
       (.I0(1'b0),
        .O(info_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_16
       (.I0(1'b0),
        .O(info_sf8[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_17
       (.I0(1'b0),
        .O(info_sf9[7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_18
       (.I0(1'b0),
        .O(info_sf9[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_19
       (.I0(1'b0),
        .O(info_sf9[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_2
       (.I0(1'b0),
        .O(self_sf7[1800]));
  LUT1 #(
    .INIT(2'h2)) 
    i_20
       (.I0(1'b0),
        .O(info_sf9[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_21
       (.I0(1'b0),
        .O(info_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_22
       (.I0(1'b0),
        .O(info_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_23
       (.I0(1'b0),
        .O(info_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_24
       (.I0(1'b0),
        .O(info_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_3
       (.I0(1'b0),
        .O(self_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_4
       (.I0(1'b0),
        .O(self_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_5
       (.I0(1'b0),
        .O(self_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_6
       (.I0(1'b0),
        .O(self_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_7
       (.I0(1'b0),
        .O(self_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_8
       (.I0(1'b0),
        .O(self_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_9
       (.I0(1'b0),
        .O(info_sf8[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst
       (.I0(self_sf7[7]),
        .O(info_sf7[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__0
       (.I0(self_sf7[6]),
        .O(info_sf7[6]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__1
       (.I0(self_sf7[5]),
        .O(info_sf7[5]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__2
       (.I0(self_sf7[4]),
        .O(info_sf7[4]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__3
       (.I0(self_sf7[3]),
        .O(info_sf7[3]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__4
       (.I0(self_sf7[2]),
        .O(info_sf7[2]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__5
       (.I0(self_sf7[1]),
        .O(info_sf7[1]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__6
       (.I0(self_sf7[0]),
        .O(info_sf7[0]));
endmodule

(* ORIG_REF_NAME = "muxer" *) (* box_type = "black_box" *) (* dont_touch = "true" *) 
module switch_elements_muxer__1
   (enable_i,
    info_o);
  input enable_i;
  output info_o;

  wire enable_i;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf7;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf8;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf9;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [1802:0]self_sf7;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf8;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf9;

  assign info_o = info_sf7[1];
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[0]),
        .S(info_sf7[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1000].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1000]),
        .S(self_sf7[1000]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1001].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1001]),
        .S(self_sf7[1001]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1002].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1002]),
        .S(self_sf7[1002]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1003].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1003]),
        .S(self_sf7[1003]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1004].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1004]),
        .S(self_sf7[1004]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1005].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1005]),
        .S(self_sf7[1005]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1006].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1006]),
        .S(self_sf7[1006]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1007].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1007]),
        .S(self_sf7[1007]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1008].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1008]),
        .S(self_sf7[1008]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1009].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1009]),
        .S(self_sf7[1009]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[100]),
        .S(self_sf7[100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1010].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1010]),
        .S(self_sf7[1010]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1011].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1011]),
        .S(self_sf7[1011]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1012].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1012]),
        .S(self_sf7[1012]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1013].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1013]),
        .S(self_sf7[1013]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1014].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1014]),
        .S(self_sf7[1014]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1015].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1015]),
        .S(self_sf7[1015]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1016].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1016]),
        .S(self_sf7[1016]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1017].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1017]),
        .S(self_sf7[1017]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1018].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1018]),
        .S(self_sf7[1018]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1019].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1019]),
        .S(self_sf7[1019]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[101]),
        .S(self_sf7[101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1020].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1020]),
        .S(self_sf7[1020]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1021].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1021]),
        .S(self_sf7[1021]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1022].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1022]),
        .S(self_sf7[1022]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1023].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1023]),
        .S(self_sf7[1023]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1024].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1024]),
        .S(self_sf7[1024]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1025].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1025]),
        .S(self_sf7[1025]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1026].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1026]),
        .S(self_sf7[1026]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1027].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1027]),
        .S(self_sf7[1027]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1028].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1028]),
        .S(self_sf7[1028]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1029].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1029]),
        .S(self_sf7[1029]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[102]),
        .S(self_sf7[102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1030].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1030]),
        .S(self_sf7[1030]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1031].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1031]),
        .S(self_sf7[1031]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1032].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1032]),
        .S(self_sf7[1032]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1033].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1033]),
        .S(self_sf7[1033]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1034].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1034]),
        .S(self_sf7[1034]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1035].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1035]),
        .S(self_sf7[1035]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1036].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1036]),
        .S(self_sf7[1036]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1037].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1037]),
        .S(self_sf7[1037]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1038].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1038]),
        .S(self_sf7[1038]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1039].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1039]),
        .S(self_sf7[1039]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[103]),
        .S(self_sf7[103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1040].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1040]),
        .S(self_sf7[1040]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1041].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1041]),
        .S(self_sf7[1041]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1042].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1042]),
        .S(self_sf7[1042]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1043].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1043]),
        .S(self_sf7[1043]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1044].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1044]),
        .S(self_sf7[1044]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1045].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1045]),
        .S(self_sf7[1045]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1046].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1046]),
        .S(self_sf7[1046]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1047].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1047]),
        .S(self_sf7[1047]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1048].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1048]),
        .S(self_sf7[1048]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1049].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1049]),
        .S(self_sf7[1049]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[104]),
        .S(self_sf7[104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1050].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1050]),
        .S(self_sf7[1050]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1051].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1051]),
        .S(self_sf7[1051]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1052].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1052]),
        .S(self_sf7[1052]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1053].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1053]),
        .S(self_sf7[1053]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1054].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1054]),
        .S(self_sf7[1054]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1055].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1055]),
        .S(self_sf7[1055]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1056].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1056]),
        .S(self_sf7[1056]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1057].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1057]),
        .S(self_sf7[1057]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1058].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1058]),
        .S(self_sf7[1058]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1059].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1059]),
        .S(self_sf7[1059]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[105]),
        .S(self_sf7[105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1060].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1060]),
        .S(self_sf7[1060]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1061].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1061]),
        .S(self_sf7[1061]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1062].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1062]),
        .S(self_sf7[1062]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1063].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1063]),
        .S(self_sf7[1063]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1064].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1064]),
        .S(self_sf7[1064]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1065].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1065]),
        .S(self_sf7[1065]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1066].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1066]),
        .S(self_sf7[1066]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1067].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1067]),
        .S(self_sf7[1067]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1068].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1068]),
        .S(self_sf7[1068]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1069].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1069]),
        .S(self_sf7[1069]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[106]),
        .S(self_sf7[106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1070].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1070]),
        .S(self_sf7[1070]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1071].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1071]),
        .S(self_sf7[1071]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1072].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1072]),
        .S(self_sf7[1072]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1073].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1073]),
        .S(self_sf7[1073]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1074].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1074]),
        .S(self_sf7[1074]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1075].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1075]),
        .S(self_sf7[1075]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1076].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1076]),
        .S(self_sf7[1076]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1077].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1077]),
        .S(self_sf7[1077]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1078].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1078]),
        .S(self_sf7[1078]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1079].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1079]),
        .S(self_sf7[1079]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[107]),
        .S(self_sf7[107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1080].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1080]),
        .S(self_sf7[1080]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1081].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1081]),
        .S(self_sf7[1081]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1082].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1082]),
        .S(self_sf7[1082]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1083].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1083]),
        .S(self_sf7[1083]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1084].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1084]),
        .S(self_sf7[1084]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1085].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1085]),
        .S(self_sf7[1085]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1086].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1086]),
        .S(self_sf7[1086]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1087].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1087]),
        .S(self_sf7[1087]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1088].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1088]),
        .S(self_sf7[1088]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1089].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1089]),
        .S(self_sf7[1089]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[108]),
        .S(self_sf7[108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1090].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1090]),
        .S(self_sf7[1090]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1091].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1091]),
        .S(self_sf7[1091]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1092].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1092]),
        .S(self_sf7[1092]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1093].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1093]),
        .S(self_sf7[1093]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1094].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1094]),
        .S(self_sf7[1094]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1095].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1095]),
        .S(self_sf7[1095]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1096].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1096]),
        .S(self_sf7[1096]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1097].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1097]),
        .S(self_sf7[1097]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1098].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1098]),
        .S(self_sf7[1098]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1099].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1099]),
        .S(self_sf7[1099]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[109]),
        .S(self_sf7[109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[10].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[10]),
        .S(self_sf7[10]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1100]),
        .S(self_sf7[1100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1101]),
        .S(self_sf7[1101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1102]),
        .S(self_sf7[1102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1103]),
        .S(self_sf7[1103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1104]),
        .S(self_sf7[1104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1105]),
        .S(self_sf7[1105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1106]),
        .S(self_sf7[1106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1107]),
        .S(self_sf7[1107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1108]),
        .S(self_sf7[1108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1109]),
        .S(self_sf7[1109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[110]),
        .S(self_sf7[110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1110]),
        .S(self_sf7[1110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1111]),
        .S(self_sf7[1111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1112]),
        .S(self_sf7[1112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1113]),
        .S(self_sf7[1113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1114]),
        .S(self_sf7[1114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1115]),
        .S(self_sf7[1115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1116]),
        .S(self_sf7[1116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1117]),
        .S(self_sf7[1117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1118]),
        .S(self_sf7[1118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1119]),
        .S(self_sf7[1119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[111]),
        .S(self_sf7[111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1120]),
        .S(self_sf7[1120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1121]),
        .S(self_sf7[1121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1122]),
        .S(self_sf7[1122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1123]),
        .S(self_sf7[1123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1124]),
        .S(self_sf7[1124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1125]),
        .S(self_sf7[1125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1126]),
        .S(self_sf7[1126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1127]),
        .S(self_sf7[1127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1128]),
        .S(self_sf7[1128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1129]),
        .S(self_sf7[1129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[112]),
        .S(self_sf7[112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1130]),
        .S(self_sf7[1130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1131]),
        .S(self_sf7[1131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1132]),
        .S(self_sf7[1132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1133]),
        .S(self_sf7[1133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1134]),
        .S(self_sf7[1134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1135]),
        .S(self_sf7[1135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1136]),
        .S(self_sf7[1136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1137]),
        .S(self_sf7[1137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1138]),
        .S(self_sf7[1138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1139]),
        .S(self_sf7[1139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[113]),
        .S(self_sf7[113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1140]),
        .S(self_sf7[1140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1141]),
        .S(self_sf7[1141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1142]),
        .S(self_sf7[1142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1143]),
        .S(self_sf7[1143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1144]),
        .S(self_sf7[1144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1145]),
        .S(self_sf7[1145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1146]),
        .S(self_sf7[1146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1147]),
        .S(self_sf7[1147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1148]),
        .S(self_sf7[1148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1149]),
        .S(self_sf7[1149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[114]),
        .S(self_sf7[114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1150]),
        .S(self_sf7[1150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1151]),
        .S(self_sf7[1151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1152]),
        .S(self_sf7[1152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1153]),
        .S(self_sf7[1153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1154]),
        .S(self_sf7[1154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1155]),
        .S(self_sf7[1155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1156]),
        .S(self_sf7[1156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1157]),
        .S(self_sf7[1157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1158]),
        .S(self_sf7[1158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1159]),
        .S(self_sf7[1159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[115]),
        .S(self_sf7[115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1160]),
        .S(self_sf7[1160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1161]),
        .S(self_sf7[1161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1162]),
        .S(self_sf7[1162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1163]),
        .S(self_sf7[1163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1164]),
        .S(self_sf7[1164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1165]),
        .S(self_sf7[1165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1166]),
        .S(self_sf7[1166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1167]),
        .S(self_sf7[1167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1168]),
        .S(self_sf7[1168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1169]),
        .S(self_sf7[1169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[116]),
        .S(self_sf7[116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1170]),
        .S(self_sf7[1170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1171]),
        .S(self_sf7[1171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1172]),
        .S(self_sf7[1172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1173]),
        .S(self_sf7[1173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1174]),
        .S(self_sf7[1174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1175]),
        .S(self_sf7[1175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1176]),
        .S(self_sf7[1176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1177]),
        .S(self_sf7[1177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1178]),
        .S(self_sf7[1178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1179]),
        .S(self_sf7[1179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[117]),
        .S(self_sf7[117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1180]),
        .S(self_sf7[1180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1181]),
        .S(self_sf7[1181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1182]),
        .S(self_sf7[1182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1183]),
        .S(self_sf7[1183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1184]),
        .S(self_sf7[1184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1185]),
        .S(self_sf7[1185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1186]),
        .S(self_sf7[1186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1187]),
        .S(self_sf7[1187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1188]),
        .S(self_sf7[1188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1189]),
        .S(self_sf7[1189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[118]),
        .S(self_sf7[118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1190]),
        .S(self_sf7[1190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1191]),
        .S(self_sf7[1191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1192]),
        .S(self_sf7[1192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1193]),
        .S(self_sf7[1193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1194]),
        .S(self_sf7[1194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1195]),
        .S(self_sf7[1195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1196]),
        .S(self_sf7[1196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1197]),
        .S(self_sf7[1197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1198]),
        .S(self_sf7[1198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1199]),
        .S(self_sf7[1199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[119]),
        .S(self_sf7[119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[11].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[11]),
        .S(self_sf7[11]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1200]),
        .S(self_sf7[1200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1201]),
        .S(self_sf7[1201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1202]),
        .S(self_sf7[1202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1203]),
        .S(self_sf7[1203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1204]),
        .S(self_sf7[1204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1205]),
        .S(self_sf7[1205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1206]),
        .S(self_sf7[1206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1207]),
        .S(self_sf7[1207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1208]),
        .S(self_sf7[1208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1209]),
        .S(self_sf7[1209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[120]),
        .S(self_sf7[120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1210]),
        .S(self_sf7[1210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1211]),
        .S(self_sf7[1211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1212]),
        .S(self_sf7[1212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1213]),
        .S(self_sf7[1213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1214]),
        .S(self_sf7[1214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1215]),
        .S(self_sf7[1215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1216]),
        .S(self_sf7[1216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1217]),
        .S(self_sf7[1217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1218]),
        .S(self_sf7[1218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1219]),
        .S(self_sf7[1219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[121]),
        .S(self_sf7[121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1220]),
        .S(self_sf7[1220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1221]),
        .S(self_sf7[1221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1222]),
        .S(self_sf7[1222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1223]),
        .S(self_sf7[1223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1224]),
        .S(self_sf7[1224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1225]),
        .S(self_sf7[1225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1226]),
        .S(self_sf7[1226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1227]),
        .S(self_sf7[1227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1228]),
        .S(self_sf7[1228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1229]),
        .S(self_sf7[1229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[122]),
        .S(self_sf7[122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1230]),
        .S(self_sf7[1230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1231]),
        .S(self_sf7[1231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1232]),
        .S(self_sf7[1232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1233]),
        .S(self_sf7[1233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1234]),
        .S(self_sf7[1234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1235]),
        .S(self_sf7[1235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1236]),
        .S(self_sf7[1236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1237]),
        .S(self_sf7[1237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1238]),
        .S(self_sf7[1238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1239]),
        .S(self_sf7[1239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[123]),
        .S(self_sf7[123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1240]),
        .S(self_sf7[1240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1241]),
        .S(self_sf7[1241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1242]),
        .S(self_sf7[1242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1243]),
        .S(self_sf7[1243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1244]),
        .S(self_sf7[1244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1245]),
        .S(self_sf7[1245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1246]),
        .S(self_sf7[1246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1247]),
        .S(self_sf7[1247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1248]),
        .S(self_sf7[1248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1249]),
        .S(self_sf7[1249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[124]),
        .S(self_sf7[124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1250]),
        .S(self_sf7[1250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1251]),
        .S(self_sf7[1251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1252]),
        .S(self_sf7[1252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1253]),
        .S(self_sf7[1253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1254]),
        .S(self_sf7[1254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1255]),
        .S(self_sf7[1255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1256]),
        .S(self_sf7[1256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1257]),
        .S(self_sf7[1257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1258]),
        .S(self_sf7[1258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1259]),
        .S(self_sf7[1259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[125]),
        .S(self_sf7[125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1260]),
        .S(self_sf7[1260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1261]),
        .S(self_sf7[1261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1262]),
        .S(self_sf7[1262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1263]),
        .S(self_sf7[1263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1264]),
        .S(self_sf7[1264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1265]),
        .S(self_sf7[1265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1266]),
        .S(self_sf7[1266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1267]),
        .S(self_sf7[1267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1268]),
        .S(self_sf7[1268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1269]),
        .S(self_sf7[1269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[126]),
        .S(self_sf7[126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1270]),
        .S(self_sf7[1270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1271]),
        .S(self_sf7[1271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1272]),
        .S(self_sf7[1272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1273]),
        .S(self_sf7[1273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1274]),
        .S(self_sf7[1274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1275]),
        .S(self_sf7[1275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1276]),
        .S(self_sf7[1276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1277]),
        .S(self_sf7[1277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1278]),
        .S(self_sf7[1278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1279]),
        .S(self_sf7[1279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[127]),
        .S(self_sf7[127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1280]),
        .S(self_sf7[1280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1281]),
        .S(self_sf7[1281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1282]),
        .S(self_sf7[1282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1283]),
        .S(self_sf7[1283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1284]),
        .S(self_sf7[1284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1285]),
        .S(self_sf7[1285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1286]),
        .S(self_sf7[1286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1287]),
        .S(self_sf7[1287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1288]),
        .S(self_sf7[1288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1289]),
        .S(self_sf7[1289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[128]),
        .S(self_sf7[128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1290]),
        .S(self_sf7[1290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1291]),
        .S(self_sf7[1291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1292]),
        .S(self_sf7[1292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1293]),
        .S(self_sf7[1293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1294]),
        .S(self_sf7[1294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1295]),
        .S(self_sf7[1295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1296]),
        .S(self_sf7[1296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1297]),
        .S(self_sf7[1297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1298]),
        .S(self_sf7[1298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1299]),
        .S(self_sf7[1299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[129]),
        .S(self_sf7[129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[12].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[12]),
        .S(self_sf7[12]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1300]),
        .S(self_sf7[1300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1301]),
        .S(self_sf7[1301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1302]),
        .S(self_sf7[1302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1303]),
        .S(self_sf7[1303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1304]),
        .S(self_sf7[1304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1305]),
        .S(self_sf7[1305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1306]),
        .S(self_sf7[1306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1307]),
        .S(self_sf7[1307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1308]),
        .S(self_sf7[1308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1309]),
        .S(self_sf7[1309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[130]),
        .S(self_sf7[130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1310]),
        .S(self_sf7[1310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1311]),
        .S(self_sf7[1311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1312]),
        .S(self_sf7[1312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1313]),
        .S(self_sf7[1313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1314]),
        .S(self_sf7[1314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1315]),
        .S(self_sf7[1315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1316]),
        .S(self_sf7[1316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1317]),
        .S(self_sf7[1317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1318]),
        .S(self_sf7[1318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1319]),
        .S(self_sf7[1319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[131]),
        .S(self_sf7[131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1320]),
        .S(self_sf7[1320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1321]),
        .S(self_sf7[1321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1322]),
        .S(self_sf7[1322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1323]),
        .S(self_sf7[1323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1324]),
        .S(self_sf7[1324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1325]),
        .S(self_sf7[1325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1326]),
        .S(self_sf7[1326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1327]),
        .S(self_sf7[1327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1328]),
        .S(self_sf7[1328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1329]),
        .S(self_sf7[1329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[132]),
        .S(self_sf7[132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1330]),
        .S(self_sf7[1330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1331]),
        .S(self_sf7[1331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1332]),
        .S(self_sf7[1332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1333]),
        .S(self_sf7[1333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1334]),
        .S(self_sf7[1334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1335]),
        .S(self_sf7[1335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1336]),
        .S(self_sf7[1336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1337]),
        .S(self_sf7[1337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1338]),
        .S(self_sf7[1338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1339]),
        .S(self_sf7[1339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[133]),
        .S(self_sf7[133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1340]),
        .S(self_sf7[1340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1341]),
        .S(self_sf7[1341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1342]),
        .S(self_sf7[1342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1343]),
        .S(self_sf7[1343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1344]),
        .S(self_sf7[1344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1345]),
        .S(self_sf7[1345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1346]),
        .S(self_sf7[1346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1347]),
        .S(self_sf7[1347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1348]),
        .S(self_sf7[1348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1349]),
        .S(self_sf7[1349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[134]),
        .S(self_sf7[134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1350]),
        .S(self_sf7[1350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1351]),
        .S(self_sf7[1351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1352]),
        .S(self_sf7[1352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1353]),
        .S(self_sf7[1353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1354]),
        .S(self_sf7[1354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1355]),
        .S(self_sf7[1355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1356]),
        .S(self_sf7[1356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1357]),
        .S(self_sf7[1357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1358]),
        .S(self_sf7[1358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1359]),
        .S(self_sf7[1359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[135]),
        .S(self_sf7[135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1360]),
        .S(self_sf7[1360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1361]),
        .S(self_sf7[1361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1362]),
        .S(self_sf7[1362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1363]),
        .S(self_sf7[1363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1364]),
        .S(self_sf7[1364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1365]),
        .S(self_sf7[1365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1366]),
        .S(self_sf7[1366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1367]),
        .S(self_sf7[1367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1368]),
        .S(self_sf7[1368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1369]),
        .S(self_sf7[1369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[136]),
        .S(self_sf7[136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1370]),
        .S(self_sf7[1370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1371]),
        .S(self_sf7[1371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1372]),
        .S(self_sf7[1372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1373]),
        .S(self_sf7[1373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1374]),
        .S(self_sf7[1374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1375]),
        .S(self_sf7[1375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1376]),
        .S(self_sf7[1376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1377]),
        .S(self_sf7[1377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1378]),
        .S(self_sf7[1378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1379]),
        .S(self_sf7[1379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[137]),
        .S(self_sf7[137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1380]),
        .S(self_sf7[1380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1381]),
        .S(self_sf7[1381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1382]),
        .S(self_sf7[1382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1383]),
        .S(self_sf7[1383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1384]),
        .S(self_sf7[1384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1385]),
        .S(self_sf7[1385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1386]),
        .S(self_sf7[1386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1387]),
        .S(self_sf7[1387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1388]),
        .S(self_sf7[1388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1389]),
        .S(self_sf7[1389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[138]),
        .S(self_sf7[138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1390]),
        .S(self_sf7[1390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1391]),
        .S(self_sf7[1391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1392]),
        .S(self_sf7[1392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1393]),
        .S(self_sf7[1393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1394]),
        .S(self_sf7[1394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1395]),
        .S(self_sf7[1395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1396]),
        .S(self_sf7[1396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1397]),
        .S(self_sf7[1397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1398]),
        .S(self_sf7[1398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1399]),
        .S(self_sf7[1399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[139]),
        .S(self_sf7[139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[13].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[13]),
        .S(self_sf7[13]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1400]),
        .S(self_sf7[1400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1401]),
        .S(self_sf7[1401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1402]),
        .S(self_sf7[1402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1403]),
        .S(self_sf7[1403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1404]),
        .S(self_sf7[1404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1405]),
        .S(self_sf7[1405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1406]),
        .S(self_sf7[1406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1407]),
        .S(self_sf7[1407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1408]),
        .S(self_sf7[1408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1409]),
        .S(self_sf7[1409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[140]),
        .S(self_sf7[140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1410]),
        .S(self_sf7[1410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1411]),
        .S(self_sf7[1411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1412]),
        .S(self_sf7[1412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1413]),
        .S(self_sf7[1413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1414]),
        .S(self_sf7[1414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1415]),
        .S(self_sf7[1415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1416]),
        .S(self_sf7[1416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1417]),
        .S(self_sf7[1417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1418]),
        .S(self_sf7[1418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1419]),
        .S(self_sf7[1419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[141]),
        .S(self_sf7[141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1420]),
        .S(self_sf7[1420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1421]),
        .S(self_sf7[1421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1422]),
        .S(self_sf7[1422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1423]),
        .S(self_sf7[1423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1424]),
        .S(self_sf7[1424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1425]),
        .S(self_sf7[1425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1426]),
        .S(self_sf7[1426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1427]),
        .S(self_sf7[1427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1428]),
        .S(self_sf7[1428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1429]),
        .S(self_sf7[1429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[142]),
        .S(self_sf7[142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1430]),
        .S(self_sf7[1430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1431]),
        .S(self_sf7[1431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1432]),
        .S(self_sf7[1432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1433]),
        .S(self_sf7[1433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1434]),
        .S(self_sf7[1434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1435]),
        .S(self_sf7[1435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1436]),
        .S(self_sf7[1436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1437]),
        .S(self_sf7[1437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1438]),
        .S(self_sf7[1438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1439]),
        .S(self_sf7[1439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[143]),
        .S(self_sf7[143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1440]),
        .S(self_sf7[1440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1441]),
        .S(self_sf7[1441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1442]),
        .S(self_sf7[1442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1443]),
        .S(self_sf7[1443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1444]),
        .S(self_sf7[1444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1445]),
        .S(self_sf7[1445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1446]),
        .S(self_sf7[1446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1447]),
        .S(self_sf7[1447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1448]),
        .S(self_sf7[1448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1449]),
        .S(self_sf7[1449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[144]),
        .S(self_sf7[144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1450]),
        .S(self_sf7[1450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1451]),
        .S(self_sf7[1451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1452]),
        .S(self_sf7[1452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1453]),
        .S(self_sf7[1453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1454]),
        .S(self_sf7[1454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1455]),
        .S(self_sf7[1455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1456]),
        .S(self_sf7[1456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1457]),
        .S(self_sf7[1457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1458]),
        .S(self_sf7[1458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1459]),
        .S(self_sf7[1459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[145]),
        .S(self_sf7[145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1460]),
        .S(self_sf7[1460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1461]),
        .S(self_sf7[1461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1462]),
        .S(self_sf7[1462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1463]),
        .S(self_sf7[1463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1464]),
        .S(self_sf7[1464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1465]),
        .S(self_sf7[1465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1466]),
        .S(self_sf7[1466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1467]),
        .S(self_sf7[1467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1468]),
        .S(self_sf7[1468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1469]),
        .S(self_sf7[1469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[146]),
        .S(self_sf7[146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1470]),
        .S(self_sf7[1470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1471]),
        .S(self_sf7[1471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1472]),
        .S(self_sf7[1472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1473]),
        .S(self_sf7[1473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1474]),
        .S(self_sf7[1474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1475]),
        .S(self_sf7[1475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1476]),
        .S(self_sf7[1476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1477]),
        .S(self_sf7[1477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1478]),
        .S(self_sf7[1478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1479]),
        .S(self_sf7[1479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[147]),
        .S(self_sf7[147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1480]),
        .S(self_sf7[1480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1481]),
        .S(self_sf7[1481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1482]),
        .S(self_sf7[1482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1483]),
        .S(self_sf7[1483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1484]),
        .S(self_sf7[1484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1485]),
        .S(self_sf7[1485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1486]),
        .S(self_sf7[1486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1487]),
        .S(self_sf7[1487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1488]),
        .S(self_sf7[1488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1489]),
        .S(self_sf7[1489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[148]),
        .S(self_sf7[148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1490]),
        .S(self_sf7[1490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1491]),
        .S(self_sf7[1491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1492]),
        .S(self_sf7[1492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1493]),
        .S(self_sf7[1493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1494]),
        .S(self_sf7[1494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1495]),
        .S(self_sf7[1495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1496]),
        .S(self_sf7[1496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1497]),
        .S(self_sf7[1497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1498]),
        .S(self_sf7[1498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1499]),
        .S(self_sf7[1499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[149]),
        .S(self_sf7[149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[14].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[14]),
        .S(self_sf7[14]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1500]),
        .S(self_sf7[1500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1501]),
        .S(self_sf7[1501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1502]),
        .S(self_sf7[1502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1503]),
        .S(self_sf7[1503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1504]),
        .S(self_sf7[1504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1505]),
        .S(self_sf7[1505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1506]),
        .S(self_sf7[1506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1507]),
        .S(self_sf7[1507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1508]),
        .S(self_sf7[1508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1509]),
        .S(self_sf7[1509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[150]),
        .S(self_sf7[150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1510]),
        .S(self_sf7[1510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1511]),
        .S(self_sf7[1511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1512]),
        .S(self_sf7[1512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1513]),
        .S(self_sf7[1513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1514]),
        .S(self_sf7[1514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1515]),
        .S(self_sf7[1515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1516]),
        .S(self_sf7[1516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1517]),
        .S(self_sf7[1517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1518]),
        .S(self_sf7[1518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1519]),
        .S(self_sf7[1519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[151]),
        .S(self_sf7[151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1520]),
        .S(self_sf7[1520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1521]),
        .S(self_sf7[1521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1522]),
        .S(self_sf7[1522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1523]),
        .S(self_sf7[1523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1524]),
        .S(self_sf7[1524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1525]),
        .S(self_sf7[1525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1526]),
        .S(self_sf7[1526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1527]),
        .S(self_sf7[1527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1528]),
        .S(self_sf7[1528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1529]),
        .S(self_sf7[1529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[152]),
        .S(self_sf7[152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1530]),
        .S(self_sf7[1530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1531]),
        .S(self_sf7[1531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1532]),
        .S(self_sf7[1532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1533]),
        .S(self_sf7[1533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1534]),
        .S(self_sf7[1534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1535]),
        .S(self_sf7[1535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1536]),
        .S(self_sf7[1536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1537]),
        .S(self_sf7[1537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1538]),
        .S(self_sf7[1538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1539]),
        .S(self_sf7[1539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[153]),
        .S(self_sf7[153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1540]),
        .S(self_sf7[1540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1541]),
        .S(self_sf7[1541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1542]),
        .S(self_sf7[1542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1543]),
        .S(self_sf7[1543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1544]),
        .S(self_sf7[1544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1545]),
        .S(self_sf7[1545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1546]),
        .S(self_sf7[1546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1547]),
        .S(self_sf7[1547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1548]),
        .S(self_sf7[1548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1549]),
        .S(self_sf7[1549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[154]),
        .S(self_sf7[154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1550]),
        .S(self_sf7[1550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1551]),
        .S(self_sf7[1551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1552]),
        .S(self_sf7[1552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1553]),
        .S(self_sf7[1553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1554]),
        .S(self_sf7[1554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1555]),
        .S(self_sf7[1555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1556]),
        .S(self_sf7[1556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1557]),
        .S(self_sf7[1557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1558]),
        .S(self_sf7[1558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1559]),
        .S(self_sf7[1559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[155]),
        .S(self_sf7[155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1560]),
        .S(self_sf7[1560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1561]),
        .S(self_sf7[1561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1562]),
        .S(self_sf7[1562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1563]),
        .S(self_sf7[1563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1564]),
        .S(self_sf7[1564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1565]),
        .S(self_sf7[1565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1566]),
        .S(self_sf7[1566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1567]),
        .S(self_sf7[1567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1568]),
        .S(self_sf7[1568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1569]),
        .S(self_sf7[1569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[156]),
        .S(self_sf7[156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1570]),
        .S(self_sf7[1570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1571]),
        .S(self_sf7[1571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1572]),
        .S(self_sf7[1572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1573]),
        .S(self_sf7[1573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1574]),
        .S(self_sf7[1574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1575]),
        .S(self_sf7[1575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1576]),
        .S(self_sf7[1576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1577]),
        .S(self_sf7[1577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1578]),
        .S(self_sf7[1578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1579]),
        .S(self_sf7[1579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[157]),
        .S(self_sf7[157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1580]),
        .S(self_sf7[1580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1581]),
        .S(self_sf7[1581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1582]),
        .S(self_sf7[1582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1583]),
        .S(self_sf7[1583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1584]),
        .S(self_sf7[1584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1585]),
        .S(self_sf7[1585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1586]),
        .S(self_sf7[1586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1587]),
        .S(self_sf7[1587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1588]),
        .S(self_sf7[1588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1589]),
        .S(self_sf7[1589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[158]),
        .S(self_sf7[158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1590]),
        .S(self_sf7[1590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1591]),
        .S(self_sf7[1591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1592]),
        .S(self_sf7[1592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1593]),
        .S(self_sf7[1593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1594]),
        .S(self_sf7[1594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1595]),
        .S(self_sf7[1595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1596]),
        .S(self_sf7[1596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1597]),
        .S(self_sf7[1597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1598]),
        .S(self_sf7[1598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1599]),
        .S(self_sf7[1599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[159]),
        .S(self_sf7[159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[15].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[15]),
        .S(self_sf7[15]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1600]),
        .S(self_sf7[1600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1601]),
        .S(self_sf7[1601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1602]),
        .S(self_sf7[1602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1603]),
        .S(self_sf7[1603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1604]),
        .S(self_sf7[1604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1605]),
        .S(self_sf7[1605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1606]),
        .S(self_sf7[1606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1607]),
        .S(self_sf7[1607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1608]),
        .S(self_sf7[1608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1609]),
        .S(self_sf7[1609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[160]),
        .S(self_sf7[160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1610]),
        .S(self_sf7[1610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1611]),
        .S(self_sf7[1611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1612]),
        .S(self_sf7[1612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1613]),
        .S(self_sf7[1613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1614]),
        .S(self_sf7[1614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1615]),
        .S(self_sf7[1615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1616]),
        .S(self_sf7[1616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1617]),
        .S(self_sf7[1617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1618]),
        .S(self_sf7[1618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1619]),
        .S(self_sf7[1619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[161]),
        .S(self_sf7[161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1620]),
        .S(self_sf7[1620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1621]),
        .S(self_sf7[1621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1622]),
        .S(self_sf7[1622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1623]),
        .S(self_sf7[1623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1624]),
        .S(self_sf7[1624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1625]),
        .S(self_sf7[1625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1626]),
        .S(self_sf7[1626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1627]),
        .S(self_sf7[1627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1628]),
        .S(self_sf7[1628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1629]),
        .S(self_sf7[1629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[162]),
        .S(self_sf7[162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1630]),
        .S(self_sf7[1630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1631]),
        .S(self_sf7[1631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1632]),
        .S(self_sf7[1632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1633]),
        .S(self_sf7[1633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1634]),
        .S(self_sf7[1634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1635]),
        .S(self_sf7[1635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1636]),
        .S(self_sf7[1636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1637]),
        .S(self_sf7[1637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1638]),
        .S(self_sf7[1638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1639]),
        .S(self_sf7[1639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[163]),
        .S(self_sf7[163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1640]),
        .S(self_sf7[1640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1641]),
        .S(self_sf7[1641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1642]),
        .S(self_sf7[1642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1643]),
        .S(self_sf7[1643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1644]),
        .S(self_sf7[1644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1645]),
        .S(self_sf7[1645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1646]),
        .S(self_sf7[1646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1647]),
        .S(self_sf7[1647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1648]),
        .S(self_sf7[1648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1649]),
        .S(self_sf7[1649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[164]),
        .S(self_sf7[164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1650]),
        .S(self_sf7[1650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1651]),
        .S(self_sf7[1651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1652]),
        .S(self_sf7[1652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1653]),
        .S(self_sf7[1653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1654]),
        .S(self_sf7[1654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1655]),
        .S(self_sf7[1655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1656]),
        .S(self_sf7[1656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1657]),
        .S(self_sf7[1657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1658]),
        .S(self_sf7[1658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1659]),
        .S(self_sf7[1659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[165]),
        .S(self_sf7[165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1660]),
        .S(self_sf7[1660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1661]),
        .S(self_sf7[1661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1662]),
        .S(self_sf7[1662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1663]),
        .S(self_sf7[1663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1664]),
        .S(self_sf7[1664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1665]),
        .S(self_sf7[1665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1666]),
        .S(self_sf7[1666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1667]),
        .S(self_sf7[1667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1668]),
        .S(self_sf7[1668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1669]),
        .S(self_sf7[1669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[166]),
        .S(self_sf7[166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1670]),
        .S(self_sf7[1670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1671]),
        .S(self_sf7[1671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1672]),
        .S(self_sf7[1672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1673]),
        .S(self_sf7[1673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1674]),
        .S(self_sf7[1674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1675]),
        .S(self_sf7[1675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1676]),
        .S(self_sf7[1676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1677]),
        .S(self_sf7[1677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1678]),
        .S(self_sf7[1678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1679]),
        .S(self_sf7[1679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[167]),
        .S(self_sf7[167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1680]),
        .S(self_sf7[1680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1681]),
        .S(self_sf7[1681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1682]),
        .S(self_sf7[1682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1683]),
        .S(self_sf7[1683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1684]),
        .S(self_sf7[1684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1685]),
        .S(self_sf7[1685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1686]),
        .S(self_sf7[1686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1687]),
        .S(self_sf7[1687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1688]),
        .S(self_sf7[1688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1689]),
        .S(self_sf7[1689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[168]),
        .S(self_sf7[168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1690]),
        .S(self_sf7[1690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1691]),
        .S(self_sf7[1691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1692]),
        .S(self_sf7[1692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1693]),
        .S(self_sf7[1693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1694]),
        .S(self_sf7[1694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1695]),
        .S(self_sf7[1695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1696]),
        .S(self_sf7[1696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1697]),
        .S(self_sf7[1697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1698]),
        .S(self_sf7[1698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1699]),
        .S(self_sf7[1699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[169]),
        .S(self_sf7[169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[16].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[16]),
        .S(self_sf7[16]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1700]),
        .S(self_sf7[1700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1701]),
        .S(self_sf7[1701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1702]),
        .S(self_sf7[1702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1703]),
        .S(self_sf7[1703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1704]),
        .S(self_sf7[1704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1705]),
        .S(self_sf7[1705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1706]),
        .S(self_sf7[1706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1707]),
        .S(self_sf7[1707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1708]),
        .S(self_sf7[1708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1709]),
        .S(self_sf7[1709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[170]),
        .S(self_sf7[170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1710]),
        .S(self_sf7[1710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1711]),
        .S(self_sf7[1711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1712]),
        .S(self_sf7[1712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1713]),
        .S(self_sf7[1713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1714]),
        .S(self_sf7[1714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1715]),
        .S(self_sf7[1715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1716]),
        .S(self_sf7[1716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1717]),
        .S(self_sf7[1717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1718]),
        .S(self_sf7[1718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1719]),
        .S(self_sf7[1719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[171]),
        .S(self_sf7[171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1720]),
        .S(self_sf7[1720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1721]),
        .S(self_sf7[1721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1722]),
        .S(self_sf7[1722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1723]),
        .S(self_sf7[1723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1724]),
        .S(self_sf7[1724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1725]),
        .S(self_sf7[1725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1726]),
        .S(self_sf7[1726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1727]),
        .S(self_sf7[1727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1728]),
        .S(self_sf7[1728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1729]),
        .S(self_sf7[1729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[172]),
        .S(self_sf7[172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1730]),
        .S(self_sf7[1730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1731]),
        .S(self_sf7[1731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1732]),
        .S(self_sf7[1732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1733]),
        .S(self_sf7[1733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1734]),
        .S(self_sf7[1734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1735]),
        .S(self_sf7[1735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1736]),
        .S(self_sf7[1736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1737]),
        .S(self_sf7[1737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1738]),
        .S(self_sf7[1738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1739]),
        .S(self_sf7[1739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[173]),
        .S(self_sf7[173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1740]),
        .S(self_sf7[1740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1741]),
        .S(self_sf7[1741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1742]),
        .S(self_sf7[1742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1743]),
        .S(self_sf7[1743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1744]),
        .S(self_sf7[1744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1745]),
        .S(self_sf7[1745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1746]),
        .S(self_sf7[1746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1747]),
        .S(self_sf7[1747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1748]),
        .S(self_sf7[1748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1749]),
        .S(self_sf7[1749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[174]),
        .S(self_sf7[174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1750]),
        .S(self_sf7[1750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1751]),
        .S(self_sf7[1751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1752]),
        .S(self_sf7[1752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1753]),
        .S(self_sf7[1753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1754]),
        .S(self_sf7[1754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1755]),
        .S(self_sf7[1755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1756]),
        .S(self_sf7[1756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1757]),
        .S(self_sf7[1757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1758]),
        .S(self_sf7[1758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1759]),
        .S(self_sf7[1759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[175]),
        .S(self_sf7[175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1760]),
        .S(self_sf7[1760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1761]),
        .S(self_sf7[1761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1762]),
        .S(self_sf7[1762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1763]),
        .S(self_sf7[1763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1764]),
        .S(self_sf7[1764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1765]),
        .S(self_sf7[1765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1766]),
        .S(self_sf7[1766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1767]),
        .S(self_sf7[1767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1768]),
        .S(self_sf7[1768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1769]),
        .S(self_sf7[1769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[176]),
        .S(self_sf7[176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1770]),
        .S(self_sf7[1770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1771]),
        .S(self_sf7[1771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1772]),
        .S(self_sf7[1772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1773]),
        .S(self_sf7[1773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1774]),
        .S(self_sf7[1774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1775]),
        .S(self_sf7[1775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1776]),
        .S(self_sf7[1776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1777]),
        .S(self_sf7[1777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1778]),
        .S(self_sf7[1778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1779]),
        .S(self_sf7[1779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[177]),
        .S(self_sf7[177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1780]),
        .S(self_sf7[1780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1781]),
        .S(self_sf7[1781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1782]),
        .S(self_sf7[1782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1783]),
        .S(self_sf7[1783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1784]),
        .S(self_sf7[1784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1785]),
        .S(self_sf7[1785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1786]),
        .S(self_sf7[1786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1787]),
        .S(self_sf7[1787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1788]),
        .S(self_sf7[1788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1789]),
        .S(self_sf7[1789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[178]),
        .S(self_sf7[178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1790]),
        .S(self_sf7[1790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1791]),
        .S(self_sf7[1791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1792]),
        .S(self_sf7[1792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1793]),
        .S(self_sf7[1793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1794]),
        .S(self_sf7[1794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1795]),
        .S(self_sf7[1795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1796]),
        .S(self_sf7[1796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1797]),
        .S(self_sf7[1797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1798]),
        .S(self_sf7[1798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1799]),
        .S(self_sf7[1799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[179]),
        .S(self_sf7[179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[17].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[17]),
        .S(self_sf7[17]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[180]),
        .S(self_sf7[180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[181]),
        .S(self_sf7[181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[182]),
        .S(self_sf7[182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[183]),
        .S(self_sf7[183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[184]),
        .S(self_sf7[184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[185]),
        .S(self_sf7[185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[186]),
        .S(self_sf7[186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[187]),
        .S(self_sf7[187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[188]),
        .S(self_sf7[188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[189]),
        .S(self_sf7[189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[18].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[18]),
        .S(self_sf7[18]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[190]),
        .S(self_sf7[190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[191]),
        .S(self_sf7[191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[192]),
        .S(self_sf7[192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[193]),
        .S(self_sf7[193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[194]),
        .S(self_sf7[194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[195]),
        .S(self_sf7[195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[196]),
        .S(self_sf7[196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[197]),
        .S(self_sf7[197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[198]),
        .S(self_sf7[198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[199]),
        .S(self_sf7[199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[19].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[19]),
        .S(self_sf7[19]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1]),
        .S(info_sf7[1]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[200]),
        .S(self_sf7[200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[201]),
        .S(self_sf7[201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[202]),
        .S(self_sf7[202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[203]),
        .S(self_sf7[203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[204]),
        .S(self_sf7[204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[205]),
        .S(self_sf7[205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[206]),
        .S(self_sf7[206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[207]),
        .S(self_sf7[207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[208]),
        .S(self_sf7[208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[209]),
        .S(self_sf7[209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[20].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[20]),
        .S(self_sf7[20]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[210]),
        .S(self_sf7[210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[211]),
        .S(self_sf7[211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[212]),
        .S(self_sf7[212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[213]),
        .S(self_sf7[213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[214]),
        .S(self_sf7[214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[215]),
        .S(self_sf7[215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[216]),
        .S(self_sf7[216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[217]),
        .S(self_sf7[217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[218]),
        .S(self_sf7[218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[219]),
        .S(self_sf7[219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[21].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[21]),
        .S(self_sf7[21]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[220]),
        .S(self_sf7[220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[221]),
        .S(self_sf7[221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[222]),
        .S(self_sf7[222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[223]),
        .S(self_sf7[223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[224]),
        .S(self_sf7[224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[225]),
        .S(self_sf7[225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[226]),
        .S(self_sf7[226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[227]),
        .S(self_sf7[227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[228]),
        .S(self_sf7[228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[229]),
        .S(self_sf7[229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[22].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[22]),
        .S(self_sf7[22]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[230]),
        .S(self_sf7[230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[231]),
        .S(self_sf7[231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[232]),
        .S(self_sf7[232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[233]),
        .S(self_sf7[233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[234]),
        .S(self_sf7[234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[235]),
        .S(self_sf7[235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[236]),
        .S(self_sf7[236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[237]),
        .S(self_sf7[237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[238]),
        .S(self_sf7[238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[239]),
        .S(self_sf7[239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[23].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[23]),
        .S(self_sf7[23]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[240]),
        .S(self_sf7[240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[241]),
        .S(self_sf7[241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[242]),
        .S(self_sf7[242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[243]),
        .S(self_sf7[243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[244]),
        .S(self_sf7[244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[245]),
        .S(self_sf7[245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[246]),
        .S(self_sf7[246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[247]),
        .S(self_sf7[247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[248]),
        .S(self_sf7[248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[249]),
        .S(self_sf7[249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[24].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[24]),
        .S(self_sf7[24]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[250]),
        .S(self_sf7[250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[251]),
        .S(self_sf7[251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[252]),
        .S(self_sf7[252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[253]),
        .S(self_sf7[253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[254]),
        .S(self_sf7[254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[255]),
        .S(self_sf7[255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[256]),
        .S(self_sf7[256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[257]),
        .S(self_sf7[257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[258]),
        .S(self_sf7[258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[259]),
        .S(self_sf7[259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[25].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[25]),
        .S(self_sf7[25]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[260]),
        .S(self_sf7[260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[261]),
        .S(self_sf7[261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[262]),
        .S(self_sf7[262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[263]),
        .S(self_sf7[263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[264]),
        .S(self_sf7[264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[265]),
        .S(self_sf7[265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[266]),
        .S(self_sf7[266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[267]),
        .S(self_sf7[267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[268]),
        .S(self_sf7[268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[269]),
        .S(self_sf7[269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[26].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[26]),
        .S(self_sf7[26]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[270]),
        .S(self_sf7[270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[271]),
        .S(self_sf7[271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[272]),
        .S(self_sf7[272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[273]),
        .S(self_sf7[273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[274]),
        .S(self_sf7[274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[275]),
        .S(self_sf7[275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[276]),
        .S(self_sf7[276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[277]),
        .S(self_sf7[277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[278]),
        .S(self_sf7[278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[279]),
        .S(self_sf7[279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[27].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[27]),
        .S(self_sf7[27]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[280]),
        .S(self_sf7[280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[281]),
        .S(self_sf7[281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[282]),
        .S(self_sf7[282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[283]),
        .S(self_sf7[283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[284]),
        .S(self_sf7[284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[285]),
        .S(self_sf7[285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[286]),
        .S(self_sf7[286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[287]),
        .S(self_sf7[287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[288]),
        .S(self_sf7[288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[289]),
        .S(self_sf7[289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[28].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[28]),
        .S(self_sf7[28]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[290]),
        .S(self_sf7[290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[291]),
        .S(self_sf7[291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[292]),
        .S(self_sf7[292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[293]),
        .S(self_sf7[293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[294]),
        .S(self_sf7[294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[295]),
        .S(self_sf7[295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[296]),
        .S(self_sf7[296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[297]),
        .S(self_sf7[297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[298]),
        .S(self_sf7[298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[299]),
        .S(self_sf7[299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[29].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[29]),
        .S(self_sf7[29]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[2].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[2]),
        .S(info_sf7[2]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[300]),
        .S(self_sf7[300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[301]),
        .S(self_sf7[301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[302]),
        .S(self_sf7[302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[303]),
        .S(self_sf7[303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[304]),
        .S(self_sf7[304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[305]),
        .S(self_sf7[305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[306]),
        .S(self_sf7[306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[307]),
        .S(self_sf7[307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[308]),
        .S(self_sf7[308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[309]),
        .S(self_sf7[309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[30].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[30]),
        .S(self_sf7[30]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[310]),
        .S(self_sf7[310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[311]),
        .S(self_sf7[311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[312]),
        .S(self_sf7[312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[313]),
        .S(self_sf7[313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[314]),
        .S(self_sf7[314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[315]),
        .S(self_sf7[315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[316]),
        .S(self_sf7[316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[317]),
        .S(self_sf7[317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[318]),
        .S(self_sf7[318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[319]),
        .S(self_sf7[319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[31].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[31]),
        .S(self_sf7[31]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[320]),
        .S(self_sf7[320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[321]),
        .S(self_sf7[321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[322]),
        .S(self_sf7[322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[323]),
        .S(self_sf7[323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[324]),
        .S(self_sf7[324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[325]),
        .S(self_sf7[325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[326]),
        .S(self_sf7[326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[327]),
        .S(self_sf7[327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[328]),
        .S(self_sf7[328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[329]),
        .S(self_sf7[329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[32].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[32]),
        .S(self_sf7[32]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[330]),
        .S(self_sf7[330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[331]),
        .S(self_sf7[331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[332]),
        .S(self_sf7[332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[333]),
        .S(self_sf7[333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[334]),
        .S(self_sf7[334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[335]),
        .S(self_sf7[335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[336]),
        .S(self_sf7[336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[337]),
        .S(self_sf7[337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[338]),
        .S(self_sf7[338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[339]),
        .S(self_sf7[339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[33].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[33]),
        .S(self_sf7[33]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[340]),
        .S(self_sf7[340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[341]),
        .S(self_sf7[341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[342]),
        .S(self_sf7[342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[343]),
        .S(self_sf7[343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[344]),
        .S(self_sf7[344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[345]),
        .S(self_sf7[345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[346]),
        .S(self_sf7[346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[347]),
        .S(self_sf7[347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[348]),
        .S(self_sf7[348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[349]),
        .S(self_sf7[349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[34].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[34]),
        .S(self_sf7[34]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[350]),
        .S(self_sf7[350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[351]),
        .S(self_sf7[351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[352]),
        .S(self_sf7[352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[353]),
        .S(self_sf7[353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[354]),
        .S(self_sf7[354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[355]),
        .S(self_sf7[355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[356]),
        .S(self_sf7[356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[357]),
        .S(self_sf7[357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[358]),
        .S(self_sf7[358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[359]),
        .S(self_sf7[359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[35].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[35]),
        .S(self_sf7[35]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[360]),
        .S(self_sf7[360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[361]),
        .S(self_sf7[361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[362]),
        .S(self_sf7[362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[363]),
        .S(self_sf7[363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[364]),
        .S(self_sf7[364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[365]),
        .S(self_sf7[365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[366]),
        .S(self_sf7[366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[367]),
        .S(self_sf7[367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[368]),
        .S(self_sf7[368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[369]),
        .S(self_sf7[369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[36].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[36]),
        .S(self_sf7[36]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[370]),
        .S(self_sf7[370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[371]),
        .S(self_sf7[371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[372]),
        .S(self_sf7[372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[373]),
        .S(self_sf7[373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[374]),
        .S(self_sf7[374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[375]),
        .S(self_sf7[375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[376]),
        .S(self_sf7[376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[377]),
        .S(self_sf7[377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[378]),
        .S(self_sf7[378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[379]),
        .S(self_sf7[379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[37].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[37]),
        .S(self_sf7[37]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[380]),
        .S(self_sf7[380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[381]),
        .S(self_sf7[381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[382]),
        .S(self_sf7[382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[383]),
        .S(self_sf7[383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[384]),
        .S(self_sf7[384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[385]),
        .S(self_sf7[385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[386]),
        .S(self_sf7[386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[387]),
        .S(self_sf7[387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[388]),
        .S(self_sf7[388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[389]),
        .S(self_sf7[389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[38].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[38]),
        .S(self_sf7[38]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[390]),
        .S(self_sf7[390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[391]),
        .S(self_sf7[391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[392]),
        .S(self_sf7[392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[393]),
        .S(self_sf7[393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[394]),
        .S(self_sf7[394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[395]),
        .S(self_sf7[395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[396]),
        .S(self_sf7[396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[397]),
        .S(self_sf7[397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[398]),
        .S(self_sf7[398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[399]),
        .S(self_sf7[399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[39].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[39]),
        .S(self_sf7[39]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[3].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[3]),
        .S(info_sf7[3]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[400]),
        .S(self_sf7[400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[401]),
        .S(self_sf7[401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[402]),
        .S(self_sf7[402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[403]),
        .S(self_sf7[403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[404]),
        .S(self_sf7[404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[405]),
        .S(self_sf7[405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[406]),
        .S(self_sf7[406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[407]),
        .S(self_sf7[407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[408]),
        .S(self_sf7[408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[409]),
        .S(self_sf7[409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[40].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[40]),
        .S(self_sf7[40]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[410]),
        .S(self_sf7[410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[411]),
        .S(self_sf7[411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[412]),
        .S(self_sf7[412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[413]),
        .S(self_sf7[413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[414]),
        .S(self_sf7[414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[415]),
        .S(self_sf7[415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[416]),
        .S(self_sf7[416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[417]),
        .S(self_sf7[417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[418]),
        .S(self_sf7[418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[419]),
        .S(self_sf7[419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[41].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[41]),
        .S(self_sf7[41]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[420]),
        .S(self_sf7[420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[421]),
        .S(self_sf7[421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[422]),
        .S(self_sf7[422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[423]),
        .S(self_sf7[423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[424]),
        .S(self_sf7[424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[425]),
        .S(self_sf7[425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[426]),
        .S(self_sf7[426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[427]),
        .S(self_sf7[427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[428]),
        .S(self_sf7[428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[429]),
        .S(self_sf7[429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[42].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[42]),
        .S(self_sf7[42]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[430]),
        .S(self_sf7[430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[431]),
        .S(self_sf7[431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[432]),
        .S(self_sf7[432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[433]),
        .S(self_sf7[433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[434]),
        .S(self_sf7[434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[435]),
        .S(self_sf7[435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[436]),
        .S(self_sf7[436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[437]),
        .S(self_sf7[437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[438]),
        .S(self_sf7[438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[439]),
        .S(self_sf7[439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[43].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[43]),
        .S(self_sf7[43]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[440]),
        .S(self_sf7[440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[441]),
        .S(self_sf7[441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[442]),
        .S(self_sf7[442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[443]),
        .S(self_sf7[443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[444]),
        .S(self_sf7[444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[445]),
        .S(self_sf7[445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[446]),
        .S(self_sf7[446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[447]),
        .S(self_sf7[447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[448]),
        .S(self_sf7[448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[449]),
        .S(self_sf7[449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[44].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[44]),
        .S(self_sf7[44]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[450]),
        .S(self_sf7[450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[451]),
        .S(self_sf7[451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[452]),
        .S(self_sf7[452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[453]),
        .S(self_sf7[453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[454]),
        .S(self_sf7[454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[455]),
        .S(self_sf7[455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[456]),
        .S(self_sf7[456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[457]),
        .S(self_sf7[457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[458]),
        .S(self_sf7[458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[459]),
        .S(self_sf7[459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[45].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[45]),
        .S(self_sf7[45]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[460]),
        .S(self_sf7[460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[461]),
        .S(self_sf7[461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[462]),
        .S(self_sf7[462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[463]),
        .S(self_sf7[463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[464]),
        .S(self_sf7[464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[465]),
        .S(self_sf7[465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[466]),
        .S(self_sf7[466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[467]),
        .S(self_sf7[467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[468]),
        .S(self_sf7[468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[469]),
        .S(self_sf7[469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[46].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[46]),
        .S(self_sf7[46]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[470]),
        .S(self_sf7[470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[471]),
        .S(self_sf7[471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[472]),
        .S(self_sf7[472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[473]),
        .S(self_sf7[473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[474]),
        .S(self_sf7[474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[475]),
        .S(self_sf7[475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[476]),
        .S(self_sf7[476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[477]),
        .S(self_sf7[477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[478]),
        .S(self_sf7[478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[479]),
        .S(self_sf7[479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[47].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[47]),
        .S(self_sf7[47]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[480]),
        .S(self_sf7[480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[481]),
        .S(self_sf7[481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[482]),
        .S(self_sf7[482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[483]),
        .S(self_sf7[483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[484]),
        .S(self_sf7[484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[485]),
        .S(self_sf7[485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[486]),
        .S(self_sf7[486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[487]),
        .S(self_sf7[487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[488]),
        .S(self_sf7[488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[489]),
        .S(self_sf7[489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[48].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[48]),
        .S(self_sf7[48]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[490]),
        .S(self_sf7[490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[491]),
        .S(self_sf7[491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[492]),
        .S(self_sf7[492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[493]),
        .S(self_sf7[493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[494]),
        .S(self_sf7[494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[495]),
        .S(self_sf7[495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[496]),
        .S(self_sf7[496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[497]),
        .S(self_sf7[497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[498]),
        .S(self_sf7[498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[499]),
        .S(self_sf7[499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[49].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[49]),
        .S(self_sf7[49]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[4].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[4]),
        .S(info_sf7[4]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[500]),
        .S(self_sf7[500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[501]),
        .S(self_sf7[501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[502]),
        .S(self_sf7[502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[503]),
        .S(self_sf7[503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[504]),
        .S(self_sf7[504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[505]),
        .S(self_sf7[505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[506]),
        .S(self_sf7[506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[507]),
        .S(self_sf7[507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[508]),
        .S(self_sf7[508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[509]),
        .S(self_sf7[509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[50].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[50]),
        .S(self_sf7[50]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[510]),
        .S(self_sf7[510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[511]),
        .S(self_sf7[511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[512]),
        .S(self_sf7[512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[513]),
        .S(self_sf7[513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[514]),
        .S(self_sf7[514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[515]),
        .S(self_sf7[515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[516]),
        .S(self_sf7[516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[517]),
        .S(self_sf7[517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[518]),
        .S(self_sf7[518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[519]),
        .S(self_sf7[519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[51].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[51]),
        .S(self_sf7[51]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[520]),
        .S(self_sf7[520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[521]),
        .S(self_sf7[521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[522]),
        .S(self_sf7[522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[523]),
        .S(self_sf7[523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[524]),
        .S(self_sf7[524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[525]),
        .S(self_sf7[525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[526]),
        .S(self_sf7[526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[527]),
        .S(self_sf7[527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[528]),
        .S(self_sf7[528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[529]),
        .S(self_sf7[529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[52].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[52]),
        .S(self_sf7[52]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[530]),
        .S(self_sf7[530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[531]),
        .S(self_sf7[531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[532]),
        .S(self_sf7[532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[533]),
        .S(self_sf7[533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[534]),
        .S(self_sf7[534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[535]),
        .S(self_sf7[535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[536]),
        .S(self_sf7[536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[537]),
        .S(self_sf7[537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[538]),
        .S(self_sf7[538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[539]),
        .S(self_sf7[539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[53].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[53]),
        .S(self_sf7[53]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[540]),
        .S(self_sf7[540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[541]),
        .S(self_sf7[541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[542]),
        .S(self_sf7[542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[543]),
        .S(self_sf7[543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[544]),
        .S(self_sf7[544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[545]),
        .S(self_sf7[545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[546]),
        .S(self_sf7[546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[547]),
        .S(self_sf7[547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[548]),
        .S(self_sf7[548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[549]),
        .S(self_sf7[549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[54].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[54]),
        .S(self_sf7[54]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[550]),
        .S(self_sf7[550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[551]),
        .S(self_sf7[551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[552]),
        .S(self_sf7[552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[553]),
        .S(self_sf7[553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[554]),
        .S(self_sf7[554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[555]),
        .S(self_sf7[555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[556]),
        .S(self_sf7[556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[557]),
        .S(self_sf7[557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[558]),
        .S(self_sf7[558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[559]),
        .S(self_sf7[559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[55].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[55]),
        .S(self_sf7[55]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[560]),
        .S(self_sf7[560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[561]),
        .S(self_sf7[561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[562]),
        .S(self_sf7[562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[563]),
        .S(self_sf7[563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[564]),
        .S(self_sf7[564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[565]),
        .S(self_sf7[565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[566]),
        .S(self_sf7[566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[567]),
        .S(self_sf7[567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[568]),
        .S(self_sf7[568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[569]),
        .S(self_sf7[569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[56].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[56]),
        .S(self_sf7[56]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[570]),
        .S(self_sf7[570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[571]),
        .S(self_sf7[571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[572]),
        .S(self_sf7[572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[573]),
        .S(self_sf7[573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[574]),
        .S(self_sf7[574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[575]),
        .S(self_sf7[575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[576]),
        .S(self_sf7[576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[577]),
        .S(self_sf7[577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[578]),
        .S(self_sf7[578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[579]),
        .S(self_sf7[579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[57].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[57]),
        .S(self_sf7[57]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[580]),
        .S(self_sf7[580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[581]),
        .S(self_sf7[581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[582]),
        .S(self_sf7[582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[583]),
        .S(self_sf7[583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[584]),
        .S(self_sf7[584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[585]),
        .S(self_sf7[585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[586]),
        .S(self_sf7[586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[587]),
        .S(self_sf7[587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[588]),
        .S(self_sf7[588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[589]),
        .S(self_sf7[589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[58].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[58]),
        .S(self_sf7[58]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[590]),
        .S(self_sf7[590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[591]),
        .S(self_sf7[591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[592]),
        .S(self_sf7[592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[593]),
        .S(self_sf7[593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[594]),
        .S(self_sf7[594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[595]),
        .S(self_sf7[595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[596]),
        .S(self_sf7[596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[597]),
        .S(self_sf7[597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[598]),
        .S(self_sf7[598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[599]),
        .S(self_sf7[599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[59].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[59]),
        .S(self_sf7[59]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[5].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[5]),
        .S(info_sf7[5]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[600]),
        .S(self_sf7[600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[601]),
        .S(self_sf7[601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[602]),
        .S(self_sf7[602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[603]),
        .S(self_sf7[603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[604]),
        .S(self_sf7[604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[605]),
        .S(self_sf7[605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[606]),
        .S(self_sf7[606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[607]),
        .S(self_sf7[607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[608]),
        .S(self_sf7[608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[609]),
        .S(self_sf7[609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[60].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[60]),
        .S(self_sf7[60]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[610]),
        .S(self_sf7[610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[611]),
        .S(self_sf7[611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[612]),
        .S(self_sf7[612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[613]),
        .S(self_sf7[613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[614]),
        .S(self_sf7[614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[615]),
        .S(self_sf7[615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[616]),
        .S(self_sf7[616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[617]),
        .S(self_sf7[617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[618]),
        .S(self_sf7[618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[619]),
        .S(self_sf7[619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[61].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[61]),
        .S(self_sf7[61]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[620]),
        .S(self_sf7[620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[621]),
        .S(self_sf7[621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[622]),
        .S(self_sf7[622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[623]),
        .S(self_sf7[623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[624]),
        .S(self_sf7[624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[625]),
        .S(self_sf7[625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[626]),
        .S(self_sf7[626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[627]),
        .S(self_sf7[627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[628]),
        .S(self_sf7[628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[629]),
        .S(self_sf7[629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[62].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[62]),
        .S(self_sf7[62]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[630]),
        .S(self_sf7[630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[631]),
        .S(self_sf7[631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[632]),
        .S(self_sf7[632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[633]),
        .S(self_sf7[633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[634]),
        .S(self_sf7[634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[635]),
        .S(self_sf7[635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[636]),
        .S(self_sf7[636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[637]),
        .S(self_sf7[637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[638]),
        .S(self_sf7[638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[639]),
        .S(self_sf7[639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[63].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[63]),
        .S(self_sf7[63]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[640]),
        .S(self_sf7[640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[641]),
        .S(self_sf7[641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[642]),
        .S(self_sf7[642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[643]),
        .S(self_sf7[643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[644]),
        .S(self_sf7[644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[645]),
        .S(self_sf7[645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[646]),
        .S(self_sf7[646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[647]),
        .S(self_sf7[647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[648]),
        .S(self_sf7[648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[649]),
        .S(self_sf7[649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[64].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[64]),
        .S(self_sf7[64]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[650]),
        .S(self_sf7[650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[651]),
        .S(self_sf7[651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[652]),
        .S(self_sf7[652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[653]),
        .S(self_sf7[653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[654]),
        .S(self_sf7[654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[655]),
        .S(self_sf7[655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[656]),
        .S(self_sf7[656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[657]),
        .S(self_sf7[657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[658]),
        .S(self_sf7[658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[659]),
        .S(self_sf7[659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[65].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[65]),
        .S(self_sf7[65]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[660]),
        .S(self_sf7[660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[661]),
        .S(self_sf7[661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[662]),
        .S(self_sf7[662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[663]),
        .S(self_sf7[663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[664]),
        .S(self_sf7[664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[665]),
        .S(self_sf7[665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[666]),
        .S(self_sf7[666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[667]),
        .S(self_sf7[667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[668]),
        .S(self_sf7[668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[669]),
        .S(self_sf7[669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[66].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[66]),
        .S(self_sf7[66]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[670]),
        .S(self_sf7[670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[671]),
        .S(self_sf7[671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[672]),
        .S(self_sf7[672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[673]),
        .S(self_sf7[673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[674]),
        .S(self_sf7[674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[675]),
        .S(self_sf7[675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[676]),
        .S(self_sf7[676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[677]),
        .S(self_sf7[677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[678]),
        .S(self_sf7[678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[679]),
        .S(self_sf7[679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[67].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[67]),
        .S(self_sf7[67]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[680]),
        .S(self_sf7[680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[681]),
        .S(self_sf7[681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[682]),
        .S(self_sf7[682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[683]),
        .S(self_sf7[683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[684]),
        .S(self_sf7[684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[685]),
        .S(self_sf7[685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[686]),
        .S(self_sf7[686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[687]),
        .S(self_sf7[687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[688]),
        .S(self_sf7[688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[689]),
        .S(self_sf7[689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[68].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[68]),
        .S(self_sf7[68]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[690]),
        .S(self_sf7[690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[691]),
        .S(self_sf7[691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[692]),
        .S(self_sf7[692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[693]),
        .S(self_sf7[693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[694]),
        .S(self_sf7[694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[695]),
        .S(self_sf7[695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[696]),
        .S(self_sf7[696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[697]),
        .S(self_sf7[697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[698]),
        .S(self_sf7[698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[699]),
        .S(self_sf7[699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[69].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[69]),
        .S(self_sf7[69]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[6].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[6]),
        .S(info_sf7[6]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[700]),
        .S(self_sf7[700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[701]),
        .S(self_sf7[701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[702]),
        .S(self_sf7[702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[703]),
        .S(self_sf7[703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[704]),
        .S(self_sf7[704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[705]),
        .S(self_sf7[705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[706]),
        .S(self_sf7[706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[707]),
        .S(self_sf7[707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[708]),
        .S(self_sf7[708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[709]),
        .S(self_sf7[709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[70].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[70]),
        .S(self_sf7[70]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[710]),
        .S(self_sf7[710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[711]),
        .S(self_sf7[711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[712]),
        .S(self_sf7[712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[713]),
        .S(self_sf7[713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[714]),
        .S(self_sf7[714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[715]),
        .S(self_sf7[715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[716]),
        .S(self_sf7[716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[717]),
        .S(self_sf7[717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[718]),
        .S(self_sf7[718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[719]),
        .S(self_sf7[719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[71].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[71]),
        .S(self_sf7[71]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[720]),
        .S(self_sf7[720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[721]),
        .S(self_sf7[721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[722]),
        .S(self_sf7[722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[723]),
        .S(self_sf7[723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[724]),
        .S(self_sf7[724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[725]),
        .S(self_sf7[725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[726]),
        .S(self_sf7[726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[727]),
        .S(self_sf7[727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[728]),
        .S(self_sf7[728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[729]),
        .S(self_sf7[729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[72].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[72]),
        .S(self_sf7[72]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[730]),
        .S(self_sf7[730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[731]),
        .S(self_sf7[731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[732]),
        .S(self_sf7[732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[733]),
        .S(self_sf7[733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[734]),
        .S(self_sf7[734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[735]),
        .S(self_sf7[735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[736]),
        .S(self_sf7[736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[737]),
        .S(self_sf7[737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[738]),
        .S(self_sf7[738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[739]),
        .S(self_sf7[739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[73].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[73]),
        .S(self_sf7[73]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[740]),
        .S(self_sf7[740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[741]),
        .S(self_sf7[741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[742]),
        .S(self_sf7[742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[743]),
        .S(self_sf7[743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[744]),
        .S(self_sf7[744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[745]),
        .S(self_sf7[745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[746]),
        .S(self_sf7[746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[747]),
        .S(self_sf7[747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[748]),
        .S(self_sf7[748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[749]),
        .S(self_sf7[749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[74].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[74]),
        .S(self_sf7[74]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[750]),
        .S(self_sf7[750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[751]),
        .S(self_sf7[751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[752]),
        .S(self_sf7[752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[753]),
        .S(self_sf7[753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[754]),
        .S(self_sf7[754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[755]),
        .S(self_sf7[755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[756]),
        .S(self_sf7[756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[757]),
        .S(self_sf7[757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[758]),
        .S(self_sf7[758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[759]),
        .S(self_sf7[759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[75].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[75]),
        .S(self_sf7[75]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[760]),
        .S(self_sf7[760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[761]),
        .S(self_sf7[761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[762]),
        .S(self_sf7[762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[763]),
        .S(self_sf7[763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[764]),
        .S(self_sf7[764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[765]),
        .S(self_sf7[765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[766]),
        .S(self_sf7[766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[767]),
        .S(self_sf7[767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[768]),
        .S(self_sf7[768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[769]),
        .S(self_sf7[769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[76].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[76]),
        .S(self_sf7[76]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[770]),
        .S(self_sf7[770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[771]),
        .S(self_sf7[771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[772]),
        .S(self_sf7[772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[773]),
        .S(self_sf7[773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[774]),
        .S(self_sf7[774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[775]),
        .S(self_sf7[775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[776]),
        .S(self_sf7[776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[777]),
        .S(self_sf7[777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[778]),
        .S(self_sf7[778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[779]),
        .S(self_sf7[779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[77].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[77]),
        .S(self_sf7[77]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[780]),
        .S(self_sf7[780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[781]),
        .S(self_sf7[781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[782]),
        .S(self_sf7[782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[783]),
        .S(self_sf7[783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[784]),
        .S(self_sf7[784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[785]),
        .S(self_sf7[785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[786]),
        .S(self_sf7[786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[787]),
        .S(self_sf7[787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[788]),
        .S(self_sf7[788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[789]),
        .S(self_sf7[789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[78].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[78]),
        .S(self_sf7[78]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[790]),
        .S(self_sf7[790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[791]),
        .S(self_sf7[791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[792]),
        .S(self_sf7[792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[793]),
        .S(self_sf7[793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[794]),
        .S(self_sf7[794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[795]),
        .S(self_sf7[795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[796]),
        .S(self_sf7[796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[797]),
        .S(self_sf7[797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[798]),
        .S(self_sf7[798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[799]),
        .S(self_sf7[799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[79].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[79]),
        .S(self_sf7[79]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[7].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[7]),
        .S(info_sf7[7]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[800].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[800]),
        .S(self_sf7[800]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[801].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[801]),
        .S(self_sf7[801]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[802].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[802]),
        .S(self_sf7[802]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[803].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[803]),
        .S(self_sf7[803]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[804].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[804]),
        .S(self_sf7[804]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[805].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[805]),
        .S(self_sf7[805]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[806].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[806]),
        .S(self_sf7[806]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[807].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[807]),
        .S(self_sf7[807]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[808].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[808]),
        .S(self_sf7[808]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[809].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[809]),
        .S(self_sf7[809]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[80].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[80]),
        .S(self_sf7[80]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[810].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[810]),
        .S(self_sf7[810]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[811].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[811]),
        .S(self_sf7[811]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[812].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[812]),
        .S(self_sf7[812]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[813].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[813]),
        .S(self_sf7[813]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[814].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[814]),
        .S(self_sf7[814]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[815].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[815]),
        .S(self_sf7[815]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[816].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[816]),
        .S(self_sf7[816]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[817].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[817]),
        .S(self_sf7[817]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[818].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[818]),
        .S(self_sf7[818]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[819].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[819]),
        .S(self_sf7[819]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[81].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[81]),
        .S(self_sf7[81]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[820].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[820]),
        .S(self_sf7[820]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[821].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[821]),
        .S(self_sf7[821]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[822].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[822]),
        .S(self_sf7[822]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[823].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[823]),
        .S(self_sf7[823]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[824].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[824]),
        .S(self_sf7[824]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[825].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[825]),
        .S(self_sf7[825]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[826].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[826]),
        .S(self_sf7[826]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[827].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[827]),
        .S(self_sf7[827]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[828].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[828]),
        .S(self_sf7[828]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[829].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[829]),
        .S(self_sf7[829]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[82].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[82]),
        .S(self_sf7[82]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[830].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[830]),
        .S(self_sf7[830]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[831].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[831]),
        .S(self_sf7[831]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[832].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[832]),
        .S(self_sf7[832]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[833].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[833]),
        .S(self_sf7[833]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[834].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[834]),
        .S(self_sf7[834]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[835].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[835]),
        .S(self_sf7[835]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[836].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[836]),
        .S(self_sf7[836]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[837].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[837]),
        .S(self_sf7[837]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[838].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[838]),
        .S(self_sf7[838]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[839].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[839]),
        .S(self_sf7[839]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[83].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[83]),
        .S(self_sf7[83]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[840].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[840]),
        .S(self_sf7[840]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[841].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[841]),
        .S(self_sf7[841]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[842].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[842]),
        .S(self_sf7[842]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[843].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[843]),
        .S(self_sf7[843]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[844].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[844]),
        .S(self_sf7[844]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[845].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[845]),
        .S(self_sf7[845]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[846].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[846]),
        .S(self_sf7[846]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[847].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[847]),
        .S(self_sf7[847]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[848].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[848]),
        .S(self_sf7[848]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[849].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[849]),
        .S(self_sf7[849]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[84].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[84]),
        .S(self_sf7[84]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[850].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[850]),
        .S(self_sf7[850]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[851].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[851]),
        .S(self_sf7[851]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[852].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[852]),
        .S(self_sf7[852]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[853].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[853]),
        .S(self_sf7[853]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[854].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[854]),
        .S(self_sf7[854]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[855].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[855]),
        .S(self_sf7[855]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[856].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[856]),
        .S(self_sf7[856]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[857].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[857]),
        .S(self_sf7[857]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[858].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[858]),
        .S(self_sf7[858]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[859].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[859]),
        .S(self_sf7[859]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[85].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[85]),
        .S(self_sf7[85]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[860].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[860]),
        .S(self_sf7[860]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[861].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[861]),
        .S(self_sf7[861]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[862].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[862]),
        .S(self_sf7[862]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[863].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[863]),
        .S(self_sf7[863]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[864].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[864]),
        .S(self_sf7[864]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[865].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[865]),
        .S(self_sf7[865]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[866].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[866]),
        .S(self_sf7[866]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[867].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[867]),
        .S(self_sf7[867]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[868].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[868]),
        .S(self_sf7[868]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[869].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[869]),
        .S(self_sf7[869]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[86].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[86]),
        .S(self_sf7[86]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[870].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[870]),
        .S(self_sf7[870]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[871].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[871]),
        .S(self_sf7[871]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[872].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[872]),
        .S(self_sf7[872]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[873].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[873]),
        .S(self_sf7[873]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[874].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[874]),
        .S(self_sf7[874]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[875].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[875]),
        .S(self_sf7[875]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[876].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[876]),
        .S(self_sf7[876]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[877].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[877]),
        .S(self_sf7[877]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[878].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[878]),
        .S(self_sf7[878]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[879].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[879]),
        .S(self_sf7[879]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[87].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[87]),
        .S(self_sf7[87]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[880].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[880]),
        .S(self_sf7[880]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[881].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[881]),
        .S(self_sf7[881]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[882].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[882]),
        .S(self_sf7[882]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[883].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[883]),
        .S(self_sf7[883]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[884].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[884]),
        .S(self_sf7[884]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[885].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[885]),
        .S(self_sf7[885]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[886].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[886]),
        .S(self_sf7[886]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[887].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[887]),
        .S(self_sf7[887]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[888].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[888]),
        .S(self_sf7[888]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[889].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[889]),
        .S(self_sf7[889]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[88].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[88]),
        .S(self_sf7[88]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[890].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[890]),
        .S(self_sf7[890]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[891].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[891]),
        .S(self_sf7[891]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[892].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[892]),
        .S(self_sf7[892]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[893].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[893]),
        .S(self_sf7[893]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[894].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[894]),
        .S(self_sf7[894]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[895].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[895]),
        .S(self_sf7[895]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[896].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[896]),
        .S(self_sf7[896]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[897].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[897]),
        .S(self_sf7[897]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[898].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[898]),
        .S(self_sf7[898]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[899].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[899]),
        .S(self_sf7[899]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[89].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[89]),
        .S(self_sf7[89]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[8].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[8]),
        .S(self_sf7[8]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[900].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[900]),
        .S(self_sf7[900]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[901].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[901]),
        .S(self_sf7[901]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[902].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[902]),
        .S(self_sf7[902]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[903].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[903]),
        .S(self_sf7[903]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[904].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[904]),
        .S(self_sf7[904]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[905].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[905]),
        .S(self_sf7[905]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[906].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[906]),
        .S(self_sf7[906]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[907].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[907]),
        .S(self_sf7[907]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[908].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[908]),
        .S(self_sf7[908]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[909].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[909]),
        .S(self_sf7[909]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[90].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[90]),
        .S(self_sf7[90]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[910].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[910]),
        .S(self_sf7[910]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[911].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[911]),
        .S(self_sf7[911]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[912].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[912]),
        .S(self_sf7[912]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[913].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[913]),
        .S(self_sf7[913]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[914].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[914]),
        .S(self_sf7[914]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[915].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[915]),
        .S(self_sf7[915]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[916].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[916]),
        .S(self_sf7[916]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[917].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[917]),
        .S(self_sf7[917]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[918].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[918]),
        .S(self_sf7[918]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[919].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[919]),
        .S(self_sf7[919]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[91].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[91]),
        .S(self_sf7[91]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[920].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[920]),
        .S(self_sf7[920]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[921].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[921]),
        .S(self_sf7[921]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[922].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[922]),
        .S(self_sf7[922]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[923].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[923]),
        .S(self_sf7[923]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[924].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[924]),
        .S(self_sf7[924]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[925].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[925]),
        .S(self_sf7[925]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[926].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[926]),
        .S(self_sf7[926]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[927].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[927]),
        .S(self_sf7[927]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[928].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[928]),
        .S(self_sf7[928]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[929].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[929]),
        .S(self_sf7[929]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[92].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[92]),
        .S(self_sf7[92]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[930].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[930]),
        .S(self_sf7[930]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[931].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[931]),
        .S(self_sf7[931]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[932].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[932]),
        .S(self_sf7[932]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[933].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[933]),
        .S(self_sf7[933]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[934].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[934]),
        .S(self_sf7[934]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[935].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[935]),
        .S(self_sf7[935]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[936].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[936]),
        .S(self_sf7[936]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[937].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[937]),
        .S(self_sf7[937]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[938].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[938]),
        .S(self_sf7[938]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[939].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[939]),
        .S(self_sf7[939]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[93].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[93]),
        .S(self_sf7[93]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[940].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[940]),
        .S(self_sf7[940]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[941].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[941]),
        .S(self_sf7[941]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[942].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[942]),
        .S(self_sf7[942]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[943].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[943]),
        .S(self_sf7[943]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[944].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[944]),
        .S(self_sf7[944]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[945].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[945]),
        .S(self_sf7[945]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[946].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[946]),
        .S(self_sf7[946]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[947].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[947]),
        .S(self_sf7[947]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[948].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[948]),
        .S(self_sf7[948]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[949].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[949]),
        .S(self_sf7[949]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[94].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[94]),
        .S(self_sf7[94]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[950].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[950]),
        .S(self_sf7[950]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[951].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[951]),
        .S(self_sf7[951]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[952].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[952]),
        .S(self_sf7[952]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[953].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[953]),
        .S(self_sf7[953]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[954].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[954]),
        .S(self_sf7[954]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[955].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[955]),
        .S(self_sf7[955]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[956].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[956]),
        .S(self_sf7[956]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[957].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[957]),
        .S(self_sf7[957]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[958].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[958]),
        .S(self_sf7[958]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[959].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[959]),
        .S(self_sf7[959]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[95].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[95]),
        .S(self_sf7[95]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[960].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[960]),
        .S(self_sf7[960]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[961].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[961]),
        .S(self_sf7[961]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[962].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[962]),
        .S(self_sf7[962]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[963].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[963]),
        .S(self_sf7[963]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[964].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[964]),
        .S(self_sf7[964]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[965].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[965]),
        .S(self_sf7[965]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[966].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[966]),
        .S(self_sf7[966]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[967].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[967]),
        .S(self_sf7[967]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[968].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[968]),
        .S(self_sf7[968]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[969].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[969]),
        .S(self_sf7[969]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[96].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[96]),
        .S(self_sf7[96]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[970].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[970]),
        .S(self_sf7[970]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[971].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[971]),
        .S(self_sf7[971]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[972].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[972]),
        .S(self_sf7[972]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[973].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[973]),
        .S(self_sf7[973]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[974].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[974]),
        .S(self_sf7[974]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[975].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[975]),
        .S(self_sf7[975]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[976].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[976]),
        .S(self_sf7[976]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[977].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[977]),
        .S(self_sf7[977]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[978].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[978]),
        .S(self_sf7[978]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[979].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[979]),
        .S(self_sf7[979]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[97].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[97]),
        .S(self_sf7[97]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[980].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[980]),
        .S(self_sf7[980]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[981].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[981]),
        .S(self_sf7[981]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[982].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[982]),
        .S(self_sf7[982]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[983].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[983]),
        .S(self_sf7[983]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[984].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[984]),
        .S(self_sf7[984]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[985].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[985]),
        .S(self_sf7[985]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[986].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[986]),
        .S(self_sf7[986]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[987].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[987]),
        .S(self_sf7[987]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[988].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[988]),
        .S(self_sf7[988]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[989].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[989]),
        .S(self_sf7[989]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[98].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[98]),
        .S(self_sf7[98]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[990].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[990]),
        .S(self_sf7[990]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[991].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[991]),
        .S(self_sf7[991]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[992].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[992]),
        .S(self_sf7[992]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[993].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[993]),
        .S(self_sf7[993]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[994].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[994]),
        .S(self_sf7[994]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[995].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[995]),
        .S(self_sf7[995]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[996].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[996]),
        .S(self_sf7[996]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[997].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[997]),
        .S(self_sf7[997]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[998].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[998]),
        .S(self_sf7[998]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[999].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[999]),
        .S(self_sf7[999]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[99].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[99]),
        .S(self_sf7[99]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[9].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[9]),
        .S(self_sf7[9]));
  (* BOX_TYPE = "black_box" *) 
  MUXF8 \activity_ROsf8[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf8[0]),
        .S(self_sf8[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF9 \activity_ROsf9[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf9[0]),
        .S(self_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_0
       (.I0(1'b0),
        .O(self_sf7[1802]));
  LUT1 #(
    .INIT(2'h2)) 
    i_1
       (.I0(1'b0),
        .O(self_sf7[1801]));
  LUT1 #(
    .INIT(2'h2)) 
    i_10
       (.I0(1'b0),
        .O(info_sf8[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_11
       (.I0(1'b0),
        .O(info_sf8[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_12
       (.I0(1'b0),
        .O(info_sf8[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_13
       (.I0(1'b0),
        .O(info_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_14
       (.I0(1'b0),
        .O(info_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_15
       (.I0(1'b0),
        .O(info_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_16
       (.I0(1'b0),
        .O(info_sf8[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_17
       (.I0(1'b0),
        .O(info_sf9[7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_18
       (.I0(1'b0),
        .O(info_sf9[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_19
       (.I0(1'b0),
        .O(info_sf9[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_2
       (.I0(1'b0),
        .O(self_sf7[1800]));
  LUT1 #(
    .INIT(2'h2)) 
    i_20
       (.I0(1'b0),
        .O(info_sf9[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_21
       (.I0(1'b0),
        .O(info_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_22
       (.I0(1'b0),
        .O(info_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_23
       (.I0(1'b0),
        .O(info_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_24
       (.I0(1'b0),
        .O(info_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_3
       (.I0(1'b0),
        .O(self_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_4
       (.I0(1'b0),
        .O(self_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_5
       (.I0(1'b0),
        .O(self_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_6
       (.I0(1'b0),
        .O(self_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_7
       (.I0(1'b0),
        .O(self_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_8
       (.I0(1'b0),
        .O(self_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_9
       (.I0(1'b0),
        .O(info_sf8[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst
       (.I0(self_sf7[7]),
        .O(info_sf7[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__0
       (.I0(self_sf7[6]),
        .O(info_sf7[6]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__1
       (.I0(self_sf7[5]),
        .O(info_sf7[5]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__2
       (.I0(self_sf7[4]),
        .O(info_sf7[4]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__3
       (.I0(self_sf7[3]),
        .O(info_sf7[3]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__4
       (.I0(self_sf7[2]),
        .O(info_sf7[2]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__5
       (.I0(self_sf7[1]),
        .O(info_sf7[1]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__6
       (.I0(self_sf7[0]),
        .O(info_sf7[0]));
endmodule

(* ORIG_REF_NAME = "muxer" *) (* box_type = "black_box" *) (* dont_touch = "true" *) 
module switch_elements_muxer__2
   (enable_i,
    info_o);
  input enable_i;
  output info_o;

  wire enable_i;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf7;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf8;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf9;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [1802:0]self_sf7;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf8;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf9;

  assign info_o = info_sf7[1];
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[0]),
        .S(info_sf7[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1000].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1000]),
        .S(self_sf7[1000]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1001].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1001]),
        .S(self_sf7[1001]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1002].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1002]),
        .S(self_sf7[1002]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1003].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1003]),
        .S(self_sf7[1003]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1004].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1004]),
        .S(self_sf7[1004]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1005].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1005]),
        .S(self_sf7[1005]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1006].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1006]),
        .S(self_sf7[1006]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1007].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1007]),
        .S(self_sf7[1007]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1008].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1008]),
        .S(self_sf7[1008]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1009].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1009]),
        .S(self_sf7[1009]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[100]),
        .S(self_sf7[100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1010].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1010]),
        .S(self_sf7[1010]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1011].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1011]),
        .S(self_sf7[1011]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1012].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1012]),
        .S(self_sf7[1012]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1013].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1013]),
        .S(self_sf7[1013]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1014].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1014]),
        .S(self_sf7[1014]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1015].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1015]),
        .S(self_sf7[1015]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1016].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1016]),
        .S(self_sf7[1016]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1017].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1017]),
        .S(self_sf7[1017]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1018].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1018]),
        .S(self_sf7[1018]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1019].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1019]),
        .S(self_sf7[1019]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[101]),
        .S(self_sf7[101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1020].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1020]),
        .S(self_sf7[1020]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1021].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1021]),
        .S(self_sf7[1021]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1022].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1022]),
        .S(self_sf7[1022]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1023].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1023]),
        .S(self_sf7[1023]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1024].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1024]),
        .S(self_sf7[1024]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1025].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1025]),
        .S(self_sf7[1025]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1026].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1026]),
        .S(self_sf7[1026]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1027].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1027]),
        .S(self_sf7[1027]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1028].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1028]),
        .S(self_sf7[1028]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1029].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1029]),
        .S(self_sf7[1029]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[102]),
        .S(self_sf7[102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1030].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1030]),
        .S(self_sf7[1030]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1031].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1031]),
        .S(self_sf7[1031]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1032].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1032]),
        .S(self_sf7[1032]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1033].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1033]),
        .S(self_sf7[1033]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1034].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1034]),
        .S(self_sf7[1034]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1035].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1035]),
        .S(self_sf7[1035]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1036].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1036]),
        .S(self_sf7[1036]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1037].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1037]),
        .S(self_sf7[1037]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1038].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1038]),
        .S(self_sf7[1038]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1039].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1039]),
        .S(self_sf7[1039]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[103]),
        .S(self_sf7[103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1040].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1040]),
        .S(self_sf7[1040]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1041].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1041]),
        .S(self_sf7[1041]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1042].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1042]),
        .S(self_sf7[1042]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1043].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1043]),
        .S(self_sf7[1043]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1044].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1044]),
        .S(self_sf7[1044]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1045].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1045]),
        .S(self_sf7[1045]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1046].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1046]),
        .S(self_sf7[1046]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1047].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1047]),
        .S(self_sf7[1047]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1048].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1048]),
        .S(self_sf7[1048]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1049].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1049]),
        .S(self_sf7[1049]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[104]),
        .S(self_sf7[104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1050].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1050]),
        .S(self_sf7[1050]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1051].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1051]),
        .S(self_sf7[1051]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1052].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1052]),
        .S(self_sf7[1052]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1053].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1053]),
        .S(self_sf7[1053]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1054].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1054]),
        .S(self_sf7[1054]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1055].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1055]),
        .S(self_sf7[1055]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1056].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1056]),
        .S(self_sf7[1056]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1057].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1057]),
        .S(self_sf7[1057]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1058].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1058]),
        .S(self_sf7[1058]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1059].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1059]),
        .S(self_sf7[1059]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[105]),
        .S(self_sf7[105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1060].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1060]),
        .S(self_sf7[1060]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1061].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1061]),
        .S(self_sf7[1061]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1062].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1062]),
        .S(self_sf7[1062]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1063].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1063]),
        .S(self_sf7[1063]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1064].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1064]),
        .S(self_sf7[1064]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1065].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1065]),
        .S(self_sf7[1065]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1066].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1066]),
        .S(self_sf7[1066]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1067].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1067]),
        .S(self_sf7[1067]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1068].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1068]),
        .S(self_sf7[1068]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1069].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1069]),
        .S(self_sf7[1069]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[106]),
        .S(self_sf7[106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1070].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1070]),
        .S(self_sf7[1070]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1071].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1071]),
        .S(self_sf7[1071]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1072].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1072]),
        .S(self_sf7[1072]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1073].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1073]),
        .S(self_sf7[1073]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1074].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1074]),
        .S(self_sf7[1074]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1075].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1075]),
        .S(self_sf7[1075]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1076].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1076]),
        .S(self_sf7[1076]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1077].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1077]),
        .S(self_sf7[1077]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1078].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1078]),
        .S(self_sf7[1078]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1079].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1079]),
        .S(self_sf7[1079]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[107]),
        .S(self_sf7[107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1080].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1080]),
        .S(self_sf7[1080]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1081].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1081]),
        .S(self_sf7[1081]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1082].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1082]),
        .S(self_sf7[1082]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1083].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1083]),
        .S(self_sf7[1083]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1084].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1084]),
        .S(self_sf7[1084]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1085].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1085]),
        .S(self_sf7[1085]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1086].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1086]),
        .S(self_sf7[1086]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1087].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1087]),
        .S(self_sf7[1087]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1088].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1088]),
        .S(self_sf7[1088]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1089].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1089]),
        .S(self_sf7[1089]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[108]),
        .S(self_sf7[108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1090].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1090]),
        .S(self_sf7[1090]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1091].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1091]),
        .S(self_sf7[1091]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1092].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1092]),
        .S(self_sf7[1092]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1093].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1093]),
        .S(self_sf7[1093]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1094].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1094]),
        .S(self_sf7[1094]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1095].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1095]),
        .S(self_sf7[1095]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1096].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1096]),
        .S(self_sf7[1096]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1097].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1097]),
        .S(self_sf7[1097]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1098].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1098]),
        .S(self_sf7[1098]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1099].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1099]),
        .S(self_sf7[1099]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[109]),
        .S(self_sf7[109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[10].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[10]),
        .S(self_sf7[10]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1100]),
        .S(self_sf7[1100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1101]),
        .S(self_sf7[1101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1102]),
        .S(self_sf7[1102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1103]),
        .S(self_sf7[1103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1104]),
        .S(self_sf7[1104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1105]),
        .S(self_sf7[1105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1106]),
        .S(self_sf7[1106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1107]),
        .S(self_sf7[1107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1108]),
        .S(self_sf7[1108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1109]),
        .S(self_sf7[1109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[110]),
        .S(self_sf7[110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1110]),
        .S(self_sf7[1110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1111]),
        .S(self_sf7[1111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1112]),
        .S(self_sf7[1112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1113]),
        .S(self_sf7[1113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1114]),
        .S(self_sf7[1114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1115]),
        .S(self_sf7[1115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1116]),
        .S(self_sf7[1116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1117]),
        .S(self_sf7[1117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1118]),
        .S(self_sf7[1118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1119]),
        .S(self_sf7[1119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[111]),
        .S(self_sf7[111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1120]),
        .S(self_sf7[1120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1121]),
        .S(self_sf7[1121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1122]),
        .S(self_sf7[1122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1123]),
        .S(self_sf7[1123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1124]),
        .S(self_sf7[1124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1125]),
        .S(self_sf7[1125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1126]),
        .S(self_sf7[1126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1127]),
        .S(self_sf7[1127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1128]),
        .S(self_sf7[1128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1129]),
        .S(self_sf7[1129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[112]),
        .S(self_sf7[112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1130]),
        .S(self_sf7[1130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1131]),
        .S(self_sf7[1131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1132]),
        .S(self_sf7[1132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1133]),
        .S(self_sf7[1133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1134]),
        .S(self_sf7[1134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1135]),
        .S(self_sf7[1135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1136]),
        .S(self_sf7[1136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1137]),
        .S(self_sf7[1137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1138]),
        .S(self_sf7[1138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1139]),
        .S(self_sf7[1139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[113]),
        .S(self_sf7[113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1140]),
        .S(self_sf7[1140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1141]),
        .S(self_sf7[1141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1142]),
        .S(self_sf7[1142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1143]),
        .S(self_sf7[1143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1144]),
        .S(self_sf7[1144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1145]),
        .S(self_sf7[1145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1146]),
        .S(self_sf7[1146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1147]),
        .S(self_sf7[1147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1148]),
        .S(self_sf7[1148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1149]),
        .S(self_sf7[1149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[114]),
        .S(self_sf7[114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1150]),
        .S(self_sf7[1150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1151]),
        .S(self_sf7[1151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1152]),
        .S(self_sf7[1152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1153]),
        .S(self_sf7[1153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1154]),
        .S(self_sf7[1154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1155]),
        .S(self_sf7[1155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1156]),
        .S(self_sf7[1156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1157]),
        .S(self_sf7[1157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1158]),
        .S(self_sf7[1158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1159]),
        .S(self_sf7[1159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[115]),
        .S(self_sf7[115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1160]),
        .S(self_sf7[1160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1161]),
        .S(self_sf7[1161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1162]),
        .S(self_sf7[1162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1163]),
        .S(self_sf7[1163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1164]),
        .S(self_sf7[1164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1165]),
        .S(self_sf7[1165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1166]),
        .S(self_sf7[1166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1167]),
        .S(self_sf7[1167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1168]),
        .S(self_sf7[1168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1169]),
        .S(self_sf7[1169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[116]),
        .S(self_sf7[116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1170]),
        .S(self_sf7[1170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1171]),
        .S(self_sf7[1171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1172]),
        .S(self_sf7[1172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1173]),
        .S(self_sf7[1173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1174]),
        .S(self_sf7[1174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1175]),
        .S(self_sf7[1175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1176]),
        .S(self_sf7[1176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1177]),
        .S(self_sf7[1177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1178]),
        .S(self_sf7[1178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1179]),
        .S(self_sf7[1179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[117]),
        .S(self_sf7[117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1180]),
        .S(self_sf7[1180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1181]),
        .S(self_sf7[1181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1182]),
        .S(self_sf7[1182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1183]),
        .S(self_sf7[1183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1184]),
        .S(self_sf7[1184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1185]),
        .S(self_sf7[1185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1186]),
        .S(self_sf7[1186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1187]),
        .S(self_sf7[1187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1188]),
        .S(self_sf7[1188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1189]),
        .S(self_sf7[1189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[118]),
        .S(self_sf7[118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1190]),
        .S(self_sf7[1190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1191]),
        .S(self_sf7[1191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1192]),
        .S(self_sf7[1192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1193]),
        .S(self_sf7[1193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1194]),
        .S(self_sf7[1194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1195]),
        .S(self_sf7[1195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1196]),
        .S(self_sf7[1196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1197]),
        .S(self_sf7[1197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1198]),
        .S(self_sf7[1198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1199]),
        .S(self_sf7[1199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[119]),
        .S(self_sf7[119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[11].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[11]),
        .S(self_sf7[11]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1200]),
        .S(self_sf7[1200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1201]),
        .S(self_sf7[1201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1202]),
        .S(self_sf7[1202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1203]),
        .S(self_sf7[1203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1204]),
        .S(self_sf7[1204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1205]),
        .S(self_sf7[1205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1206]),
        .S(self_sf7[1206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1207]),
        .S(self_sf7[1207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1208]),
        .S(self_sf7[1208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1209]),
        .S(self_sf7[1209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[120]),
        .S(self_sf7[120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1210]),
        .S(self_sf7[1210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1211]),
        .S(self_sf7[1211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1212]),
        .S(self_sf7[1212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1213]),
        .S(self_sf7[1213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1214]),
        .S(self_sf7[1214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1215]),
        .S(self_sf7[1215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1216]),
        .S(self_sf7[1216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1217]),
        .S(self_sf7[1217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1218]),
        .S(self_sf7[1218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1219]),
        .S(self_sf7[1219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[121]),
        .S(self_sf7[121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1220]),
        .S(self_sf7[1220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1221]),
        .S(self_sf7[1221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1222]),
        .S(self_sf7[1222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1223]),
        .S(self_sf7[1223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1224]),
        .S(self_sf7[1224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1225]),
        .S(self_sf7[1225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1226]),
        .S(self_sf7[1226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1227]),
        .S(self_sf7[1227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1228]),
        .S(self_sf7[1228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1229]),
        .S(self_sf7[1229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[122]),
        .S(self_sf7[122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1230]),
        .S(self_sf7[1230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1231]),
        .S(self_sf7[1231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1232]),
        .S(self_sf7[1232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1233]),
        .S(self_sf7[1233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1234]),
        .S(self_sf7[1234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1235]),
        .S(self_sf7[1235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1236]),
        .S(self_sf7[1236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1237]),
        .S(self_sf7[1237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1238]),
        .S(self_sf7[1238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1239]),
        .S(self_sf7[1239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[123]),
        .S(self_sf7[123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1240]),
        .S(self_sf7[1240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1241]),
        .S(self_sf7[1241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1242]),
        .S(self_sf7[1242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1243]),
        .S(self_sf7[1243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1244]),
        .S(self_sf7[1244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1245]),
        .S(self_sf7[1245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1246]),
        .S(self_sf7[1246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1247]),
        .S(self_sf7[1247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1248]),
        .S(self_sf7[1248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1249]),
        .S(self_sf7[1249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[124]),
        .S(self_sf7[124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1250]),
        .S(self_sf7[1250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1251]),
        .S(self_sf7[1251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1252]),
        .S(self_sf7[1252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1253]),
        .S(self_sf7[1253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1254]),
        .S(self_sf7[1254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1255]),
        .S(self_sf7[1255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1256]),
        .S(self_sf7[1256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1257]),
        .S(self_sf7[1257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1258]),
        .S(self_sf7[1258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1259]),
        .S(self_sf7[1259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[125]),
        .S(self_sf7[125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1260]),
        .S(self_sf7[1260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1261]),
        .S(self_sf7[1261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1262]),
        .S(self_sf7[1262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1263]),
        .S(self_sf7[1263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1264]),
        .S(self_sf7[1264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1265]),
        .S(self_sf7[1265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1266]),
        .S(self_sf7[1266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1267]),
        .S(self_sf7[1267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1268]),
        .S(self_sf7[1268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1269]),
        .S(self_sf7[1269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[126]),
        .S(self_sf7[126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1270]),
        .S(self_sf7[1270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1271]),
        .S(self_sf7[1271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1272]),
        .S(self_sf7[1272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1273]),
        .S(self_sf7[1273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1274]),
        .S(self_sf7[1274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1275]),
        .S(self_sf7[1275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1276]),
        .S(self_sf7[1276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1277]),
        .S(self_sf7[1277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1278]),
        .S(self_sf7[1278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1279]),
        .S(self_sf7[1279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[127]),
        .S(self_sf7[127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1280]),
        .S(self_sf7[1280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1281]),
        .S(self_sf7[1281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1282]),
        .S(self_sf7[1282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1283]),
        .S(self_sf7[1283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1284]),
        .S(self_sf7[1284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1285]),
        .S(self_sf7[1285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1286]),
        .S(self_sf7[1286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1287]),
        .S(self_sf7[1287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1288]),
        .S(self_sf7[1288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1289]),
        .S(self_sf7[1289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[128]),
        .S(self_sf7[128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1290]),
        .S(self_sf7[1290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1291]),
        .S(self_sf7[1291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1292]),
        .S(self_sf7[1292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1293]),
        .S(self_sf7[1293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1294]),
        .S(self_sf7[1294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1295]),
        .S(self_sf7[1295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1296]),
        .S(self_sf7[1296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1297]),
        .S(self_sf7[1297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1298]),
        .S(self_sf7[1298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1299]),
        .S(self_sf7[1299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[129]),
        .S(self_sf7[129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[12].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[12]),
        .S(self_sf7[12]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1300]),
        .S(self_sf7[1300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1301]),
        .S(self_sf7[1301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1302]),
        .S(self_sf7[1302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1303]),
        .S(self_sf7[1303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1304]),
        .S(self_sf7[1304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1305]),
        .S(self_sf7[1305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1306]),
        .S(self_sf7[1306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1307]),
        .S(self_sf7[1307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1308]),
        .S(self_sf7[1308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1309]),
        .S(self_sf7[1309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[130]),
        .S(self_sf7[130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1310]),
        .S(self_sf7[1310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1311]),
        .S(self_sf7[1311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1312]),
        .S(self_sf7[1312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1313]),
        .S(self_sf7[1313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1314]),
        .S(self_sf7[1314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1315]),
        .S(self_sf7[1315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1316]),
        .S(self_sf7[1316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1317]),
        .S(self_sf7[1317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1318]),
        .S(self_sf7[1318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1319]),
        .S(self_sf7[1319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[131]),
        .S(self_sf7[131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1320]),
        .S(self_sf7[1320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1321]),
        .S(self_sf7[1321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1322]),
        .S(self_sf7[1322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1323]),
        .S(self_sf7[1323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1324]),
        .S(self_sf7[1324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1325]),
        .S(self_sf7[1325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1326]),
        .S(self_sf7[1326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1327]),
        .S(self_sf7[1327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1328]),
        .S(self_sf7[1328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1329]),
        .S(self_sf7[1329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[132]),
        .S(self_sf7[132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1330]),
        .S(self_sf7[1330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1331]),
        .S(self_sf7[1331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1332]),
        .S(self_sf7[1332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1333]),
        .S(self_sf7[1333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1334]),
        .S(self_sf7[1334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1335]),
        .S(self_sf7[1335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1336]),
        .S(self_sf7[1336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1337]),
        .S(self_sf7[1337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1338]),
        .S(self_sf7[1338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1339]),
        .S(self_sf7[1339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[133]),
        .S(self_sf7[133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1340]),
        .S(self_sf7[1340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1341]),
        .S(self_sf7[1341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1342]),
        .S(self_sf7[1342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1343]),
        .S(self_sf7[1343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1344]),
        .S(self_sf7[1344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1345]),
        .S(self_sf7[1345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1346]),
        .S(self_sf7[1346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1347]),
        .S(self_sf7[1347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1348]),
        .S(self_sf7[1348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1349]),
        .S(self_sf7[1349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[134]),
        .S(self_sf7[134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1350]),
        .S(self_sf7[1350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1351]),
        .S(self_sf7[1351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1352]),
        .S(self_sf7[1352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1353]),
        .S(self_sf7[1353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1354]),
        .S(self_sf7[1354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1355]),
        .S(self_sf7[1355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1356]),
        .S(self_sf7[1356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1357]),
        .S(self_sf7[1357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1358]),
        .S(self_sf7[1358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1359]),
        .S(self_sf7[1359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[135]),
        .S(self_sf7[135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1360]),
        .S(self_sf7[1360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1361]),
        .S(self_sf7[1361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1362]),
        .S(self_sf7[1362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1363]),
        .S(self_sf7[1363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1364]),
        .S(self_sf7[1364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1365]),
        .S(self_sf7[1365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1366]),
        .S(self_sf7[1366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1367]),
        .S(self_sf7[1367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1368]),
        .S(self_sf7[1368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1369]),
        .S(self_sf7[1369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[136]),
        .S(self_sf7[136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1370]),
        .S(self_sf7[1370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1371]),
        .S(self_sf7[1371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1372]),
        .S(self_sf7[1372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1373]),
        .S(self_sf7[1373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1374]),
        .S(self_sf7[1374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1375]),
        .S(self_sf7[1375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1376]),
        .S(self_sf7[1376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1377]),
        .S(self_sf7[1377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1378]),
        .S(self_sf7[1378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1379]),
        .S(self_sf7[1379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[137]),
        .S(self_sf7[137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1380]),
        .S(self_sf7[1380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1381]),
        .S(self_sf7[1381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1382]),
        .S(self_sf7[1382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1383]),
        .S(self_sf7[1383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1384]),
        .S(self_sf7[1384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1385]),
        .S(self_sf7[1385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1386]),
        .S(self_sf7[1386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1387]),
        .S(self_sf7[1387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1388]),
        .S(self_sf7[1388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1389]),
        .S(self_sf7[1389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[138]),
        .S(self_sf7[138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1390]),
        .S(self_sf7[1390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1391]),
        .S(self_sf7[1391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1392]),
        .S(self_sf7[1392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1393]),
        .S(self_sf7[1393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1394]),
        .S(self_sf7[1394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1395]),
        .S(self_sf7[1395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1396]),
        .S(self_sf7[1396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1397]),
        .S(self_sf7[1397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1398]),
        .S(self_sf7[1398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1399]),
        .S(self_sf7[1399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[139]),
        .S(self_sf7[139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[13].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[13]),
        .S(self_sf7[13]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1400]),
        .S(self_sf7[1400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1401]),
        .S(self_sf7[1401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1402]),
        .S(self_sf7[1402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1403]),
        .S(self_sf7[1403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1404]),
        .S(self_sf7[1404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1405]),
        .S(self_sf7[1405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1406]),
        .S(self_sf7[1406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1407]),
        .S(self_sf7[1407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1408]),
        .S(self_sf7[1408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1409]),
        .S(self_sf7[1409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[140]),
        .S(self_sf7[140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1410]),
        .S(self_sf7[1410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1411]),
        .S(self_sf7[1411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1412]),
        .S(self_sf7[1412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1413]),
        .S(self_sf7[1413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1414]),
        .S(self_sf7[1414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1415]),
        .S(self_sf7[1415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1416]),
        .S(self_sf7[1416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1417]),
        .S(self_sf7[1417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1418]),
        .S(self_sf7[1418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1419]),
        .S(self_sf7[1419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[141]),
        .S(self_sf7[141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1420]),
        .S(self_sf7[1420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1421]),
        .S(self_sf7[1421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1422]),
        .S(self_sf7[1422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1423]),
        .S(self_sf7[1423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1424]),
        .S(self_sf7[1424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1425]),
        .S(self_sf7[1425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1426]),
        .S(self_sf7[1426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1427]),
        .S(self_sf7[1427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1428]),
        .S(self_sf7[1428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1429]),
        .S(self_sf7[1429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[142]),
        .S(self_sf7[142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1430]),
        .S(self_sf7[1430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1431]),
        .S(self_sf7[1431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1432]),
        .S(self_sf7[1432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1433]),
        .S(self_sf7[1433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1434]),
        .S(self_sf7[1434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1435]),
        .S(self_sf7[1435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1436]),
        .S(self_sf7[1436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1437]),
        .S(self_sf7[1437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1438]),
        .S(self_sf7[1438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1439]),
        .S(self_sf7[1439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[143]),
        .S(self_sf7[143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1440]),
        .S(self_sf7[1440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1441]),
        .S(self_sf7[1441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1442]),
        .S(self_sf7[1442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1443]),
        .S(self_sf7[1443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1444]),
        .S(self_sf7[1444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1445]),
        .S(self_sf7[1445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1446]),
        .S(self_sf7[1446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1447]),
        .S(self_sf7[1447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1448]),
        .S(self_sf7[1448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1449]),
        .S(self_sf7[1449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[144]),
        .S(self_sf7[144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1450]),
        .S(self_sf7[1450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1451]),
        .S(self_sf7[1451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1452]),
        .S(self_sf7[1452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1453]),
        .S(self_sf7[1453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1454]),
        .S(self_sf7[1454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1455]),
        .S(self_sf7[1455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1456]),
        .S(self_sf7[1456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1457]),
        .S(self_sf7[1457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1458]),
        .S(self_sf7[1458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1459]),
        .S(self_sf7[1459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[145]),
        .S(self_sf7[145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1460]),
        .S(self_sf7[1460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1461]),
        .S(self_sf7[1461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1462]),
        .S(self_sf7[1462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1463]),
        .S(self_sf7[1463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1464]),
        .S(self_sf7[1464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1465]),
        .S(self_sf7[1465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1466]),
        .S(self_sf7[1466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1467]),
        .S(self_sf7[1467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1468]),
        .S(self_sf7[1468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1469]),
        .S(self_sf7[1469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[146]),
        .S(self_sf7[146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1470]),
        .S(self_sf7[1470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1471]),
        .S(self_sf7[1471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1472]),
        .S(self_sf7[1472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1473]),
        .S(self_sf7[1473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1474]),
        .S(self_sf7[1474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1475]),
        .S(self_sf7[1475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1476]),
        .S(self_sf7[1476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1477]),
        .S(self_sf7[1477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1478]),
        .S(self_sf7[1478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1479]),
        .S(self_sf7[1479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[147]),
        .S(self_sf7[147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1480]),
        .S(self_sf7[1480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1481]),
        .S(self_sf7[1481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1482]),
        .S(self_sf7[1482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1483]),
        .S(self_sf7[1483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1484]),
        .S(self_sf7[1484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1485]),
        .S(self_sf7[1485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1486]),
        .S(self_sf7[1486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1487]),
        .S(self_sf7[1487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1488]),
        .S(self_sf7[1488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1489]),
        .S(self_sf7[1489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[148]),
        .S(self_sf7[148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1490]),
        .S(self_sf7[1490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1491]),
        .S(self_sf7[1491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1492]),
        .S(self_sf7[1492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1493]),
        .S(self_sf7[1493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1494]),
        .S(self_sf7[1494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1495]),
        .S(self_sf7[1495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1496]),
        .S(self_sf7[1496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1497]),
        .S(self_sf7[1497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1498]),
        .S(self_sf7[1498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1499]),
        .S(self_sf7[1499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[149]),
        .S(self_sf7[149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[14].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[14]),
        .S(self_sf7[14]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1500]),
        .S(self_sf7[1500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1501]),
        .S(self_sf7[1501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1502]),
        .S(self_sf7[1502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1503]),
        .S(self_sf7[1503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1504]),
        .S(self_sf7[1504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1505]),
        .S(self_sf7[1505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1506]),
        .S(self_sf7[1506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1507]),
        .S(self_sf7[1507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1508]),
        .S(self_sf7[1508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1509]),
        .S(self_sf7[1509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[150]),
        .S(self_sf7[150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1510]),
        .S(self_sf7[1510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1511]),
        .S(self_sf7[1511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1512]),
        .S(self_sf7[1512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1513]),
        .S(self_sf7[1513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1514]),
        .S(self_sf7[1514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1515]),
        .S(self_sf7[1515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1516]),
        .S(self_sf7[1516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1517]),
        .S(self_sf7[1517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1518]),
        .S(self_sf7[1518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1519]),
        .S(self_sf7[1519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[151]),
        .S(self_sf7[151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1520]),
        .S(self_sf7[1520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1521]),
        .S(self_sf7[1521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1522]),
        .S(self_sf7[1522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1523]),
        .S(self_sf7[1523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1524]),
        .S(self_sf7[1524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1525]),
        .S(self_sf7[1525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1526]),
        .S(self_sf7[1526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1527]),
        .S(self_sf7[1527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1528]),
        .S(self_sf7[1528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1529]),
        .S(self_sf7[1529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[152]),
        .S(self_sf7[152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1530]),
        .S(self_sf7[1530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1531]),
        .S(self_sf7[1531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1532]),
        .S(self_sf7[1532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1533]),
        .S(self_sf7[1533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1534]),
        .S(self_sf7[1534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1535]),
        .S(self_sf7[1535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1536]),
        .S(self_sf7[1536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1537]),
        .S(self_sf7[1537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1538]),
        .S(self_sf7[1538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1539]),
        .S(self_sf7[1539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[153]),
        .S(self_sf7[153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1540]),
        .S(self_sf7[1540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1541]),
        .S(self_sf7[1541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1542]),
        .S(self_sf7[1542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1543]),
        .S(self_sf7[1543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1544]),
        .S(self_sf7[1544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1545]),
        .S(self_sf7[1545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1546]),
        .S(self_sf7[1546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1547]),
        .S(self_sf7[1547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1548]),
        .S(self_sf7[1548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1549]),
        .S(self_sf7[1549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[154]),
        .S(self_sf7[154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1550]),
        .S(self_sf7[1550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1551]),
        .S(self_sf7[1551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1552]),
        .S(self_sf7[1552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1553]),
        .S(self_sf7[1553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1554]),
        .S(self_sf7[1554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1555]),
        .S(self_sf7[1555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1556]),
        .S(self_sf7[1556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1557]),
        .S(self_sf7[1557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1558]),
        .S(self_sf7[1558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1559]),
        .S(self_sf7[1559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[155]),
        .S(self_sf7[155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1560]),
        .S(self_sf7[1560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1561]),
        .S(self_sf7[1561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1562]),
        .S(self_sf7[1562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1563]),
        .S(self_sf7[1563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1564]),
        .S(self_sf7[1564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1565]),
        .S(self_sf7[1565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1566]),
        .S(self_sf7[1566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1567]),
        .S(self_sf7[1567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1568]),
        .S(self_sf7[1568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1569]),
        .S(self_sf7[1569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[156]),
        .S(self_sf7[156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1570]),
        .S(self_sf7[1570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1571]),
        .S(self_sf7[1571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1572]),
        .S(self_sf7[1572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1573]),
        .S(self_sf7[1573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1574]),
        .S(self_sf7[1574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1575]),
        .S(self_sf7[1575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1576]),
        .S(self_sf7[1576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1577]),
        .S(self_sf7[1577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1578]),
        .S(self_sf7[1578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1579]),
        .S(self_sf7[1579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[157]),
        .S(self_sf7[157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1580]),
        .S(self_sf7[1580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1581]),
        .S(self_sf7[1581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1582]),
        .S(self_sf7[1582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1583]),
        .S(self_sf7[1583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1584]),
        .S(self_sf7[1584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1585]),
        .S(self_sf7[1585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1586]),
        .S(self_sf7[1586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1587]),
        .S(self_sf7[1587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1588]),
        .S(self_sf7[1588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1589]),
        .S(self_sf7[1589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[158]),
        .S(self_sf7[158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1590]),
        .S(self_sf7[1590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1591]),
        .S(self_sf7[1591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1592]),
        .S(self_sf7[1592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1593]),
        .S(self_sf7[1593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1594]),
        .S(self_sf7[1594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1595]),
        .S(self_sf7[1595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1596]),
        .S(self_sf7[1596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1597]),
        .S(self_sf7[1597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1598]),
        .S(self_sf7[1598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1599]),
        .S(self_sf7[1599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[159]),
        .S(self_sf7[159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[15].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[15]),
        .S(self_sf7[15]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1600]),
        .S(self_sf7[1600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1601]),
        .S(self_sf7[1601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1602]),
        .S(self_sf7[1602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1603]),
        .S(self_sf7[1603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1604]),
        .S(self_sf7[1604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1605]),
        .S(self_sf7[1605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1606]),
        .S(self_sf7[1606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1607]),
        .S(self_sf7[1607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1608]),
        .S(self_sf7[1608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1609]),
        .S(self_sf7[1609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[160]),
        .S(self_sf7[160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1610]),
        .S(self_sf7[1610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1611]),
        .S(self_sf7[1611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1612]),
        .S(self_sf7[1612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1613]),
        .S(self_sf7[1613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1614]),
        .S(self_sf7[1614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1615]),
        .S(self_sf7[1615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1616]),
        .S(self_sf7[1616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1617]),
        .S(self_sf7[1617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1618]),
        .S(self_sf7[1618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1619]),
        .S(self_sf7[1619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[161]),
        .S(self_sf7[161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1620]),
        .S(self_sf7[1620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1621]),
        .S(self_sf7[1621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1622]),
        .S(self_sf7[1622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1623]),
        .S(self_sf7[1623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1624]),
        .S(self_sf7[1624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1625]),
        .S(self_sf7[1625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1626]),
        .S(self_sf7[1626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1627]),
        .S(self_sf7[1627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1628]),
        .S(self_sf7[1628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1629]),
        .S(self_sf7[1629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[162]),
        .S(self_sf7[162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1630]),
        .S(self_sf7[1630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1631]),
        .S(self_sf7[1631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1632]),
        .S(self_sf7[1632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1633]),
        .S(self_sf7[1633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1634]),
        .S(self_sf7[1634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1635]),
        .S(self_sf7[1635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1636]),
        .S(self_sf7[1636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1637]),
        .S(self_sf7[1637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1638]),
        .S(self_sf7[1638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1639]),
        .S(self_sf7[1639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[163]),
        .S(self_sf7[163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1640]),
        .S(self_sf7[1640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1641]),
        .S(self_sf7[1641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1642]),
        .S(self_sf7[1642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1643]),
        .S(self_sf7[1643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1644]),
        .S(self_sf7[1644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1645]),
        .S(self_sf7[1645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1646]),
        .S(self_sf7[1646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1647]),
        .S(self_sf7[1647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1648]),
        .S(self_sf7[1648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1649]),
        .S(self_sf7[1649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[164]),
        .S(self_sf7[164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1650]),
        .S(self_sf7[1650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1651]),
        .S(self_sf7[1651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1652]),
        .S(self_sf7[1652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1653]),
        .S(self_sf7[1653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1654]),
        .S(self_sf7[1654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1655]),
        .S(self_sf7[1655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1656]),
        .S(self_sf7[1656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1657]),
        .S(self_sf7[1657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1658]),
        .S(self_sf7[1658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1659]),
        .S(self_sf7[1659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[165]),
        .S(self_sf7[165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1660]),
        .S(self_sf7[1660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1661]),
        .S(self_sf7[1661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1662]),
        .S(self_sf7[1662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1663]),
        .S(self_sf7[1663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1664]),
        .S(self_sf7[1664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1665]),
        .S(self_sf7[1665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1666]),
        .S(self_sf7[1666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1667]),
        .S(self_sf7[1667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1668]),
        .S(self_sf7[1668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1669]),
        .S(self_sf7[1669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[166]),
        .S(self_sf7[166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1670]),
        .S(self_sf7[1670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1671]),
        .S(self_sf7[1671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1672]),
        .S(self_sf7[1672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1673]),
        .S(self_sf7[1673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1674]),
        .S(self_sf7[1674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1675]),
        .S(self_sf7[1675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1676]),
        .S(self_sf7[1676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1677]),
        .S(self_sf7[1677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1678]),
        .S(self_sf7[1678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1679]),
        .S(self_sf7[1679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[167]),
        .S(self_sf7[167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1680]),
        .S(self_sf7[1680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1681]),
        .S(self_sf7[1681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1682]),
        .S(self_sf7[1682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1683]),
        .S(self_sf7[1683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1684]),
        .S(self_sf7[1684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1685]),
        .S(self_sf7[1685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1686]),
        .S(self_sf7[1686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1687]),
        .S(self_sf7[1687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1688]),
        .S(self_sf7[1688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1689]),
        .S(self_sf7[1689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[168]),
        .S(self_sf7[168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1690]),
        .S(self_sf7[1690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1691]),
        .S(self_sf7[1691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1692]),
        .S(self_sf7[1692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1693]),
        .S(self_sf7[1693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1694]),
        .S(self_sf7[1694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1695]),
        .S(self_sf7[1695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1696]),
        .S(self_sf7[1696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1697]),
        .S(self_sf7[1697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1698]),
        .S(self_sf7[1698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1699]),
        .S(self_sf7[1699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[169]),
        .S(self_sf7[169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[16].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[16]),
        .S(self_sf7[16]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1700]),
        .S(self_sf7[1700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1701]),
        .S(self_sf7[1701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1702]),
        .S(self_sf7[1702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1703]),
        .S(self_sf7[1703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1704]),
        .S(self_sf7[1704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1705]),
        .S(self_sf7[1705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1706]),
        .S(self_sf7[1706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1707]),
        .S(self_sf7[1707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1708]),
        .S(self_sf7[1708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1709]),
        .S(self_sf7[1709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[170]),
        .S(self_sf7[170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1710]),
        .S(self_sf7[1710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1711]),
        .S(self_sf7[1711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1712]),
        .S(self_sf7[1712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1713]),
        .S(self_sf7[1713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1714]),
        .S(self_sf7[1714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1715]),
        .S(self_sf7[1715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1716]),
        .S(self_sf7[1716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1717]),
        .S(self_sf7[1717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1718]),
        .S(self_sf7[1718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1719]),
        .S(self_sf7[1719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[171]),
        .S(self_sf7[171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1720]),
        .S(self_sf7[1720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1721]),
        .S(self_sf7[1721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1722]),
        .S(self_sf7[1722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1723]),
        .S(self_sf7[1723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1724]),
        .S(self_sf7[1724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1725]),
        .S(self_sf7[1725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1726]),
        .S(self_sf7[1726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1727]),
        .S(self_sf7[1727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1728]),
        .S(self_sf7[1728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1729]),
        .S(self_sf7[1729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[172]),
        .S(self_sf7[172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1730]),
        .S(self_sf7[1730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1731]),
        .S(self_sf7[1731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1732]),
        .S(self_sf7[1732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1733]),
        .S(self_sf7[1733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1734]),
        .S(self_sf7[1734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1735]),
        .S(self_sf7[1735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1736]),
        .S(self_sf7[1736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1737]),
        .S(self_sf7[1737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1738]),
        .S(self_sf7[1738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1739]),
        .S(self_sf7[1739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[173]),
        .S(self_sf7[173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1740]),
        .S(self_sf7[1740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1741]),
        .S(self_sf7[1741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1742]),
        .S(self_sf7[1742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1743]),
        .S(self_sf7[1743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1744]),
        .S(self_sf7[1744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1745]),
        .S(self_sf7[1745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1746]),
        .S(self_sf7[1746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1747]),
        .S(self_sf7[1747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1748]),
        .S(self_sf7[1748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1749]),
        .S(self_sf7[1749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[174]),
        .S(self_sf7[174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1750]),
        .S(self_sf7[1750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1751]),
        .S(self_sf7[1751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1752]),
        .S(self_sf7[1752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1753]),
        .S(self_sf7[1753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1754]),
        .S(self_sf7[1754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1755]),
        .S(self_sf7[1755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1756]),
        .S(self_sf7[1756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1757]),
        .S(self_sf7[1757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1758]),
        .S(self_sf7[1758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1759]),
        .S(self_sf7[1759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[175]),
        .S(self_sf7[175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1760]),
        .S(self_sf7[1760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1761]),
        .S(self_sf7[1761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1762]),
        .S(self_sf7[1762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1763]),
        .S(self_sf7[1763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1764]),
        .S(self_sf7[1764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1765]),
        .S(self_sf7[1765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1766]),
        .S(self_sf7[1766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1767]),
        .S(self_sf7[1767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1768]),
        .S(self_sf7[1768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1769]),
        .S(self_sf7[1769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[176]),
        .S(self_sf7[176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1770]),
        .S(self_sf7[1770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1771]),
        .S(self_sf7[1771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1772]),
        .S(self_sf7[1772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1773]),
        .S(self_sf7[1773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1774]),
        .S(self_sf7[1774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1775]),
        .S(self_sf7[1775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1776]),
        .S(self_sf7[1776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1777]),
        .S(self_sf7[1777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1778]),
        .S(self_sf7[1778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1779]),
        .S(self_sf7[1779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[177]),
        .S(self_sf7[177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1780]),
        .S(self_sf7[1780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1781]),
        .S(self_sf7[1781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1782]),
        .S(self_sf7[1782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1783]),
        .S(self_sf7[1783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1784]),
        .S(self_sf7[1784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1785]),
        .S(self_sf7[1785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1786]),
        .S(self_sf7[1786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1787]),
        .S(self_sf7[1787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1788]),
        .S(self_sf7[1788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1789]),
        .S(self_sf7[1789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[178]),
        .S(self_sf7[178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1790]),
        .S(self_sf7[1790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1791]),
        .S(self_sf7[1791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1792]),
        .S(self_sf7[1792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1793]),
        .S(self_sf7[1793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1794]),
        .S(self_sf7[1794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1795]),
        .S(self_sf7[1795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1796]),
        .S(self_sf7[1796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1797]),
        .S(self_sf7[1797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1798]),
        .S(self_sf7[1798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1799]),
        .S(self_sf7[1799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[179]),
        .S(self_sf7[179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[17].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[17]),
        .S(self_sf7[17]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[180]),
        .S(self_sf7[180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[181]),
        .S(self_sf7[181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[182]),
        .S(self_sf7[182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[183]),
        .S(self_sf7[183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[184]),
        .S(self_sf7[184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[185]),
        .S(self_sf7[185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[186]),
        .S(self_sf7[186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[187]),
        .S(self_sf7[187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[188]),
        .S(self_sf7[188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[189]),
        .S(self_sf7[189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[18].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[18]),
        .S(self_sf7[18]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[190]),
        .S(self_sf7[190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[191]),
        .S(self_sf7[191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[192]),
        .S(self_sf7[192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[193]),
        .S(self_sf7[193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[194]),
        .S(self_sf7[194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[195]),
        .S(self_sf7[195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[196]),
        .S(self_sf7[196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[197]),
        .S(self_sf7[197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[198]),
        .S(self_sf7[198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[199]),
        .S(self_sf7[199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[19].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[19]),
        .S(self_sf7[19]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1]),
        .S(info_sf7[1]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[200]),
        .S(self_sf7[200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[201]),
        .S(self_sf7[201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[202]),
        .S(self_sf7[202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[203]),
        .S(self_sf7[203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[204]),
        .S(self_sf7[204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[205]),
        .S(self_sf7[205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[206]),
        .S(self_sf7[206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[207]),
        .S(self_sf7[207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[208]),
        .S(self_sf7[208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[209]),
        .S(self_sf7[209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[20].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[20]),
        .S(self_sf7[20]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[210]),
        .S(self_sf7[210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[211]),
        .S(self_sf7[211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[212]),
        .S(self_sf7[212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[213]),
        .S(self_sf7[213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[214]),
        .S(self_sf7[214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[215]),
        .S(self_sf7[215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[216]),
        .S(self_sf7[216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[217]),
        .S(self_sf7[217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[218]),
        .S(self_sf7[218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[219]),
        .S(self_sf7[219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[21].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[21]),
        .S(self_sf7[21]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[220]),
        .S(self_sf7[220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[221]),
        .S(self_sf7[221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[222]),
        .S(self_sf7[222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[223]),
        .S(self_sf7[223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[224]),
        .S(self_sf7[224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[225]),
        .S(self_sf7[225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[226]),
        .S(self_sf7[226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[227]),
        .S(self_sf7[227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[228]),
        .S(self_sf7[228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[229]),
        .S(self_sf7[229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[22].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[22]),
        .S(self_sf7[22]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[230]),
        .S(self_sf7[230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[231]),
        .S(self_sf7[231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[232]),
        .S(self_sf7[232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[233]),
        .S(self_sf7[233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[234]),
        .S(self_sf7[234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[235]),
        .S(self_sf7[235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[236]),
        .S(self_sf7[236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[237]),
        .S(self_sf7[237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[238]),
        .S(self_sf7[238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[239]),
        .S(self_sf7[239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[23].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[23]),
        .S(self_sf7[23]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[240]),
        .S(self_sf7[240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[241]),
        .S(self_sf7[241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[242]),
        .S(self_sf7[242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[243]),
        .S(self_sf7[243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[244]),
        .S(self_sf7[244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[245]),
        .S(self_sf7[245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[246]),
        .S(self_sf7[246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[247]),
        .S(self_sf7[247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[248]),
        .S(self_sf7[248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[249]),
        .S(self_sf7[249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[24].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[24]),
        .S(self_sf7[24]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[250]),
        .S(self_sf7[250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[251]),
        .S(self_sf7[251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[252]),
        .S(self_sf7[252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[253]),
        .S(self_sf7[253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[254]),
        .S(self_sf7[254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[255]),
        .S(self_sf7[255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[256]),
        .S(self_sf7[256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[257]),
        .S(self_sf7[257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[258]),
        .S(self_sf7[258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[259]),
        .S(self_sf7[259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[25].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[25]),
        .S(self_sf7[25]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[260]),
        .S(self_sf7[260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[261]),
        .S(self_sf7[261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[262]),
        .S(self_sf7[262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[263]),
        .S(self_sf7[263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[264]),
        .S(self_sf7[264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[265]),
        .S(self_sf7[265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[266]),
        .S(self_sf7[266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[267]),
        .S(self_sf7[267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[268]),
        .S(self_sf7[268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[269]),
        .S(self_sf7[269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[26].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[26]),
        .S(self_sf7[26]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[270]),
        .S(self_sf7[270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[271]),
        .S(self_sf7[271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[272]),
        .S(self_sf7[272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[273]),
        .S(self_sf7[273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[274]),
        .S(self_sf7[274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[275]),
        .S(self_sf7[275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[276]),
        .S(self_sf7[276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[277]),
        .S(self_sf7[277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[278]),
        .S(self_sf7[278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[279]),
        .S(self_sf7[279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[27].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[27]),
        .S(self_sf7[27]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[280]),
        .S(self_sf7[280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[281]),
        .S(self_sf7[281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[282]),
        .S(self_sf7[282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[283]),
        .S(self_sf7[283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[284]),
        .S(self_sf7[284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[285]),
        .S(self_sf7[285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[286]),
        .S(self_sf7[286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[287]),
        .S(self_sf7[287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[288]),
        .S(self_sf7[288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[289]),
        .S(self_sf7[289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[28].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[28]),
        .S(self_sf7[28]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[290]),
        .S(self_sf7[290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[291]),
        .S(self_sf7[291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[292]),
        .S(self_sf7[292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[293]),
        .S(self_sf7[293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[294]),
        .S(self_sf7[294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[295]),
        .S(self_sf7[295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[296]),
        .S(self_sf7[296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[297]),
        .S(self_sf7[297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[298]),
        .S(self_sf7[298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[299]),
        .S(self_sf7[299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[29].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[29]),
        .S(self_sf7[29]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[2].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[2]),
        .S(info_sf7[2]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[300]),
        .S(self_sf7[300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[301]),
        .S(self_sf7[301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[302]),
        .S(self_sf7[302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[303]),
        .S(self_sf7[303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[304]),
        .S(self_sf7[304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[305]),
        .S(self_sf7[305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[306]),
        .S(self_sf7[306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[307]),
        .S(self_sf7[307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[308]),
        .S(self_sf7[308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[309]),
        .S(self_sf7[309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[30].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[30]),
        .S(self_sf7[30]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[310]),
        .S(self_sf7[310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[311]),
        .S(self_sf7[311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[312]),
        .S(self_sf7[312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[313]),
        .S(self_sf7[313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[314]),
        .S(self_sf7[314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[315]),
        .S(self_sf7[315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[316]),
        .S(self_sf7[316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[317]),
        .S(self_sf7[317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[318]),
        .S(self_sf7[318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[319]),
        .S(self_sf7[319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[31].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[31]),
        .S(self_sf7[31]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[320]),
        .S(self_sf7[320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[321]),
        .S(self_sf7[321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[322]),
        .S(self_sf7[322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[323]),
        .S(self_sf7[323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[324]),
        .S(self_sf7[324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[325]),
        .S(self_sf7[325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[326]),
        .S(self_sf7[326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[327]),
        .S(self_sf7[327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[328]),
        .S(self_sf7[328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[329]),
        .S(self_sf7[329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[32].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[32]),
        .S(self_sf7[32]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[330]),
        .S(self_sf7[330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[331]),
        .S(self_sf7[331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[332]),
        .S(self_sf7[332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[333]),
        .S(self_sf7[333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[334]),
        .S(self_sf7[334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[335]),
        .S(self_sf7[335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[336]),
        .S(self_sf7[336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[337]),
        .S(self_sf7[337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[338]),
        .S(self_sf7[338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[339]),
        .S(self_sf7[339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[33].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[33]),
        .S(self_sf7[33]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[340]),
        .S(self_sf7[340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[341]),
        .S(self_sf7[341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[342]),
        .S(self_sf7[342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[343]),
        .S(self_sf7[343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[344]),
        .S(self_sf7[344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[345]),
        .S(self_sf7[345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[346]),
        .S(self_sf7[346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[347]),
        .S(self_sf7[347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[348]),
        .S(self_sf7[348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[349]),
        .S(self_sf7[349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[34].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[34]),
        .S(self_sf7[34]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[350]),
        .S(self_sf7[350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[351]),
        .S(self_sf7[351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[352]),
        .S(self_sf7[352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[353]),
        .S(self_sf7[353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[354]),
        .S(self_sf7[354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[355]),
        .S(self_sf7[355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[356]),
        .S(self_sf7[356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[357]),
        .S(self_sf7[357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[358]),
        .S(self_sf7[358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[359]),
        .S(self_sf7[359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[35].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[35]),
        .S(self_sf7[35]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[360]),
        .S(self_sf7[360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[361]),
        .S(self_sf7[361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[362]),
        .S(self_sf7[362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[363]),
        .S(self_sf7[363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[364]),
        .S(self_sf7[364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[365]),
        .S(self_sf7[365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[366]),
        .S(self_sf7[366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[367]),
        .S(self_sf7[367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[368]),
        .S(self_sf7[368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[369]),
        .S(self_sf7[369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[36].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[36]),
        .S(self_sf7[36]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[370]),
        .S(self_sf7[370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[371]),
        .S(self_sf7[371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[372]),
        .S(self_sf7[372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[373]),
        .S(self_sf7[373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[374]),
        .S(self_sf7[374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[375]),
        .S(self_sf7[375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[376]),
        .S(self_sf7[376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[377]),
        .S(self_sf7[377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[378]),
        .S(self_sf7[378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[379]),
        .S(self_sf7[379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[37].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[37]),
        .S(self_sf7[37]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[380]),
        .S(self_sf7[380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[381]),
        .S(self_sf7[381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[382]),
        .S(self_sf7[382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[383]),
        .S(self_sf7[383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[384]),
        .S(self_sf7[384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[385]),
        .S(self_sf7[385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[386]),
        .S(self_sf7[386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[387]),
        .S(self_sf7[387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[388]),
        .S(self_sf7[388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[389]),
        .S(self_sf7[389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[38].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[38]),
        .S(self_sf7[38]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[390]),
        .S(self_sf7[390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[391]),
        .S(self_sf7[391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[392]),
        .S(self_sf7[392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[393]),
        .S(self_sf7[393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[394]),
        .S(self_sf7[394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[395]),
        .S(self_sf7[395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[396]),
        .S(self_sf7[396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[397]),
        .S(self_sf7[397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[398]),
        .S(self_sf7[398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[399]),
        .S(self_sf7[399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[39].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[39]),
        .S(self_sf7[39]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[3].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[3]),
        .S(info_sf7[3]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[400]),
        .S(self_sf7[400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[401]),
        .S(self_sf7[401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[402]),
        .S(self_sf7[402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[403]),
        .S(self_sf7[403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[404]),
        .S(self_sf7[404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[405]),
        .S(self_sf7[405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[406]),
        .S(self_sf7[406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[407]),
        .S(self_sf7[407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[408]),
        .S(self_sf7[408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[409]),
        .S(self_sf7[409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[40].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[40]),
        .S(self_sf7[40]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[410]),
        .S(self_sf7[410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[411]),
        .S(self_sf7[411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[412]),
        .S(self_sf7[412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[413]),
        .S(self_sf7[413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[414]),
        .S(self_sf7[414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[415]),
        .S(self_sf7[415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[416]),
        .S(self_sf7[416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[417]),
        .S(self_sf7[417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[418]),
        .S(self_sf7[418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[419]),
        .S(self_sf7[419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[41].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[41]),
        .S(self_sf7[41]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[420]),
        .S(self_sf7[420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[421]),
        .S(self_sf7[421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[422]),
        .S(self_sf7[422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[423]),
        .S(self_sf7[423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[424]),
        .S(self_sf7[424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[425]),
        .S(self_sf7[425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[426]),
        .S(self_sf7[426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[427]),
        .S(self_sf7[427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[428]),
        .S(self_sf7[428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[429]),
        .S(self_sf7[429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[42].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[42]),
        .S(self_sf7[42]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[430]),
        .S(self_sf7[430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[431]),
        .S(self_sf7[431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[432]),
        .S(self_sf7[432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[433]),
        .S(self_sf7[433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[434]),
        .S(self_sf7[434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[435]),
        .S(self_sf7[435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[436]),
        .S(self_sf7[436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[437]),
        .S(self_sf7[437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[438]),
        .S(self_sf7[438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[439]),
        .S(self_sf7[439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[43].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[43]),
        .S(self_sf7[43]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[440]),
        .S(self_sf7[440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[441]),
        .S(self_sf7[441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[442]),
        .S(self_sf7[442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[443]),
        .S(self_sf7[443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[444]),
        .S(self_sf7[444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[445]),
        .S(self_sf7[445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[446]),
        .S(self_sf7[446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[447]),
        .S(self_sf7[447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[448]),
        .S(self_sf7[448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[449]),
        .S(self_sf7[449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[44].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[44]),
        .S(self_sf7[44]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[450]),
        .S(self_sf7[450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[451]),
        .S(self_sf7[451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[452]),
        .S(self_sf7[452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[453]),
        .S(self_sf7[453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[454]),
        .S(self_sf7[454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[455]),
        .S(self_sf7[455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[456]),
        .S(self_sf7[456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[457]),
        .S(self_sf7[457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[458]),
        .S(self_sf7[458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[459]),
        .S(self_sf7[459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[45].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[45]),
        .S(self_sf7[45]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[460]),
        .S(self_sf7[460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[461]),
        .S(self_sf7[461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[462]),
        .S(self_sf7[462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[463]),
        .S(self_sf7[463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[464]),
        .S(self_sf7[464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[465]),
        .S(self_sf7[465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[466]),
        .S(self_sf7[466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[467]),
        .S(self_sf7[467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[468]),
        .S(self_sf7[468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[469]),
        .S(self_sf7[469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[46].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[46]),
        .S(self_sf7[46]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[470]),
        .S(self_sf7[470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[471]),
        .S(self_sf7[471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[472]),
        .S(self_sf7[472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[473]),
        .S(self_sf7[473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[474]),
        .S(self_sf7[474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[475]),
        .S(self_sf7[475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[476]),
        .S(self_sf7[476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[477]),
        .S(self_sf7[477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[478]),
        .S(self_sf7[478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[479]),
        .S(self_sf7[479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[47].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[47]),
        .S(self_sf7[47]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[480]),
        .S(self_sf7[480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[481]),
        .S(self_sf7[481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[482]),
        .S(self_sf7[482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[483]),
        .S(self_sf7[483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[484]),
        .S(self_sf7[484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[485]),
        .S(self_sf7[485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[486]),
        .S(self_sf7[486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[487]),
        .S(self_sf7[487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[488]),
        .S(self_sf7[488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[489]),
        .S(self_sf7[489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[48].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[48]),
        .S(self_sf7[48]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[490]),
        .S(self_sf7[490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[491]),
        .S(self_sf7[491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[492]),
        .S(self_sf7[492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[493]),
        .S(self_sf7[493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[494]),
        .S(self_sf7[494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[495]),
        .S(self_sf7[495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[496]),
        .S(self_sf7[496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[497]),
        .S(self_sf7[497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[498]),
        .S(self_sf7[498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[499]),
        .S(self_sf7[499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[49].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[49]),
        .S(self_sf7[49]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[4].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[4]),
        .S(info_sf7[4]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[500]),
        .S(self_sf7[500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[501]),
        .S(self_sf7[501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[502]),
        .S(self_sf7[502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[503]),
        .S(self_sf7[503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[504]),
        .S(self_sf7[504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[505]),
        .S(self_sf7[505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[506]),
        .S(self_sf7[506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[507]),
        .S(self_sf7[507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[508]),
        .S(self_sf7[508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[509]),
        .S(self_sf7[509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[50].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[50]),
        .S(self_sf7[50]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[510]),
        .S(self_sf7[510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[511]),
        .S(self_sf7[511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[512]),
        .S(self_sf7[512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[513]),
        .S(self_sf7[513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[514]),
        .S(self_sf7[514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[515]),
        .S(self_sf7[515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[516]),
        .S(self_sf7[516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[517]),
        .S(self_sf7[517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[518]),
        .S(self_sf7[518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[519]),
        .S(self_sf7[519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[51].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[51]),
        .S(self_sf7[51]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[520]),
        .S(self_sf7[520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[521]),
        .S(self_sf7[521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[522]),
        .S(self_sf7[522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[523]),
        .S(self_sf7[523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[524]),
        .S(self_sf7[524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[525]),
        .S(self_sf7[525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[526]),
        .S(self_sf7[526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[527]),
        .S(self_sf7[527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[528]),
        .S(self_sf7[528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[529]),
        .S(self_sf7[529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[52].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[52]),
        .S(self_sf7[52]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[530]),
        .S(self_sf7[530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[531]),
        .S(self_sf7[531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[532]),
        .S(self_sf7[532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[533]),
        .S(self_sf7[533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[534]),
        .S(self_sf7[534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[535]),
        .S(self_sf7[535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[536]),
        .S(self_sf7[536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[537]),
        .S(self_sf7[537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[538]),
        .S(self_sf7[538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[539]),
        .S(self_sf7[539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[53].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[53]),
        .S(self_sf7[53]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[540]),
        .S(self_sf7[540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[541]),
        .S(self_sf7[541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[542]),
        .S(self_sf7[542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[543]),
        .S(self_sf7[543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[544]),
        .S(self_sf7[544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[545]),
        .S(self_sf7[545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[546]),
        .S(self_sf7[546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[547]),
        .S(self_sf7[547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[548]),
        .S(self_sf7[548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[549]),
        .S(self_sf7[549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[54].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[54]),
        .S(self_sf7[54]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[550]),
        .S(self_sf7[550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[551]),
        .S(self_sf7[551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[552]),
        .S(self_sf7[552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[553]),
        .S(self_sf7[553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[554]),
        .S(self_sf7[554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[555]),
        .S(self_sf7[555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[556]),
        .S(self_sf7[556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[557]),
        .S(self_sf7[557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[558]),
        .S(self_sf7[558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[559]),
        .S(self_sf7[559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[55].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[55]),
        .S(self_sf7[55]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[560]),
        .S(self_sf7[560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[561]),
        .S(self_sf7[561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[562]),
        .S(self_sf7[562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[563]),
        .S(self_sf7[563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[564]),
        .S(self_sf7[564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[565]),
        .S(self_sf7[565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[566]),
        .S(self_sf7[566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[567]),
        .S(self_sf7[567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[568]),
        .S(self_sf7[568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[569]),
        .S(self_sf7[569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[56].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[56]),
        .S(self_sf7[56]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[570]),
        .S(self_sf7[570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[571]),
        .S(self_sf7[571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[572]),
        .S(self_sf7[572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[573]),
        .S(self_sf7[573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[574]),
        .S(self_sf7[574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[575]),
        .S(self_sf7[575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[576]),
        .S(self_sf7[576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[577]),
        .S(self_sf7[577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[578]),
        .S(self_sf7[578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[579]),
        .S(self_sf7[579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[57].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[57]),
        .S(self_sf7[57]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[580]),
        .S(self_sf7[580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[581]),
        .S(self_sf7[581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[582]),
        .S(self_sf7[582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[583]),
        .S(self_sf7[583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[584]),
        .S(self_sf7[584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[585]),
        .S(self_sf7[585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[586]),
        .S(self_sf7[586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[587]),
        .S(self_sf7[587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[588]),
        .S(self_sf7[588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[589]),
        .S(self_sf7[589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[58].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[58]),
        .S(self_sf7[58]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[590]),
        .S(self_sf7[590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[591]),
        .S(self_sf7[591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[592]),
        .S(self_sf7[592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[593]),
        .S(self_sf7[593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[594]),
        .S(self_sf7[594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[595]),
        .S(self_sf7[595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[596]),
        .S(self_sf7[596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[597]),
        .S(self_sf7[597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[598]),
        .S(self_sf7[598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[599]),
        .S(self_sf7[599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[59].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[59]),
        .S(self_sf7[59]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[5].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[5]),
        .S(info_sf7[5]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[600]),
        .S(self_sf7[600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[601]),
        .S(self_sf7[601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[602]),
        .S(self_sf7[602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[603]),
        .S(self_sf7[603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[604]),
        .S(self_sf7[604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[605]),
        .S(self_sf7[605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[606]),
        .S(self_sf7[606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[607]),
        .S(self_sf7[607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[608]),
        .S(self_sf7[608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[609]),
        .S(self_sf7[609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[60].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[60]),
        .S(self_sf7[60]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[610]),
        .S(self_sf7[610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[611]),
        .S(self_sf7[611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[612]),
        .S(self_sf7[612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[613]),
        .S(self_sf7[613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[614]),
        .S(self_sf7[614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[615]),
        .S(self_sf7[615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[616]),
        .S(self_sf7[616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[617]),
        .S(self_sf7[617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[618]),
        .S(self_sf7[618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[619]),
        .S(self_sf7[619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[61].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[61]),
        .S(self_sf7[61]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[620]),
        .S(self_sf7[620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[621]),
        .S(self_sf7[621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[622]),
        .S(self_sf7[622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[623]),
        .S(self_sf7[623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[624]),
        .S(self_sf7[624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[625]),
        .S(self_sf7[625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[626]),
        .S(self_sf7[626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[627]),
        .S(self_sf7[627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[628]),
        .S(self_sf7[628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[629]),
        .S(self_sf7[629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[62].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[62]),
        .S(self_sf7[62]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[630]),
        .S(self_sf7[630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[631]),
        .S(self_sf7[631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[632]),
        .S(self_sf7[632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[633]),
        .S(self_sf7[633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[634]),
        .S(self_sf7[634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[635]),
        .S(self_sf7[635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[636]),
        .S(self_sf7[636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[637]),
        .S(self_sf7[637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[638]),
        .S(self_sf7[638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[639]),
        .S(self_sf7[639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[63].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[63]),
        .S(self_sf7[63]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[640]),
        .S(self_sf7[640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[641]),
        .S(self_sf7[641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[642]),
        .S(self_sf7[642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[643]),
        .S(self_sf7[643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[644]),
        .S(self_sf7[644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[645]),
        .S(self_sf7[645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[646]),
        .S(self_sf7[646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[647]),
        .S(self_sf7[647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[648]),
        .S(self_sf7[648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[649]),
        .S(self_sf7[649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[64].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[64]),
        .S(self_sf7[64]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[650]),
        .S(self_sf7[650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[651]),
        .S(self_sf7[651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[652]),
        .S(self_sf7[652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[653]),
        .S(self_sf7[653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[654]),
        .S(self_sf7[654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[655]),
        .S(self_sf7[655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[656]),
        .S(self_sf7[656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[657]),
        .S(self_sf7[657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[658]),
        .S(self_sf7[658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[659]),
        .S(self_sf7[659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[65].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[65]),
        .S(self_sf7[65]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[660]),
        .S(self_sf7[660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[661]),
        .S(self_sf7[661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[662]),
        .S(self_sf7[662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[663]),
        .S(self_sf7[663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[664]),
        .S(self_sf7[664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[665]),
        .S(self_sf7[665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[666]),
        .S(self_sf7[666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[667]),
        .S(self_sf7[667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[668]),
        .S(self_sf7[668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[669]),
        .S(self_sf7[669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[66].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[66]),
        .S(self_sf7[66]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[670]),
        .S(self_sf7[670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[671]),
        .S(self_sf7[671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[672]),
        .S(self_sf7[672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[673]),
        .S(self_sf7[673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[674]),
        .S(self_sf7[674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[675]),
        .S(self_sf7[675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[676]),
        .S(self_sf7[676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[677]),
        .S(self_sf7[677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[678]),
        .S(self_sf7[678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[679]),
        .S(self_sf7[679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[67].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[67]),
        .S(self_sf7[67]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[680]),
        .S(self_sf7[680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[681]),
        .S(self_sf7[681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[682]),
        .S(self_sf7[682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[683]),
        .S(self_sf7[683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[684]),
        .S(self_sf7[684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[685]),
        .S(self_sf7[685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[686]),
        .S(self_sf7[686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[687]),
        .S(self_sf7[687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[688]),
        .S(self_sf7[688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[689]),
        .S(self_sf7[689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[68].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[68]),
        .S(self_sf7[68]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[690]),
        .S(self_sf7[690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[691]),
        .S(self_sf7[691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[692]),
        .S(self_sf7[692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[693]),
        .S(self_sf7[693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[694]),
        .S(self_sf7[694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[695]),
        .S(self_sf7[695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[696]),
        .S(self_sf7[696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[697]),
        .S(self_sf7[697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[698]),
        .S(self_sf7[698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[699]),
        .S(self_sf7[699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[69].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[69]),
        .S(self_sf7[69]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[6].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[6]),
        .S(info_sf7[6]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[700]),
        .S(self_sf7[700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[701]),
        .S(self_sf7[701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[702]),
        .S(self_sf7[702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[703]),
        .S(self_sf7[703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[704]),
        .S(self_sf7[704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[705]),
        .S(self_sf7[705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[706]),
        .S(self_sf7[706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[707]),
        .S(self_sf7[707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[708]),
        .S(self_sf7[708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[709]),
        .S(self_sf7[709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[70].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[70]),
        .S(self_sf7[70]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[710]),
        .S(self_sf7[710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[711]),
        .S(self_sf7[711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[712]),
        .S(self_sf7[712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[713]),
        .S(self_sf7[713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[714]),
        .S(self_sf7[714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[715]),
        .S(self_sf7[715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[716]),
        .S(self_sf7[716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[717]),
        .S(self_sf7[717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[718]),
        .S(self_sf7[718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[719]),
        .S(self_sf7[719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[71].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[71]),
        .S(self_sf7[71]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[720]),
        .S(self_sf7[720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[721]),
        .S(self_sf7[721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[722]),
        .S(self_sf7[722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[723]),
        .S(self_sf7[723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[724]),
        .S(self_sf7[724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[725]),
        .S(self_sf7[725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[726]),
        .S(self_sf7[726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[727]),
        .S(self_sf7[727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[728]),
        .S(self_sf7[728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[729]),
        .S(self_sf7[729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[72].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[72]),
        .S(self_sf7[72]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[730]),
        .S(self_sf7[730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[731]),
        .S(self_sf7[731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[732]),
        .S(self_sf7[732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[733]),
        .S(self_sf7[733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[734]),
        .S(self_sf7[734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[735]),
        .S(self_sf7[735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[736]),
        .S(self_sf7[736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[737]),
        .S(self_sf7[737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[738]),
        .S(self_sf7[738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[739]),
        .S(self_sf7[739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[73].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[73]),
        .S(self_sf7[73]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[740]),
        .S(self_sf7[740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[741]),
        .S(self_sf7[741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[742]),
        .S(self_sf7[742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[743]),
        .S(self_sf7[743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[744]),
        .S(self_sf7[744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[745]),
        .S(self_sf7[745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[746]),
        .S(self_sf7[746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[747]),
        .S(self_sf7[747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[748]),
        .S(self_sf7[748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[749]),
        .S(self_sf7[749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[74].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[74]),
        .S(self_sf7[74]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[750]),
        .S(self_sf7[750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[751]),
        .S(self_sf7[751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[752]),
        .S(self_sf7[752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[753]),
        .S(self_sf7[753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[754]),
        .S(self_sf7[754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[755]),
        .S(self_sf7[755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[756]),
        .S(self_sf7[756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[757]),
        .S(self_sf7[757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[758]),
        .S(self_sf7[758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[759]),
        .S(self_sf7[759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[75].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[75]),
        .S(self_sf7[75]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[760]),
        .S(self_sf7[760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[761]),
        .S(self_sf7[761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[762]),
        .S(self_sf7[762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[763]),
        .S(self_sf7[763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[764]),
        .S(self_sf7[764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[765]),
        .S(self_sf7[765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[766]),
        .S(self_sf7[766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[767]),
        .S(self_sf7[767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[768]),
        .S(self_sf7[768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[769]),
        .S(self_sf7[769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[76].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[76]),
        .S(self_sf7[76]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[770]),
        .S(self_sf7[770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[771]),
        .S(self_sf7[771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[772]),
        .S(self_sf7[772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[773]),
        .S(self_sf7[773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[774]),
        .S(self_sf7[774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[775]),
        .S(self_sf7[775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[776]),
        .S(self_sf7[776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[777]),
        .S(self_sf7[777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[778]),
        .S(self_sf7[778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[779]),
        .S(self_sf7[779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[77].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[77]),
        .S(self_sf7[77]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[780]),
        .S(self_sf7[780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[781]),
        .S(self_sf7[781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[782]),
        .S(self_sf7[782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[783]),
        .S(self_sf7[783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[784]),
        .S(self_sf7[784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[785]),
        .S(self_sf7[785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[786]),
        .S(self_sf7[786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[787]),
        .S(self_sf7[787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[788]),
        .S(self_sf7[788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[789]),
        .S(self_sf7[789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[78].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[78]),
        .S(self_sf7[78]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[790]),
        .S(self_sf7[790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[791]),
        .S(self_sf7[791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[792]),
        .S(self_sf7[792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[793]),
        .S(self_sf7[793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[794]),
        .S(self_sf7[794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[795]),
        .S(self_sf7[795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[796]),
        .S(self_sf7[796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[797]),
        .S(self_sf7[797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[798]),
        .S(self_sf7[798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[799]),
        .S(self_sf7[799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[79].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[79]),
        .S(self_sf7[79]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[7].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[7]),
        .S(info_sf7[7]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[800].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[800]),
        .S(self_sf7[800]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[801].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[801]),
        .S(self_sf7[801]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[802].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[802]),
        .S(self_sf7[802]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[803].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[803]),
        .S(self_sf7[803]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[804].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[804]),
        .S(self_sf7[804]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[805].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[805]),
        .S(self_sf7[805]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[806].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[806]),
        .S(self_sf7[806]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[807].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[807]),
        .S(self_sf7[807]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[808].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[808]),
        .S(self_sf7[808]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[809].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[809]),
        .S(self_sf7[809]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[80].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[80]),
        .S(self_sf7[80]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[810].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[810]),
        .S(self_sf7[810]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[811].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[811]),
        .S(self_sf7[811]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[812].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[812]),
        .S(self_sf7[812]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[813].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[813]),
        .S(self_sf7[813]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[814].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[814]),
        .S(self_sf7[814]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[815].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[815]),
        .S(self_sf7[815]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[816].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[816]),
        .S(self_sf7[816]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[817].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[817]),
        .S(self_sf7[817]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[818].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[818]),
        .S(self_sf7[818]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[819].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[819]),
        .S(self_sf7[819]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[81].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[81]),
        .S(self_sf7[81]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[820].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[820]),
        .S(self_sf7[820]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[821].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[821]),
        .S(self_sf7[821]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[822].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[822]),
        .S(self_sf7[822]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[823].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[823]),
        .S(self_sf7[823]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[824].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[824]),
        .S(self_sf7[824]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[825].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[825]),
        .S(self_sf7[825]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[826].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[826]),
        .S(self_sf7[826]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[827].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[827]),
        .S(self_sf7[827]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[828].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[828]),
        .S(self_sf7[828]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[829].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[829]),
        .S(self_sf7[829]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[82].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[82]),
        .S(self_sf7[82]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[830].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[830]),
        .S(self_sf7[830]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[831].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[831]),
        .S(self_sf7[831]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[832].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[832]),
        .S(self_sf7[832]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[833].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[833]),
        .S(self_sf7[833]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[834].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[834]),
        .S(self_sf7[834]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[835].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[835]),
        .S(self_sf7[835]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[836].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[836]),
        .S(self_sf7[836]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[837].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[837]),
        .S(self_sf7[837]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[838].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[838]),
        .S(self_sf7[838]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[839].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[839]),
        .S(self_sf7[839]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[83].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[83]),
        .S(self_sf7[83]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[840].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[840]),
        .S(self_sf7[840]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[841].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[841]),
        .S(self_sf7[841]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[842].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[842]),
        .S(self_sf7[842]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[843].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[843]),
        .S(self_sf7[843]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[844].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[844]),
        .S(self_sf7[844]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[845].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[845]),
        .S(self_sf7[845]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[846].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[846]),
        .S(self_sf7[846]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[847].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[847]),
        .S(self_sf7[847]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[848].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[848]),
        .S(self_sf7[848]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[849].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[849]),
        .S(self_sf7[849]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[84].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[84]),
        .S(self_sf7[84]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[850].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[850]),
        .S(self_sf7[850]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[851].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[851]),
        .S(self_sf7[851]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[852].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[852]),
        .S(self_sf7[852]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[853].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[853]),
        .S(self_sf7[853]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[854].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[854]),
        .S(self_sf7[854]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[855].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[855]),
        .S(self_sf7[855]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[856].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[856]),
        .S(self_sf7[856]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[857].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[857]),
        .S(self_sf7[857]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[858].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[858]),
        .S(self_sf7[858]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[859].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[859]),
        .S(self_sf7[859]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[85].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[85]),
        .S(self_sf7[85]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[860].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[860]),
        .S(self_sf7[860]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[861].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[861]),
        .S(self_sf7[861]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[862].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[862]),
        .S(self_sf7[862]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[863].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[863]),
        .S(self_sf7[863]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[864].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[864]),
        .S(self_sf7[864]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[865].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[865]),
        .S(self_sf7[865]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[866].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[866]),
        .S(self_sf7[866]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[867].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[867]),
        .S(self_sf7[867]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[868].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[868]),
        .S(self_sf7[868]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[869].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[869]),
        .S(self_sf7[869]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[86].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[86]),
        .S(self_sf7[86]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[870].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[870]),
        .S(self_sf7[870]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[871].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[871]),
        .S(self_sf7[871]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[872].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[872]),
        .S(self_sf7[872]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[873].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[873]),
        .S(self_sf7[873]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[874].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[874]),
        .S(self_sf7[874]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[875].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[875]),
        .S(self_sf7[875]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[876].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[876]),
        .S(self_sf7[876]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[877].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[877]),
        .S(self_sf7[877]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[878].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[878]),
        .S(self_sf7[878]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[879].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[879]),
        .S(self_sf7[879]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[87].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[87]),
        .S(self_sf7[87]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[880].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[880]),
        .S(self_sf7[880]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[881].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[881]),
        .S(self_sf7[881]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[882].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[882]),
        .S(self_sf7[882]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[883].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[883]),
        .S(self_sf7[883]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[884].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[884]),
        .S(self_sf7[884]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[885].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[885]),
        .S(self_sf7[885]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[886].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[886]),
        .S(self_sf7[886]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[887].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[887]),
        .S(self_sf7[887]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[888].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[888]),
        .S(self_sf7[888]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[889].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[889]),
        .S(self_sf7[889]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[88].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[88]),
        .S(self_sf7[88]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[890].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[890]),
        .S(self_sf7[890]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[891].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[891]),
        .S(self_sf7[891]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[892].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[892]),
        .S(self_sf7[892]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[893].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[893]),
        .S(self_sf7[893]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[894].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[894]),
        .S(self_sf7[894]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[895].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[895]),
        .S(self_sf7[895]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[896].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[896]),
        .S(self_sf7[896]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[897].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[897]),
        .S(self_sf7[897]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[898].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[898]),
        .S(self_sf7[898]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[899].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[899]),
        .S(self_sf7[899]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[89].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[89]),
        .S(self_sf7[89]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[8].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[8]),
        .S(self_sf7[8]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[900].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[900]),
        .S(self_sf7[900]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[901].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[901]),
        .S(self_sf7[901]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[902].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[902]),
        .S(self_sf7[902]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[903].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[903]),
        .S(self_sf7[903]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[904].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[904]),
        .S(self_sf7[904]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[905].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[905]),
        .S(self_sf7[905]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[906].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[906]),
        .S(self_sf7[906]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[907].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[907]),
        .S(self_sf7[907]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[908].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[908]),
        .S(self_sf7[908]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[909].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[909]),
        .S(self_sf7[909]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[90].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[90]),
        .S(self_sf7[90]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[910].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[910]),
        .S(self_sf7[910]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[911].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[911]),
        .S(self_sf7[911]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[912].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[912]),
        .S(self_sf7[912]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[913].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[913]),
        .S(self_sf7[913]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[914].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[914]),
        .S(self_sf7[914]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[915].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[915]),
        .S(self_sf7[915]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[916].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[916]),
        .S(self_sf7[916]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[917].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[917]),
        .S(self_sf7[917]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[918].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[918]),
        .S(self_sf7[918]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[919].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[919]),
        .S(self_sf7[919]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[91].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[91]),
        .S(self_sf7[91]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[920].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[920]),
        .S(self_sf7[920]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[921].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[921]),
        .S(self_sf7[921]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[922].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[922]),
        .S(self_sf7[922]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[923].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[923]),
        .S(self_sf7[923]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[924].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[924]),
        .S(self_sf7[924]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[925].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[925]),
        .S(self_sf7[925]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[926].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[926]),
        .S(self_sf7[926]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[927].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[927]),
        .S(self_sf7[927]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[928].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[928]),
        .S(self_sf7[928]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[929].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[929]),
        .S(self_sf7[929]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[92].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[92]),
        .S(self_sf7[92]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[930].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[930]),
        .S(self_sf7[930]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[931].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[931]),
        .S(self_sf7[931]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[932].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[932]),
        .S(self_sf7[932]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[933].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[933]),
        .S(self_sf7[933]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[934].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[934]),
        .S(self_sf7[934]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[935].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[935]),
        .S(self_sf7[935]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[936].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[936]),
        .S(self_sf7[936]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[937].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[937]),
        .S(self_sf7[937]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[938].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[938]),
        .S(self_sf7[938]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[939].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[939]),
        .S(self_sf7[939]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[93].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[93]),
        .S(self_sf7[93]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[940].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[940]),
        .S(self_sf7[940]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[941].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[941]),
        .S(self_sf7[941]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[942].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[942]),
        .S(self_sf7[942]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[943].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[943]),
        .S(self_sf7[943]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[944].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[944]),
        .S(self_sf7[944]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[945].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[945]),
        .S(self_sf7[945]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[946].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[946]),
        .S(self_sf7[946]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[947].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[947]),
        .S(self_sf7[947]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[948].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[948]),
        .S(self_sf7[948]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[949].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[949]),
        .S(self_sf7[949]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[94].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[94]),
        .S(self_sf7[94]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[950].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[950]),
        .S(self_sf7[950]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[951].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[951]),
        .S(self_sf7[951]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[952].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[952]),
        .S(self_sf7[952]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[953].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[953]),
        .S(self_sf7[953]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[954].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[954]),
        .S(self_sf7[954]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[955].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[955]),
        .S(self_sf7[955]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[956].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[956]),
        .S(self_sf7[956]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[957].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[957]),
        .S(self_sf7[957]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[958].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[958]),
        .S(self_sf7[958]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[959].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[959]),
        .S(self_sf7[959]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[95].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[95]),
        .S(self_sf7[95]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[960].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[960]),
        .S(self_sf7[960]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[961].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[961]),
        .S(self_sf7[961]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[962].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[962]),
        .S(self_sf7[962]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[963].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[963]),
        .S(self_sf7[963]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[964].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[964]),
        .S(self_sf7[964]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[965].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[965]),
        .S(self_sf7[965]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[966].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[966]),
        .S(self_sf7[966]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[967].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[967]),
        .S(self_sf7[967]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[968].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[968]),
        .S(self_sf7[968]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[969].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[969]),
        .S(self_sf7[969]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[96].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[96]),
        .S(self_sf7[96]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[970].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[970]),
        .S(self_sf7[970]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[971].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[971]),
        .S(self_sf7[971]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[972].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[972]),
        .S(self_sf7[972]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[973].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[973]),
        .S(self_sf7[973]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[974].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[974]),
        .S(self_sf7[974]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[975].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[975]),
        .S(self_sf7[975]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[976].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[976]),
        .S(self_sf7[976]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[977].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[977]),
        .S(self_sf7[977]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[978].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[978]),
        .S(self_sf7[978]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[979].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[979]),
        .S(self_sf7[979]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[97].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[97]),
        .S(self_sf7[97]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[980].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[980]),
        .S(self_sf7[980]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[981].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[981]),
        .S(self_sf7[981]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[982].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[982]),
        .S(self_sf7[982]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[983].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[983]),
        .S(self_sf7[983]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[984].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[984]),
        .S(self_sf7[984]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[985].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[985]),
        .S(self_sf7[985]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[986].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[986]),
        .S(self_sf7[986]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[987].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[987]),
        .S(self_sf7[987]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[988].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[988]),
        .S(self_sf7[988]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[989].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[989]),
        .S(self_sf7[989]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[98].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[98]),
        .S(self_sf7[98]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[990].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[990]),
        .S(self_sf7[990]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[991].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[991]),
        .S(self_sf7[991]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[992].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[992]),
        .S(self_sf7[992]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[993].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[993]),
        .S(self_sf7[993]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[994].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[994]),
        .S(self_sf7[994]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[995].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[995]),
        .S(self_sf7[995]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[996].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[996]),
        .S(self_sf7[996]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[997].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[997]),
        .S(self_sf7[997]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[998].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[998]),
        .S(self_sf7[998]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[999].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[999]),
        .S(self_sf7[999]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[99].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[99]),
        .S(self_sf7[99]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[9].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[9]),
        .S(self_sf7[9]));
  (* BOX_TYPE = "black_box" *) 
  MUXF8 \activity_ROsf8[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf8[0]),
        .S(self_sf8[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF9 \activity_ROsf9[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf9[0]),
        .S(self_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_0
       (.I0(1'b0),
        .O(self_sf7[1802]));
  LUT1 #(
    .INIT(2'h2)) 
    i_1
       (.I0(1'b0),
        .O(self_sf7[1801]));
  LUT1 #(
    .INIT(2'h2)) 
    i_10
       (.I0(1'b0),
        .O(info_sf8[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_11
       (.I0(1'b0),
        .O(info_sf8[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_12
       (.I0(1'b0),
        .O(info_sf8[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_13
       (.I0(1'b0),
        .O(info_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_14
       (.I0(1'b0),
        .O(info_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_15
       (.I0(1'b0),
        .O(info_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_16
       (.I0(1'b0),
        .O(info_sf8[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_17
       (.I0(1'b0),
        .O(info_sf9[7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_18
       (.I0(1'b0),
        .O(info_sf9[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_19
       (.I0(1'b0),
        .O(info_sf9[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_2
       (.I0(1'b0),
        .O(self_sf7[1800]));
  LUT1 #(
    .INIT(2'h2)) 
    i_20
       (.I0(1'b0),
        .O(info_sf9[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_21
       (.I0(1'b0),
        .O(info_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_22
       (.I0(1'b0),
        .O(info_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_23
       (.I0(1'b0),
        .O(info_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_24
       (.I0(1'b0),
        .O(info_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_3
       (.I0(1'b0),
        .O(self_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_4
       (.I0(1'b0),
        .O(self_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_5
       (.I0(1'b0),
        .O(self_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_6
       (.I0(1'b0),
        .O(self_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_7
       (.I0(1'b0),
        .O(self_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_8
       (.I0(1'b0),
        .O(self_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_9
       (.I0(1'b0),
        .O(info_sf8[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst
       (.I0(self_sf7[7]),
        .O(info_sf7[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__0
       (.I0(self_sf7[6]),
        .O(info_sf7[6]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__1
       (.I0(self_sf7[5]),
        .O(info_sf7[5]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__2
       (.I0(self_sf7[4]),
        .O(info_sf7[4]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__3
       (.I0(self_sf7[3]),
        .O(info_sf7[3]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__4
       (.I0(self_sf7[2]),
        .O(info_sf7[2]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__5
       (.I0(self_sf7[1]),
        .O(info_sf7[1]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__6
       (.I0(self_sf7[0]),
        .O(info_sf7[0]));
endmodule

(* ORIG_REF_NAME = "muxer" *) (* box_type = "black_box" *) (* dont_touch = "true" *) 
module switch_elements_muxer__3
   (enable_i,
    info_o);
  input enable_i;
  output info_o;

  wire enable_i;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf7;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf8;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf9;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [1802:0]self_sf7;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf8;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf9;

  assign info_o = info_sf7[1];
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[0]),
        .S(info_sf7[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1000].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1000]),
        .S(self_sf7[1000]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1001].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1001]),
        .S(self_sf7[1001]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1002].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1002]),
        .S(self_sf7[1002]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1003].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1003]),
        .S(self_sf7[1003]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1004].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1004]),
        .S(self_sf7[1004]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1005].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1005]),
        .S(self_sf7[1005]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1006].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1006]),
        .S(self_sf7[1006]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1007].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1007]),
        .S(self_sf7[1007]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1008].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1008]),
        .S(self_sf7[1008]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1009].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1009]),
        .S(self_sf7[1009]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[100]),
        .S(self_sf7[100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1010].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1010]),
        .S(self_sf7[1010]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1011].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1011]),
        .S(self_sf7[1011]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1012].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1012]),
        .S(self_sf7[1012]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1013].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1013]),
        .S(self_sf7[1013]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1014].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1014]),
        .S(self_sf7[1014]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1015].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1015]),
        .S(self_sf7[1015]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1016].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1016]),
        .S(self_sf7[1016]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1017].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1017]),
        .S(self_sf7[1017]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1018].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1018]),
        .S(self_sf7[1018]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1019].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1019]),
        .S(self_sf7[1019]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[101]),
        .S(self_sf7[101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1020].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1020]),
        .S(self_sf7[1020]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1021].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1021]),
        .S(self_sf7[1021]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1022].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1022]),
        .S(self_sf7[1022]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1023].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1023]),
        .S(self_sf7[1023]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1024].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1024]),
        .S(self_sf7[1024]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1025].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1025]),
        .S(self_sf7[1025]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1026].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1026]),
        .S(self_sf7[1026]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1027].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1027]),
        .S(self_sf7[1027]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1028].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1028]),
        .S(self_sf7[1028]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1029].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1029]),
        .S(self_sf7[1029]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[102]),
        .S(self_sf7[102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1030].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1030]),
        .S(self_sf7[1030]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1031].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1031]),
        .S(self_sf7[1031]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1032].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1032]),
        .S(self_sf7[1032]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1033].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1033]),
        .S(self_sf7[1033]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1034].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1034]),
        .S(self_sf7[1034]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1035].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1035]),
        .S(self_sf7[1035]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1036].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1036]),
        .S(self_sf7[1036]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1037].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1037]),
        .S(self_sf7[1037]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1038].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1038]),
        .S(self_sf7[1038]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1039].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1039]),
        .S(self_sf7[1039]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[103]),
        .S(self_sf7[103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1040].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1040]),
        .S(self_sf7[1040]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1041].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1041]),
        .S(self_sf7[1041]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1042].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1042]),
        .S(self_sf7[1042]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1043].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1043]),
        .S(self_sf7[1043]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1044].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1044]),
        .S(self_sf7[1044]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1045].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1045]),
        .S(self_sf7[1045]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1046].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1046]),
        .S(self_sf7[1046]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1047].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1047]),
        .S(self_sf7[1047]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1048].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1048]),
        .S(self_sf7[1048]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1049].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1049]),
        .S(self_sf7[1049]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[104]),
        .S(self_sf7[104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1050].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1050]),
        .S(self_sf7[1050]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1051].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1051]),
        .S(self_sf7[1051]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1052].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1052]),
        .S(self_sf7[1052]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1053].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1053]),
        .S(self_sf7[1053]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1054].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1054]),
        .S(self_sf7[1054]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1055].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1055]),
        .S(self_sf7[1055]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1056].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1056]),
        .S(self_sf7[1056]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1057].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1057]),
        .S(self_sf7[1057]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1058].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1058]),
        .S(self_sf7[1058]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1059].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1059]),
        .S(self_sf7[1059]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[105]),
        .S(self_sf7[105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1060].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1060]),
        .S(self_sf7[1060]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1061].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1061]),
        .S(self_sf7[1061]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1062].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1062]),
        .S(self_sf7[1062]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1063].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1063]),
        .S(self_sf7[1063]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1064].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1064]),
        .S(self_sf7[1064]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1065].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1065]),
        .S(self_sf7[1065]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1066].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1066]),
        .S(self_sf7[1066]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1067].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1067]),
        .S(self_sf7[1067]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1068].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1068]),
        .S(self_sf7[1068]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1069].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1069]),
        .S(self_sf7[1069]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[106]),
        .S(self_sf7[106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1070].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1070]),
        .S(self_sf7[1070]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1071].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1071]),
        .S(self_sf7[1071]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1072].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1072]),
        .S(self_sf7[1072]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1073].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1073]),
        .S(self_sf7[1073]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1074].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1074]),
        .S(self_sf7[1074]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1075].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1075]),
        .S(self_sf7[1075]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1076].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1076]),
        .S(self_sf7[1076]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1077].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1077]),
        .S(self_sf7[1077]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1078].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1078]),
        .S(self_sf7[1078]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1079].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1079]),
        .S(self_sf7[1079]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[107]),
        .S(self_sf7[107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1080].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1080]),
        .S(self_sf7[1080]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1081].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1081]),
        .S(self_sf7[1081]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1082].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1082]),
        .S(self_sf7[1082]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1083].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1083]),
        .S(self_sf7[1083]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1084].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1084]),
        .S(self_sf7[1084]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1085].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1085]),
        .S(self_sf7[1085]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1086].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1086]),
        .S(self_sf7[1086]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1087].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1087]),
        .S(self_sf7[1087]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1088].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1088]),
        .S(self_sf7[1088]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1089].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1089]),
        .S(self_sf7[1089]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[108]),
        .S(self_sf7[108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1090].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1090]),
        .S(self_sf7[1090]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1091].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1091]),
        .S(self_sf7[1091]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1092].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1092]),
        .S(self_sf7[1092]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1093].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1093]),
        .S(self_sf7[1093]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1094].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1094]),
        .S(self_sf7[1094]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1095].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1095]),
        .S(self_sf7[1095]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1096].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1096]),
        .S(self_sf7[1096]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1097].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1097]),
        .S(self_sf7[1097]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1098].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1098]),
        .S(self_sf7[1098]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1099].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1099]),
        .S(self_sf7[1099]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[109]),
        .S(self_sf7[109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[10].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[10]),
        .S(self_sf7[10]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1100]),
        .S(self_sf7[1100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1101]),
        .S(self_sf7[1101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1102]),
        .S(self_sf7[1102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1103]),
        .S(self_sf7[1103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1104]),
        .S(self_sf7[1104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1105]),
        .S(self_sf7[1105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1106]),
        .S(self_sf7[1106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1107]),
        .S(self_sf7[1107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1108]),
        .S(self_sf7[1108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1109]),
        .S(self_sf7[1109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[110]),
        .S(self_sf7[110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1110]),
        .S(self_sf7[1110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1111]),
        .S(self_sf7[1111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1112]),
        .S(self_sf7[1112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1113]),
        .S(self_sf7[1113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1114]),
        .S(self_sf7[1114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1115]),
        .S(self_sf7[1115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1116]),
        .S(self_sf7[1116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1117]),
        .S(self_sf7[1117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1118]),
        .S(self_sf7[1118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1119]),
        .S(self_sf7[1119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[111]),
        .S(self_sf7[111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1120]),
        .S(self_sf7[1120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1121]),
        .S(self_sf7[1121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1122]),
        .S(self_sf7[1122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1123]),
        .S(self_sf7[1123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1124]),
        .S(self_sf7[1124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1125]),
        .S(self_sf7[1125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1126]),
        .S(self_sf7[1126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1127]),
        .S(self_sf7[1127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1128]),
        .S(self_sf7[1128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1129]),
        .S(self_sf7[1129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[112]),
        .S(self_sf7[112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1130]),
        .S(self_sf7[1130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1131]),
        .S(self_sf7[1131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1132]),
        .S(self_sf7[1132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1133]),
        .S(self_sf7[1133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1134]),
        .S(self_sf7[1134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1135]),
        .S(self_sf7[1135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1136]),
        .S(self_sf7[1136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1137]),
        .S(self_sf7[1137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1138]),
        .S(self_sf7[1138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1139]),
        .S(self_sf7[1139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[113]),
        .S(self_sf7[113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1140]),
        .S(self_sf7[1140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1141]),
        .S(self_sf7[1141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1142]),
        .S(self_sf7[1142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1143]),
        .S(self_sf7[1143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1144]),
        .S(self_sf7[1144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1145]),
        .S(self_sf7[1145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1146]),
        .S(self_sf7[1146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1147]),
        .S(self_sf7[1147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1148]),
        .S(self_sf7[1148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1149]),
        .S(self_sf7[1149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[114]),
        .S(self_sf7[114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1150]),
        .S(self_sf7[1150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1151]),
        .S(self_sf7[1151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1152]),
        .S(self_sf7[1152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1153]),
        .S(self_sf7[1153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1154]),
        .S(self_sf7[1154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1155]),
        .S(self_sf7[1155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1156]),
        .S(self_sf7[1156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1157]),
        .S(self_sf7[1157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1158]),
        .S(self_sf7[1158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1159]),
        .S(self_sf7[1159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[115]),
        .S(self_sf7[115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1160]),
        .S(self_sf7[1160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1161]),
        .S(self_sf7[1161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1162]),
        .S(self_sf7[1162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1163]),
        .S(self_sf7[1163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1164]),
        .S(self_sf7[1164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1165]),
        .S(self_sf7[1165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1166]),
        .S(self_sf7[1166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1167]),
        .S(self_sf7[1167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1168]),
        .S(self_sf7[1168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1169]),
        .S(self_sf7[1169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[116]),
        .S(self_sf7[116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1170]),
        .S(self_sf7[1170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1171]),
        .S(self_sf7[1171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1172]),
        .S(self_sf7[1172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1173]),
        .S(self_sf7[1173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1174]),
        .S(self_sf7[1174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1175]),
        .S(self_sf7[1175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1176]),
        .S(self_sf7[1176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1177]),
        .S(self_sf7[1177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1178]),
        .S(self_sf7[1178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1179]),
        .S(self_sf7[1179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[117]),
        .S(self_sf7[117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1180]),
        .S(self_sf7[1180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1181]),
        .S(self_sf7[1181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1182]),
        .S(self_sf7[1182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1183]),
        .S(self_sf7[1183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1184]),
        .S(self_sf7[1184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1185]),
        .S(self_sf7[1185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1186]),
        .S(self_sf7[1186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1187]),
        .S(self_sf7[1187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1188]),
        .S(self_sf7[1188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1189]),
        .S(self_sf7[1189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[118]),
        .S(self_sf7[118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1190]),
        .S(self_sf7[1190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1191]),
        .S(self_sf7[1191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1192]),
        .S(self_sf7[1192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1193]),
        .S(self_sf7[1193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1194]),
        .S(self_sf7[1194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1195]),
        .S(self_sf7[1195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1196]),
        .S(self_sf7[1196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1197]),
        .S(self_sf7[1197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1198]),
        .S(self_sf7[1198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1199]),
        .S(self_sf7[1199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[119]),
        .S(self_sf7[119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[11].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[11]),
        .S(self_sf7[11]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1200]),
        .S(self_sf7[1200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1201]),
        .S(self_sf7[1201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1202]),
        .S(self_sf7[1202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1203]),
        .S(self_sf7[1203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1204]),
        .S(self_sf7[1204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1205]),
        .S(self_sf7[1205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1206]),
        .S(self_sf7[1206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1207]),
        .S(self_sf7[1207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1208]),
        .S(self_sf7[1208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1209]),
        .S(self_sf7[1209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[120]),
        .S(self_sf7[120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1210]),
        .S(self_sf7[1210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1211]),
        .S(self_sf7[1211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1212]),
        .S(self_sf7[1212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1213]),
        .S(self_sf7[1213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1214]),
        .S(self_sf7[1214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1215]),
        .S(self_sf7[1215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1216]),
        .S(self_sf7[1216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1217]),
        .S(self_sf7[1217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1218]),
        .S(self_sf7[1218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1219]),
        .S(self_sf7[1219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[121]),
        .S(self_sf7[121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1220]),
        .S(self_sf7[1220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1221]),
        .S(self_sf7[1221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1222]),
        .S(self_sf7[1222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1223]),
        .S(self_sf7[1223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1224]),
        .S(self_sf7[1224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1225]),
        .S(self_sf7[1225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1226]),
        .S(self_sf7[1226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1227]),
        .S(self_sf7[1227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1228]),
        .S(self_sf7[1228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1229]),
        .S(self_sf7[1229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[122]),
        .S(self_sf7[122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1230]),
        .S(self_sf7[1230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1231]),
        .S(self_sf7[1231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1232]),
        .S(self_sf7[1232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1233]),
        .S(self_sf7[1233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1234]),
        .S(self_sf7[1234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1235]),
        .S(self_sf7[1235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1236]),
        .S(self_sf7[1236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1237]),
        .S(self_sf7[1237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1238]),
        .S(self_sf7[1238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1239]),
        .S(self_sf7[1239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[123]),
        .S(self_sf7[123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1240]),
        .S(self_sf7[1240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1241]),
        .S(self_sf7[1241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1242]),
        .S(self_sf7[1242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1243]),
        .S(self_sf7[1243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1244]),
        .S(self_sf7[1244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1245]),
        .S(self_sf7[1245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1246]),
        .S(self_sf7[1246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1247]),
        .S(self_sf7[1247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1248]),
        .S(self_sf7[1248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1249]),
        .S(self_sf7[1249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[124]),
        .S(self_sf7[124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1250]),
        .S(self_sf7[1250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1251]),
        .S(self_sf7[1251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1252]),
        .S(self_sf7[1252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1253]),
        .S(self_sf7[1253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1254]),
        .S(self_sf7[1254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1255]),
        .S(self_sf7[1255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1256]),
        .S(self_sf7[1256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1257]),
        .S(self_sf7[1257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1258]),
        .S(self_sf7[1258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1259]),
        .S(self_sf7[1259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[125]),
        .S(self_sf7[125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1260]),
        .S(self_sf7[1260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1261]),
        .S(self_sf7[1261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1262]),
        .S(self_sf7[1262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1263]),
        .S(self_sf7[1263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1264]),
        .S(self_sf7[1264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1265]),
        .S(self_sf7[1265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1266]),
        .S(self_sf7[1266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1267]),
        .S(self_sf7[1267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1268]),
        .S(self_sf7[1268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1269]),
        .S(self_sf7[1269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[126]),
        .S(self_sf7[126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1270]),
        .S(self_sf7[1270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1271]),
        .S(self_sf7[1271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1272]),
        .S(self_sf7[1272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1273]),
        .S(self_sf7[1273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1274]),
        .S(self_sf7[1274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1275]),
        .S(self_sf7[1275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1276]),
        .S(self_sf7[1276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1277]),
        .S(self_sf7[1277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1278]),
        .S(self_sf7[1278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1279]),
        .S(self_sf7[1279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[127]),
        .S(self_sf7[127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1280]),
        .S(self_sf7[1280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1281]),
        .S(self_sf7[1281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1282]),
        .S(self_sf7[1282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1283]),
        .S(self_sf7[1283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1284]),
        .S(self_sf7[1284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1285]),
        .S(self_sf7[1285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1286]),
        .S(self_sf7[1286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1287]),
        .S(self_sf7[1287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1288]),
        .S(self_sf7[1288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1289]),
        .S(self_sf7[1289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[128]),
        .S(self_sf7[128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1290]),
        .S(self_sf7[1290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1291]),
        .S(self_sf7[1291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1292]),
        .S(self_sf7[1292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1293]),
        .S(self_sf7[1293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1294]),
        .S(self_sf7[1294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1295]),
        .S(self_sf7[1295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1296]),
        .S(self_sf7[1296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1297]),
        .S(self_sf7[1297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1298]),
        .S(self_sf7[1298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1299]),
        .S(self_sf7[1299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[129]),
        .S(self_sf7[129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[12].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[12]),
        .S(self_sf7[12]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1300]),
        .S(self_sf7[1300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1301]),
        .S(self_sf7[1301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1302]),
        .S(self_sf7[1302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1303]),
        .S(self_sf7[1303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1304]),
        .S(self_sf7[1304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1305]),
        .S(self_sf7[1305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1306]),
        .S(self_sf7[1306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1307]),
        .S(self_sf7[1307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1308]),
        .S(self_sf7[1308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1309]),
        .S(self_sf7[1309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[130]),
        .S(self_sf7[130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1310]),
        .S(self_sf7[1310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1311]),
        .S(self_sf7[1311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1312]),
        .S(self_sf7[1312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1313]),
        .S(self_sf7[1313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1314]),
        .S(self_sf7[1314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1315]),
        .S(self_sf7[1315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1316]),
        .S(self_sf7[1316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1317]),
        .S(self_sf7[1317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1318]),
        .S(self_sf7[1318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1319]),
        .S(self_sf7[1319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[131]),
        .S(self_sf7[131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1320]),
        .S(self_sf7[1320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1321]),
        .S(self_sf7[1321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1322]),
        .S(self_sf7[1322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1323]),
        .S(self_sf7[1323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1324]),
        .S(self_sf7[1324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1325]),
        .S(self_sf7[1325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1326]),
        .S(self_sf7[1326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1327]),
        .S(self_sf7[1327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1328]),
        .S(self_sf7[1328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1329]),
        .S(self_sf7[1329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[132]),
        .S(self_sf7[132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1330]),
        .S(self_sf7[1330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1331]),
        .S(self_sf7[1331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1332]),
        .S(self_sf7[1332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1333]),
        .S(self_sf7[1333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1334]),
        .S(self_sf7[1334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1335]),
        .S(self_sf7[1335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1336]),
        .S(self_sf7[1336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1337]),
        .S(self_sf7[1337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1338]),
        .S(self_sf7[1338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1339]),
        .S(self_sf7[1339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[133]),
        .S(self_sf7[133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1340]),
        .S(self_sf7[1340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1341]),
        .S(self_sf7[1341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1342]),
        .S(self_sf7[1342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1343]),
        .S(self_sf7[1343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1344]),
        .S(self_sf7[1344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1345]),
        .S(self_sf7[1345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1346]),
        .S(self_sf7[1346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1347]),
        .S(self_sf7[1347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1348]),
        .S(self_sf7[1348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1349]),
        .S(self_sf7[1349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[134]),
        .S(self_sf7[134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1350]),
        .S(self_sf7[1350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1351]),
        .S(self_sf7[1351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1352]),
        .S(self_sf7[1352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1353]),
        .S(self_sf7[1353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1354]),
        .S(self_sf7[1354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1355]),
        .S(self_sf7[1355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1356]),
        .S(self_sf7[1356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1357]),
        .S(self_sf7[1357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1358]),
        .S(self_sf7[1358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1359]),
        .S(self_sf7[1359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[135]),
        .S(self_sf7[135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1360]),
        .S(self_sf7[1360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1361]),
        .S(self_sf7[1361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1362]),
        .S(self_sf7[1362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1363]),
        .S(self_sf7[1363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1364]),
        .S(self_sf7[1364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1365]),
        .S(self_sf7[1365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1366]),
        .S(self_sf7[1366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1367]),
        .S(self_sf7[1367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1368]),
        .S(self_sf7[1368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1369]),
        .S(self_sf7[1369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[136]),
        .S(self_sf7[136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1370]),
        .S(self_sf7[1370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1371]),
        .S(self_sf7[1371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1372]),
        .S(self_sf7[1372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1373]),
        .S(self_sf7[1373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1374]),
        .S(self_sf7[1374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1375]),
        .S(self_sf7[1375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1376]),
        .S(self_sf7[1376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1377]),
        .S(self_sf7[1377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1378]),
        .S(self_sf7[1378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1379]),
        .S(self_sf7[1379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[137]),
        .S(self_sf7[137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1380]),
        .S(self_sf7[1380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1381]),
        .S(self_sf7[1381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1382]),
        .S(self_sf7[1382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1383]),
        .S(self_sf7[1383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1384]),
        .S(self_sf7[1384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1385]),
        .S(self_sf7[1385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1386]),
        .S(self_sf7[1386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1387]),
        .S(self_sf7[1387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1388]),
        .S(self_sf7[1388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1389]),
        .S(self_sf7[1389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[138]),
        .S(self_sf7[138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1390]),
        .S(self_sf7[1390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1391]),
        .S(self_sf7[1391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1392]),
        .S(self_sf7[1392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1393]),
        .S(self_sf7[1393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1394]),
        .S(self_sf7[1394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1395]),
        .S(self_sf7[1395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1396]),
        .S(self_sf7[1396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1397]),
        .S(self_sf7[1397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1398]),
        .S(self_sf7[1398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1399]),
        .S(self_sf7[1399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[139]),
        .S(self_sf7[139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[13].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[13]),
        .S(self_sf7[13]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1400]),
        .S(self_sf7[1400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1401]),
        .S(self_sf7[1401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1402]),
        .S(self_sf7[1402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1403]),
        .S(self_sf7[1403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1404]),
        .S(self_sf7[1404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1405]),
        .S(self_sf7[1405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1406]),
        .S(self_sf7[1406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1407]),
        .S(self_sf7[1407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1408]),
        .S(self_sf7[1408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1409]),
        .S(self_sf7[1409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[140]),
        .S(self_sf7[140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1410]),
        .S(self_sf7[1410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1411]),
        .S(self_sf7[1411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1412]),
        .S(self_sf7[1412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1413]),
        .S(self_sf7[1413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1414]),
        .S(self_sf7[1414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1415]),
        .S(self_sf7[1415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1416]),
        .S(self_sf7[1416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1417]),
        .S(self_sf7[1417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1418]),
        .S(self_sf7[1418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1419]),
        .S(self_sf7[1419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[141]),
        .S(self_sf7[141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1420]),
        .S(self_sf7[1420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1421]),
        .S(self_sf7[1421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1422]),
        .S(self_sf7[1422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1423]),
        .S(self_sf7[1423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1424]),
        .S(self_sf7[1424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1425]),
        .S(self_sf7[1425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1426]),
        .S(self_sf7[1426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1427]),
        .S(self_sf7[1427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1428]),
        .S(self_sf7[1428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1429]),
        .S(self_sf7[1429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[142]),
        .S(self_sf7[142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1430]),
        .S(self_sf7[1430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1431]),
        .S(self_sf7[1431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1432]),
        .S(self_sf7[1432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1433]),
        .S(self_sf7[1433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1434]),
        .S(self_sf7[1434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1435]),
        .S(self_sf7[1435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1436]),
        .S(self_sf7[1436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1437]),
        .S(self_sf7[1437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1438]),
        .S(self_sf7[1438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1439]),
        .S(self_sf7[1439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[143]),
        .S(self_sf7[143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1440]),
        .S(self_sf7[1440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1441]),
        .S(self_sf7[1441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1442]),
        .S(self_sf7[1442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1443]),
        .S(self_sf7[1443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1444]),
        .S(self_sf7[1444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1445]),
        .S(self_sf7[1445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1446]),
        .S(self_sf7[1446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1447]),
        .S(self_sf7[1447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1448]),
        .S(self_sf7[1448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1449]),
        .S(self_sf7[1449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[144]),
        .S(self_sf7[144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1450]),
        .S(self_sf7[1450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1451]),
        .S(self_sf7[1451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1452]),
        .S(self_sf7[1452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1453]),
        .S(self_sf7[1453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1454]),
        .S(self_sf7[1454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1455]),
        .S(self_sf7[1455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1456]),
        .S(self_sf7[1456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1457]),
        .S(self_sf7[1457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1458]),
        .S(self_sf7[1458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1459]),
        .S(self_sf7[1459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[145]),
        .S(self_sf7[145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1460]),
        .S(self_sf7[1460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1461]),
        .S(self_sf7[1461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1462]),
        .S(self_sf7[1462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1463]),
        .S(self_sf7[1463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1464]),
        .S(self_sf7[1464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1465]),
        .S(self_sf7[1465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1466]),
        .S(self_sf7[1466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1467]),
        .S(self_sf7[1467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1468]),
        .S(self_sf7[1468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1469]),
        .S(self_sf7[1469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[146]),
        .S(self_sf7[146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1470]),
        .S(self_sf7[1470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1471]),
        .S(self_sf7[1471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1472]),
        .S(self_sf7[1472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1473]),
        .S(self_sf7[1473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1474]),
        .S(self_sf7[1474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1475]),
        .S(self_sf7[1475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1476]),
        .S(self_sf7[1476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1477]),
        .S(self_sf7[1477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1478]),
        .S(self_sf7[1478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1479]),
        .S(self_sf7[1479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[147]),
        .S(self_sf7[147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1480]),
        .S(self_sf7[1480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1481]),
        .S(self_sf7[1481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1482]),
        .S(self_sf7[1482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1483]),
        .S(self_sf7[1483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1484]),
        .S(self_sf7[1484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1485]),
        .S(self_sf7[1485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1486]),
        .S(self_sf7[1486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1487]),
        .S(self_sf7[1487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1488]),
        .S(self_sf7[1488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1489]),
        .S(self_sf7[1489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[148]),
        .S(self_sf7[148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1490]),
        .S(self_sf7[1490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1491]),
        .S(self_sf7[1491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1492]),
        .S(self_sf7[1492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1493]),
        .S(self_sf7[1493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1494]),
        .S(self_sf7[1494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1495]),
        .S(self_sf7[1495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1496]),
        .S(self_sf7[1496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1497]),
        .S(self_sf7[1497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1498]),
        .S(self_sf7[1498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1499]),
        .S(self_sf7[1499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[149]),
        .S(self_sf7[149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[14].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[14]),
        .S(self_sf7[14]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1500]),
        .S(self_sf7[1500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1501]),
        .S(self_sf7[1501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1502]),
        .S(self_sf7[1502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1503]),
        .S(self_sf7[1503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1504]),
        .S(self_sf7[1504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1505]),
        .S(self_sf7[1505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1506]),
        .S(self_sf7[1506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1507]),
        .S(self_sf7[1507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1508]),
        .S(self_sf7[1508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1509]),
        .S(self_sf7[1509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[150]),
        .S(self_sf7[150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1510]),
        .S(self_sf7[1510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1511]),
        .S(self_sf7[1511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1512]),
        .S(self_sf7[1512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1513]),
        .S(self_sf7[1513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1514]),
        .S(self_sf7[1514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1515]),
        .S(self_sf7[1515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1516]),
        .S(self_sf7[1516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1517]),
        .S(self_sf7[1517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1518]),
        .S(self_sf7[1518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1519]),
        .S(self_sf7[1519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[151]),
        .S(self_sf7[151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1520]),
        .S(self_sf7[1520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1521]),
        .S(self_sf7[1521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1522]),
        .S(self_sf7[1522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1523]),
        .S(self_sf7[1523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1524]),
        .S(self_sf7[1524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1525]),
        .S(self_sf7[1525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1526]),
        .S(self_sf7[1526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1527]),
        .S(self_sf7[1527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1528]),
        .S(self_sf7[1528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1529]),
        .S(self_sf7[1529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[152]),
        .S(self_sf7[152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1530]),
        .S(self_sf7[1530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1531]),
        .S(self_sf7[1531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1532]),
        .S(self_sf7[1532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1533]),
        .S(self_sf7[1533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1534]),
        .S(self_sf7[1534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1535]),
        .S(self_sf7[1535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1536]),
        .S(self_sf7[1536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1537]),
        .S(self_sf7[1537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1538]),
        .S(self_sf7[1538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1539]),
        .S(self_sf7[1539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[153]),
        .S(self_sf7[153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1540]),
        .S(self_sf7[1540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1541]),
        .S(self_sf7[1541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1542]),
        .S(self_sf7[1542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1543]),
        .S(self_sf7[1543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1544]),
        .S(self_sf7[1544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1545]),
        .S(self_sf7[1545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1546]),
        .S(self_sf7[1546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1547]),
        .S(self_sf7[1547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1548]),
        .S(self_sf7[1548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1549]),
        .S(self_sf7[1549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[154]),
        .S(self_sf7[154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1550]),
        .S(self_sf7[1550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1551]),
        .S(self_sf7[1551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1552]),
        .S(self_sf7[1552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1553]),
        .S(self_sf7[1553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1554]),
        .S(self_sf7[1554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1555]),
        .S(self_sf7[1555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1556]),
        .S(self_sf7[1556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1557]),
        .S(self_sf7[1557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1558]),
        .S(self_sf7[1558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1559]),
        .S(self_sf7[1559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[155]),
        .S(self_sf7[155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1560]),
        .S(self_sf7[1560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1561]),
        .S(self_sf7[1561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1562]),
        .S(self_sf7[1562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1563]),
        .S(self_sf7[1563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1564]),
        .S(self_sf7[1564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1565]),
        .S(self_sf7[1565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1566]),
        .S(self_sf7[1566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1567]),
        .S(self_sf7[1567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1568]),
        .S(self_sf7[1568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1569]),
        .S(self_sf7[1569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[156]),
        .S(self_sf7[156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1570]),
        .S(self_sf7[1570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1571]),
        .S(self_sf7[1571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1572]),
        .S(self_sf7[1572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1573]),
        .S(self_sf7[1573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1574]),
        .S(self_sf7[1574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1575]),
        .S(self_sf7[1575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1576]),
        .S(self_sf7[1576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1577]),
        .S(self_sf7[1577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1578]),
        .S(self_sf7[1578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1579]),
        .S(self_sf7[1579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[157]),
        .S(self_sf7[157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1580]),
        .S(self_sf7[1580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1581]),
        .S(self_sf7[1581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1582]),
        .S(self_sf7[1582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1583]),
        .S(self_sf7[1583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1584]),
        .S(self_sf7[1584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1585]),
        .S(self_sf7[1585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1586]),
        .S(self_sf7[1586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1587]),
        .S(self_sf7[1587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1588]),
        .S(self_sf7[1588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1589]),
        .S(self_sf7[1589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[158]),
        .S(self_sf7[158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1590]),
        .S(self_sf7[1590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1591]),
        .S(self_sf7[1591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1592]),
        .S(self_sf7[1592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1593]),
        .S(self_sf7[1593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1594]),
        .S(self_sf7[1594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1595]),
        .S(self_sf7[1595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1596]),
        .S(self_sf7[1596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1597]),
        .S(self_sf7[1597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1598]),
        .S(self_sf7[1598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1599]),
        .S(self_sf7[1599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[159]),
        .S(self_sf7[159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[15].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[15]),
        .S(self_sf7[15]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1600]),
        .S(self_sf7[1600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1601]),
        .S(self_sf7[1601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1602]),
        .S(self_sf7[1602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1603]),
        .S(self_sf7[1603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1604]),
        .S(self_sf7[1604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1605]),
        .S(self_sf7[1605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1606]),
        .S(self_sf7[1606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1607]),
        .S(self_sf7[1607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1608]),
        .S(self_sf7[1608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1609]),
        .S(self_sf7[1609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[160]),
        .S(self_sf7[160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1610]),
        .S(self_sf7[1610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1611]),
        .S(self_sf7[1611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1612]),
        .S(self_sf7[1612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1613]),
        .S(self_sf7[1613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1614]),
        .S(self_sf7[1614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1615]),
        .S(self_sf7[1615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1616]),
        .S(self_sf7[1616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1617]),
        .S(self_sf7[1617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1618]),
        .S(self_sf7[1618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1619]),
        .S(self_sf7[1619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[161]),
        .S(self_sf7[161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1620]),
        .S(self_sf7[1620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1621]),
        .S(self_sf7[1621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1622]),
        .S(self_sf7[1622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1623]),
        .S(self_sf7[1623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1624]),
        .S(self_sf7[1624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1625]),
        .S(self_sf7[1625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1626]),
        .S(self_sf7[1626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1627]),
        .S(self_sf7[1627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1628]),
        .S(self_sf7[1628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1629]),
        .S(self_sf7[1629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[162]),
        .S(self_sf7[162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1630]),
        .S(self_sf7[1630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1631]),
        .S(self_sf7[1631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1632]),
        .S(self_sf7[1632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1633]),
        .S(self_sf7[1633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1634]),
        .S(self_sf7[1634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1635]),
        .S(self_sf7[1635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1636]),
        .S(self_sf7[1636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1637]),
        .S(self_sf7[1637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1638]),
        .S(self_sf7[1638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1639]),
        .S(self_sf7[1639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[163]),
        .S(self_sf7[163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1640]),
        .S(self_sf7[1640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1641]),
        .S(self_sf7[1641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1642]),
        .S(self_sf7[1642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1643]),
        .S(self_sf7[1643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1644]),
        .S(self_sf7[1644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1645]),
        .S(self_sf7[1645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1646]),
        .S(self_sf7[1646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1647]),
        .S(self_sf7[1647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1648]),
        .S(self_sf7[1648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1649]),
        .S(self_sf7[1649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[164]),
        .S(self_sf7[164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1650]),
        .S(self_sf7[1650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1651]),
        .S(self_sf7[1651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1652]),
        .S(self_sf7[1652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1653]),
        .S(self_sf7[1653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1654]),
        .S(self_sf7[1654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1655]),
        .S(self_sf7[1655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1656]),
        .S(self_sf7[1656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1657]),
        .S(self_sf7[1657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1658]),
        .S(self_sf7[1658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1659]),
        .S(self_sf7[1659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[165]),
        .S(self_sf7[165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1660]),
        .S(self_sf7[1660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1661]),
        .S(self_sf7[1661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1662]),
        .S(self_sf7[1662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1663]),
        .S(self_sf7[1663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1664]),
        .S(self_sf7[1664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1665]),
        .S(self_sf7[1665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1666]),
        .S(self_sf7[1666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1667]),
        .S(self_sf7[1667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1668]),
        .S(self_sf7[1668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1669]),
        .S(self_sf7[1669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[166]),
        .S(self_sf7[166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1670]),
        .S(self_sf7[1670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1671]),
        .S(self_sf7[1671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1672]),
        .S(self_sf7[1672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1673]),
        .S(self_sf7[1673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1674]),
        .S(self_sf7[1674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1675]),
        .S(self_sf7[1675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1676]),
        .S(self_sf7[1676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1677]),
        .S(self_sf7[1677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1678]),
        .S(self_sf7[1678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1679]),
        .S(self_sf7[1679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[167]),
        .S(self_sf7[167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1680]),
        .S(self_sf7[1680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1681]),
        .S(self_sf7[1681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1682]),
        .S(self_sf7[1682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1683]),
        .S(self_sf7[1683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1684]),
        .S(self_sf7[1684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1685]),
        .S(self_sf7[1685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1686]),
        .S(self_sf7[1686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1687]),
        .S(self_sf7[1687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1688]),
        .S(self_sf7[1688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1689]),
        .S(self_sf7[1689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[168]),
        .S(self_sf7[168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1690]),
        .S(self_sf7[1690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1691]),
        .S(self_sf7[1691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1692]),
        .S(self_sf7[1692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1693]),
        .S(self_sf7[1693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1694]),
        .S(self_sf7[1694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1695]),
        .S(self_sf7[1695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1696]),
        .S(self_sf7[1696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1697]),
        .S(self_sf7[1697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1698]),
        .S(self_sf7[1698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1699]),
        .S(self_sf7[1699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[169]),
        .S(self_sf7[169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[16].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[16]),
        .S(self_sf7[16]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1700]),
        .S(self_sf7[1700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1701]),
        .S(self_sf7[1701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1702]),
        .S(self_sf7[1702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1703]),
        .S(self_sf7[1703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1704]),
        .S(self_sf7[1704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1705]),
        .S(self_sf7[1705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1706]),
        .S(self_sf7[1706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1707]),
        .S(self_sf7[1707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1708]),
        .S(self_sf7[1708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1709]),
        .S(self_sf7[1709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[170]),
        .S(self_sf7[170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1710]),
        .S(self_sf7[1710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1711]),
        .S(self_sf7[1711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1712]),
        .S(self_sf7[1712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1713]),
        .S(self_sf7[1713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1714]),
        .S(self_sf7[1714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1715]),
        .S(self_sf7[1715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1716]),
        .S(self_sf7[1716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1717]),
        .S(self_sf7[1717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1718]),
        .S(self_sf7[1718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1719]),
        .S(self_sf7[1719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[171]),
        .S(self_sf7[171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1720]),
        .S(self_sf7[1720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1721]),
        .S(self_sf7[1721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1722]),
        .S(self_sf7[1722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1723]),
        .S(self_sf7[1723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1724]),
        .S(self_sf7[1724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1725]),
        .S(self_sf7[1725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1726]),
        .S(self_sf7[1726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1727]),
        .S(self_sf7[1727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1728]),
        .S(self_sf7[1728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1729]),
        .S(self_sf7[1729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[172]),
        .S(self_sf7[172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1730]),
        .S(self_sf7[1730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1731]),
        .S(self_sf7[1731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1732]),
        .S(self_sf7[1732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1733]),
        .S(self_sf7[1733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1734]),
        .S(self_sf7[1734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1735]),
        .S(self_sf7[1735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1736]),
        .S(self_sf7[1736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1737]),
        .S(self_sf7[1737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1738]),
        .S(self_sf7[1738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1739]),
        .S(self_sf7[1739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[173]),
        .S(self_sf7[173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1740]),
        .S(self_sf7[1740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1741]),
        .S(self_sf7[1741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1742]),
        .S(self_sf7[1742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1743]),
        .S(self_sf7[1743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1744]),
        .S(self_sf7[1744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1745]),
        .S(self_sf7[1745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1746]),
        .S(self_sf7[1746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1747]),
        .S(self_sf7[1747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1748]),
        .S(self_sf7[1748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1749]),
        .S(self_sf7[1749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[174]),
        .S(self_sf7[174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1750]),
        .S(self_sf7[1750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1751]),
        .S(self_sf7[1751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1752]),
        .S(self_sf7[1752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1753]),
        .S(self_sf7[1753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1754]),
        .S(self_sf7[1754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1755]),
        .S(self_sf7[1755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1756]),
        .S(self_sf7[1756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1757]),
        .S(self_sf7[1757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1758]),
        .S(self_sf7[1758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1759]),
        .S(self_sf7[1759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[175]),
        .S(self_sf7[175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1760]),
        .S(self_sf7[1760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1761]),
        .S(self_sf7[1761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1762]),
        .S(self_sf7[1762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1763]),
        .S(self_sf7[1763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1764]),
        .S(self_sf7[1764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1765]),
        .S(self_sf7[1765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1766]),
        .S(self_sf7[1766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1767]),
        .S(self_sf7[1767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1768]),
        .S(self_sf7[1768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1769]),
        .S(self_sf7[1769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[176]),
        .S(self_sf7[176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1770]),
        .S(self_sf7[1770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1771]),
        .S(self_sf7[1771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1772]),
        .S(self_sf7[1772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1773]),
        .S(self_sf7[1773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1774]),
        .S(self_sf7[1774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1775]),
        .S(self_sf7[1775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1776]),
        .S(self_sf7[1776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1777]),
        .S(self_sf7[1777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1778]),
        .S(self_sf7[1778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1779]),
        .S(self_sf7[1779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[177]),
        .S(self_sf7[177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1780]),
        .S(self_sf7[1780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1781]),
        .S(self_sf7[1781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1782]),
        .S(self_sf7[1782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1783]),
        .S(self_sf7[1783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1784]),
        .S(self_sf7[1784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1785]),
        .S(self_sf7[1785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1786]),
        .S(self_sf7[1786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1787]),
        .S(self_sf7[1787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1788]),
        .S(self_sf7[1788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1789]),
        .S(self_sf7[1789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[178]),
        .S(self_sf7[178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1790]),
        .S(self_sf7[1790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1791]),
        .S(self_sf7[1791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1792]),
        .S(self_sf7[1792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1793]),
        .S(self_sf7[1793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1794]),
        .S(self_sf7[1794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1795]),
        .S(self_sf7[1795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1796]),
        .S(self_sf7[1796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1797]),
        .S(self_sf7[1797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1798]),
        .S(self_sf7[1798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1799]),
        .S(self_sf7[1799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[179]),
        .S(self_sf7[179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[17].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[17]),
        .S(self_sf7[17]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[180]),
        .S(self_sf7[180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[181]),
        .S(self_sf7[181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[182]),
        .S(self_sf7[182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[183]),
        .S(self_sf7[183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[184]),
        .S(self_sf7[184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[185]),
        .S(self_sf7[185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[186]),
        .S(self_sf7[186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[187]),
        .S(self_sf7[187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[188]),
        .S(self_sf7[188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[189]),
        .S(self_sf7[189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[18].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[18]),
        .S(self_sf7[18]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[190]),
        .S(self_sf7[190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[191]),
        .S(self_sf7[191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[192]),
        .S(self_sf7[192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[193]),
        .S(self_sf7[193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[194]),
        .S(self_sf7[194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[195]),
        .S(self_sf7[195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[196]),
        .S(self_sf7[196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[197]),
        .S(self_sf7[197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[198]),
        .S(self_sf7[198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[199]),
        .S(self_sf7[199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[19].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[19]),
        .S(self_sf7[19]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1]),
        .S(info_sf7[1]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[200]),
        .S(self_sf7[200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[201]),
        .S(self_sf7[201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[202]),
        .S(self_sf7[202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[203]),
        .S(self_sf7[203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[204]),
        .S(self_sf7[204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[205]),
        .S(self_sf7[205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[206]),
        .S(self_sf7[206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[207]),
        .S(self_sf7[207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[208]),
        .S(self_sf7[208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[209]),
        .S(self_sf7[209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[20].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[20]),
        .S(self_sf7[20]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[210]),
        .S(self_sf7[210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[211]),
        .S(self_sf7[211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[212]),
        .S(self_sf7[212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[213]),
        .S(self_sf7[213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[214]),
        .S(self_sf7[214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[215]),
        .S(self_sf7[215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[216]),
        .S(self_sf7[216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[217]),
        .S(self_sf7[217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[218]),
        .S(self_sf7[218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[219]),
        .S(self_sf7[219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[21].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[21]),
        .S(self_sf7[21]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[220]),
        .S(self_sf7[220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[221]),
        .S(self_sf7[221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[222]),
        .S(self_sf7[222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[223]),
        .S(self_sf7[223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[224]),
        .S(self_sf7[224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[225]),
        .S(self_sf7[225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[226]),
        .S(self_sf7[226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[227]),
        .S(self_sf7[227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[228]),
        .S(self_sf7[228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[229]),
        .S(self_sf7[229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[22].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[22]),
        .S(self_sf7[22]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[230]),
        .S(self_sf7[230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[231]),
        .S(self_sf7[231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[232]),
        .S(self_sf7[232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[233]),
        .S(self_sf7[233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[234]),
        .S(self_sf7[234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[235]),
        .S(self_sf7[235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[236]),
        .S(self_sf7[236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[237]),
        .S(self_sf7[237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[238]),
        .S(self_sf7[238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[239]),
        .S(self_sf7[239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[23].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[23]),
        .S(self_sf7[23]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[240]),
        .S(self_sf7[240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[241]),
        .S(self_sf7[241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[242]),
        .S(self_sf7[242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[243]),
        .S(self_sf7[243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[244]),
        .S(self_sf7[244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[245]),
        .S(self_sf7[245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[246]),
        .S(self_sf7[246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[247]),
        .S(self_sf7[247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[248]),
        .S(self_sf7[248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[249]),
        .S(self_sf7[249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[24].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[24]),
        .S(self_sf7[24]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[250]),
        .S(self_sf7[250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[251]),
        .S(self_sf7[251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[252]),
        .S(self_sf7[252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[253]),
        .S(self_sf7[253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[254]),
        .S(self_sf7[254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[255]),
        .S(self_sf7[255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[256]),
        .S(self_sf7[256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[257]),
        .S(self_sf7[257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[258]),
        .S(self_sf7[258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[259]),
        .S(self_sf7[259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[25].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[25]),
        .S(self_sf7[25]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[260]),
        .S(self_sf7[260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[261]),
        .S(self_sf7[261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[262]),
        .S(self_sf7[262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[263]),
        .S(self_sf7[263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[264]),
        .S(self_sf7[264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[265]),
        .S(self_sf7[265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[266]),
        .S(self_sf7[266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[267]),
        .S(self_sf7[267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[268]),
        .S(self_sf7[268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[269]),
        .S(self_sf7[269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[26].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[26]),
        .S(self_sf7[26]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[270]),
        .S(self_sf7[270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[271]),
        .S(self_sf7[271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[272]),
        .S(self_sf7[272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[273]),
        .S(self_sf7[273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[274]),
        .S(self_sf7[274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[275]),
        .S(self_sf7[275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[276]),
        .S(self_sf7[276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[277]),
        .S(self_sf7[277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[278]),
        .S(self_sf7[278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[279]),
        .S(self_sf7[279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[27].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[27]),
        .S(self_sf7[27]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[280]),
        .S(self_sf7[280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[281]),
        .S(self_sf7[281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[282]),
        .S(self_sf7[282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[283]),
        .S(self_sf7[283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[284]),
        .S(self_sf7[284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[285]),
        .S(self_sf7[285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[286]),
        .S(self_sf7[286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[287]),
        .S(self_sf7[287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[288]),
        .S(self_sf7[288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[289]),
        .S(self_sf7[289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[28].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[28]),
        .S(self_sf7[28]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[290]),
        .S(self_sf7[290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[291]),
        .S(self_sf7[291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[292]),
        .S(self_sf7[292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[293]),
        .S(self_sf7[293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[294]),
        .S(self_sf7[294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[295]),
        .S(self_sf7[295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[296]),
        .S(self_sf7[296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[297]),
        .S(self_sf7[297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[298]),
        .S(self_sf7[298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[299]),
        .S(self_sf7[299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[29].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[29]),
        .S(self_sf7[29]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[2].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[2]),
        .S(info_sf7[2]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[300]),
        .S(self_sf7[300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[301]),
        .S(self_sf7[301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[302]),
        .S(self_sf7[302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[303]),
        .S(self_sf7[303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[304]),
        .S(self_sf7[304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[305]),
        .S(self_sf7[305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[306]),
        .S(self_sf7[306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[307]),
        .S(self_sf7[307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[308]),
        .S(self_sf7[308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[309]),
        .S(self_sf7[309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[30].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[30]),
        .S(self_sf7[30]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[310]),
        .S(self_sf7[310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[311]),
        .S(self_sf7[311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[312]),
        .S(self_sf7[312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[313]),
        .S(self_sf7[313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[314]),
        .S(self_sf7[314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[315]),
        .S(self_sf7[315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[316]),
        .S(self_sf7[316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[317]),
        .S(self_sf7[317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[318]),
        .S(self_sf7[318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[319]),
        .S(self_sf7[319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[31].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[31]),
        .S(self_sf7[31]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[320]),
        .S(self_sf7[320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[321]),
        .S(self_sf7[321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[322]),
        .S(self_sf7[322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[323]),
        .S(self_sf7[323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[324]),
        .S(self_sf7[324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[325]),
        .S(self_sf7[325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[326]),
        .S(self_sf7[326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[327]),
        .S(self_sf7[327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[328]),
        .S(self_sf7[328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[329]),
        .S(self_sf7[329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[32].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[32]),
        .S(self_sf7[32]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[330]),
        .S(self_sf7[330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[331]),
        .S(self_sf7[331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[332]),
        .S(self_sf7[332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[333]),
        .S(self_sf7[333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[334]),
        .S(self_sf7[334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[335]),
        .S(self_sf7[335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[336]),
        .S(self_sf7[336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[337]),
        .S(self_sf7[337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[338]),
        .S(self_sf7[338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[339]),
        .S(self_sf7[339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[33].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[33]),
        .S(self_sf7[33]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[340]),
        .S(self_sf7[340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[341]),
        .S(self_sf7[341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[342]),
        .S(self_sf7[342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[343]),
        .S(self_sf7[343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[344]),
        .S(self_sf7[344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[345]),
        .S(self_sf7[345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[346]),
        .S(self_sf7[346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[347]),
        .S(self_sf7[347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[348]),
        .S(self_sf7[348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[349]),
        .S(self_sf7[349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[34].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[34]),
        .S(self_sf7[34]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[350]),
        .S(self_sf7[350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[351]),
        .S(self_sf7[351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[352]),
        .S(self_sf7[352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[353]),
        .S(self_sf7[353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[354]),
        .S(self_sf7[354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[355]),
        .S(self_sf7[355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[356]),
        .S(self_sf7[356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[357]),
        .S(self_sf7[357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[358]),
        .S(self_sf7[358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[359]),
        .S(self_sf7[359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[35].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[35]),
        .S(self_sf7[35]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[360]),
        .S(self_sf7[360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[361]),
        .S(self_sf7[361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[362]),
        .S(self_sf7[362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[363]),
        .S(self_sf7[363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[364]),
        .S(self_sf7[364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[365]),
        .S(self_sf7[365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[366]),
        .S(self_sf7[366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[367]),
        .S(self_sf7[367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[368]),
        .S(self_sf7[368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[369]),
        .S(self_sf7[369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[36].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[36]),
        .S(self_sf7[36]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[370]),
        .S(self_sf7[370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[371]),
        .S(self_sf7[371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[372]),
        .S(self_sf7[372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[373]),
        .S(self_sf7[373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[374]),
        .S(self_sf7[374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[375]),
        .S(self_sf7[375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[376]),
        .S(self_sf7[376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[377]),
        .S(self_sf7[377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[378]),
        .S(self_sf7[378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[379]),
        .S(self_sf7[379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[37].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[37]),
        .S(self_sf7[37]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[380]),
        .S(self_sf7[380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[381]),
        .S(self_sf7[381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[382]),
        .S(self_sf7[382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[383]),
        .S(self_sf7[383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[384]),
        .S(self_sf7[384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[385]),
        .S(self_sf7[385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[386]),
        .S(self_sf7[386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[387]),
        .S(self_sf7[387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[388]),
        .S(self_sf7[388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[389]),
        .S(self_sf7[389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[38].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[38]),
        .S(self_sf7[38]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[390]),
        .S(self_sf7[390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[391]),
        .S(self_sf7[391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[392]),
        .S(self_sf7[392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[393]),
        .S(self_sf7[393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[394]),
        .S(self_sf7[394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[395]),
        .S(self_sf7[395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[396]),
        .S(self_sf7[396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[397]),
        .S(self_sf7[397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[398]),
        .S(self_sf7[398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[399]),
        .S(self_sf7[399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[39].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[39]),
        .S(self_sf7[39]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[3].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[3]),
        .S(info_sf7[3]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[400]),
        .S(self_sf7[400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[401]),
        .S(self_sf7[401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[402]),
        .S(self_sf7[402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[403]),
        .S(self_sf7[403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[404]),
        .S(self_sf7[404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[405]),
        .S(self_sf7[405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[406]),
        .S(self_sf7[406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[407]),
        .S(self_sf7[407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[408]),
        .S(self_sf7[408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[409]),
        .S(self_sf7[409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[40].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[40]),
        .S(self_sf7[40]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[410]),
        .S(self_sf7[410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[411]),
        .S(self_sf7[411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[412]),
        .S(self_sf7[412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[413]),
        .S(self_sf7[413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[414]),
        .S(self_sf7[414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[415]),
        .S(self_sf7[415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[416]),
        .S(self_sf7[416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[417]),
        .S(self_sf7[417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[418]),
        .S(self_sf7[418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[419]),
        .S(self_sf7[419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[41].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[41]),
        .S(self_sf7[41]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[420]),
        .S(self_sf7[420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[421]),
        .S(self_sf7[421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[422]),
        .S(self_sf7[422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[423]),
        .S(self_sf7[423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[424]),
        .S(self_sf7[424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[425]),
        .S(self_sf7[425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[426]),
        .S(self_sf7[426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[427]),
        .S(self_sf7[427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[428]),
        .S(self_sf7[428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[429]),
        .S(self_sf7[429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[42].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[42]),
        .S(self_sf7[42]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[430]),
        .S(self_sf7[430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[431]),
        .S(self_sf7[431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[432]),
        .S(self_sf7[432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[433]),
        .S(self_sf7[433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[434]),
        .S(self_sf7[434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[435]),
        .S(self_sf7[435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[436]),
        .S(self_sf7[436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[437]),
        .S(self_sf7[437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[438]),
        .S(self_sf7[438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[439]),
        .S(self_sf7[439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[43].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[43]),
        .S(self_sf7[43]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[440]),
        .S(self_sf7[440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[441]),
        .S(self_sf7[441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[442]),
        .S(self_sf7[442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[443]),
        .S(self_sf7[443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[444]),
        .S(self_sf7[444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[445]),
        .S(self_sf7[445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[446]),
        .S(self_sf7[446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[447]),
        .S(self_sf7[447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[448]),
        .S(self_sf7[448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[449]),
        .S(self_sf7[449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[44].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[44]),
        .S(self_sf7[44]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[450]),
        .S(self_sf7[450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[451]),
        .S(self_sf7[451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[452]),
        .S(self_sf7[452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[453]),
        .S(self_sf7[453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[454]),
        .S(self_sf7[454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[455]),
        .S(self_sf7[455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[456]),
        .S(self_sf7[456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[457]),
        .S(self_sf7[457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[458]),
        .S(self_sf7[458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[459]),
        .S(self_sf7[459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[45].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[45]),
        .S(self_sf7[45]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[460]),
        .S(self_sf7[460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[461]),
        .S(self_sf7[461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[462]),
        .S(self_sf7[462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[463]),
        .S(self_sf7[463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[464]),
        .S(self_sf7[464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[465]),
        .S(self_sf7[465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[466]),
        .S(self_sf7[466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[467]),
        .S(self_sf7[467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[468]),
        .S(self_sf7[468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[469]),
        .S(self_sf7[469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[46].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[46]),
        .S(self_sf7[46]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[470]),
        .S(self_sf7[470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[471]),
        .S(self_sf7[471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[472]),
        .S(self_sf7[472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[473]),
        .S(self_sf7[473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[474]),
        .S(self_sf7[474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[475]),
        .S(self_sf7[475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[476]),
        .S(self_sf7[476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[477]),
        .S(self_sf7[477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[478]),
        .S(self_sf7[478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[479]),
        .S(self_sf7[479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[47].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[47]),
        .S(self_sf7[47]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[480]),
        .S(self_sf7[480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[481]),
        .S(self_sf7[481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[482]),
        .S(self_sf7[482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[483]),
        .S(self_sf7[483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[484]),
        .S(self_sf7[484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[485]),
        .S(self_sf7[485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[486]),
        .S(self_sf7[486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[487]),
        .S(self_sf7[487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[488]),
        .S(self_sf7[488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[489]),
        .S(self_sf7[489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[48].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[48]),
        .S(self_sf7[48]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[490]),
        .S(self_sf7[490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[491]),
        .S(self_sf7[491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[492]),
        .S(self_sf7[492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[493]),
        .S(self_sf7[493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[494]),
        .S(self_sf7[494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[495]),
        .S(self_sf7[495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[496]),
        .S(self_sf7[496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[497]),
        .S(self_sf7[497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[498]),
        .S(self_sf7[498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[499]),
        .S(self_sf7[499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[49].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[49]),
        .S(self_sf7[49]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[4].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[4]),
        .S(info_sf7[4]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[500]),
        .S(self_sf7[500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[501]),
        .S(self_sf7[501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[502]),
        .S(self_sf7[502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[503]),
        .S(self_sf7[503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[504]),
        .S(self_sf7[504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[505]),
        .S(self_sf7[505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[506]),
        .S(self_sf7[506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[507]),
        .S(self_sf7[507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[508]),
        .S(self_sf7[508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[509]),
        .S(self_sf7[509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[50].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[50]),
        .S(self_sf7[50]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[510]),
        .S(self_sf7[510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[511]),
        .S(self_sf7[511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[512]),
        .S(self_sf7[512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[513]),
        .S(self_sf7[513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[514]),
        .S(self_sf7[514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[515]),
        .S(self_sf7[515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[516]),
        .S(self_sf7[516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[517]),
        .S(self_sf7[517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[518]),
        .S(self_sf7[518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[519]),
        .S(self_sf7[519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[51].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[51]),
        .S(self_sf7[51]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[520]),
        .S(self_sf7[520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[521]),
        .S(self_sf7[521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[522]),
        .S(self_sf7[522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[523]),
        .S(self_sf7[523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[524]),
        .S(self_sf7[524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[525]),
        .S(self_sf7[525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[526]),
        .S(self_sf7[526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[527]),
        .S(self_sf7[527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[528]),
        .S(self_sf7[528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[529]),
        .S(self_sf7[529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[52].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[52]),
        .S(self_sf7[52]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[530]),
        .S(self_sf7[530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[531]),
        .S(self_sf7[531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[532]),
        .S(self_sf7[532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[533]),
        .S(self_sf7[533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[534]),
        .S(self_sf7[534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[535]),
        .S(self_sf7[535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[536]),
        .S(self_sf7[536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[537]),
        .S(self_sf7[537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[538]),
        .S(self_sf7[538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[539]),
        .S(self_sf7[539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[53].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[53]),
        .S(self_sf7[53]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[540]),
        .S(self_sf7[540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[541]),
        .S(self_sf7[541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[542]),
        .S(self_sf7[542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[543]),
        .S(self_sf7[543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[544]),
        .S(self_sf7[544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[545]),
        .S(self_sf7[545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[546]),
        .S(self_sf7[546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[547]),
        .S(self_sf7[547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[548]),
        .S(self_sf7[548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[549]),
        .S(self_sf7[549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[54].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[54]),
        .S(self_sf7[54]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[550]),
        .S(self_sf7[550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[551]),
        .S(self_sf7[551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[552]),
        .S(self_sf7[552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[553]),
        .S(self_sf7[553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[554]),
        .S(self_sf7[554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[555]),
        .S(self_sf7[555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[556]),
        .S(self_sf7[556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[557]),
        .S(self_sf7[557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[558]),
        .S(self_sf7[558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[559]),
        .S(self_sf7[559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[55].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[55]),
        .S(self_sf7[55]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[560]),
        .S(self_sf7[560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[561]),
        .S(self_sf7[561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[562]),
        .S(self_sf7[562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[563]),
        .S(self_sf7[563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[564]),
        .S(self_sf7[564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[565]),
        .S(self_sf7[565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[566]),
        .S(self_sf7[566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[567]),
        .S(self_sf7[567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[568]),
        .S(self_sf7[568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[569]),
        .S(self_sf7[569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[56].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[56]),
        .S(self_sf7[56]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[570]),
        .S(self_sf7[570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[571]),
        .S(self_sf7[571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[572]),
        .S(self_sf7[572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[573]),
        .S(self_sf7[573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[574]),
        .S(self_sf7[574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[575]),
        .S(self_sf7[575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[576]),
        .S(self_sf7[576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[577]),
        .S(self_sf7[577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[578]),
        .S(self_sf7[578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[579]),
        .S(self_sf7[579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[57].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[57]),
        .S(self_sf7[57]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[580]),
        .S(self_sf7[580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[581]),
        .S(self_sf7[581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[582]),
        .S(self_sf7[582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[583]),
        .S(self_sf7[583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[584]),
        .S(self_sf7[584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[585]),
        .S(self_sf7[585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[586]),
        .S(self_sf7[586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[587]),
        .S(self_sf7[587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[588]),
        .S(self_sf7[588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[589]),
        .S(self_sf7[589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[58].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[58]),
        .S(self_sf7[58]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[590]),
        .S(self_sf7[590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[591]),
        .S(self_sf7[591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[592]),
        .S(self_sf7[592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[593]),
        .S(self_sf7[593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[594]),
        .S(self_sf7[594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[595]),
        .S(self_sf7[595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[596]),
        .S(self_sf7[596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[597]),
        .S(self_sf7[597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[598]),
        .S(self_sf7[598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[599]),
        .S(self_sf7[599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[59].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[59]),
        .S(self_sf7[59]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[5].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[5]),
        .S(info_sf7[5]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[600]),
        .S(self_sf7[600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[601]),
        .S(self_sf7[601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[602]),
        .S(self_sf7[602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[603]),
        .S(self_sf7[603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[604]),
        .S(self_sf7[604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[605]),
        .S(self_sf7[605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[606]),
        .S(self_sf7[606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[607]),
        .S(self_sf7[607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[608]),
        .S(self_sf7[608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[609]),
        .S(self_sf7[609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[60].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[60]),
        .S(self_sf7[60]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[610]),
        .S(self_sf7[610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[611]),
        .S(self_sf7[611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[612]),
        .S(self_sf7[612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[613]),
        .S(self_sf7[613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[614]),
        .S(self_sf7[614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[615]),
        .S(self_sf7[615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[616]),
        .S(self_sf7[616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[617]),
        .S(self_sf7[617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[618]),
        .S(self_sf7[618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[619]),
        .S(self_sf7[619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[61].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[61]),
        .S(self_sf7[61]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[620]),
        .S(self_sf7[620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[621]),
        .S(self_sf7[621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[622]),
        .S(self_sf7[622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[623]),
        .S(self_sf7[623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[624]),
        .S(self_sf7[624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[625]),
        .S(self_sf7[625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[626]),
        .S(self_sf7[626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[627]),
        .S(self_sf7[627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[628]),
        .S(self_sf7[628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[629]),
        .S(self_sf7[629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[62].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[62]),
        .S(self_sf7[62]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[630]),
        .S(self_sf7[630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[631]),
        .S(self_sf7[631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[632]),
        .S(self_sf7[632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[633]),
        .S(self_sf7[633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[634]),
        .S(self_sf7[634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[635]),
        .S(self_sf7[635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[636]),
        .S(self_sf7[636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[637]),
        .S(self_sf7[637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[638]),
        .S(self_sf7[638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[639]),
        .S(self_sf7[639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[63].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[63]),
        .S(self_sf7[63]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[640]),
        .S(self_sf7[640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[641]),
        .S(self_sf7[641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[642]),
        .S(self_sf7[642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[643]),
        .S(self_sf7[643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[644]),
        .S(self_sf7[644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[645]),
        .S(self_sf7[645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[646]),
        .S(self_sf7[646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[647]),
        .S(self_sf7[647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[648]),
        .S(self_sf7[648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[649]),
        .S(self_sf7[649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[64].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[64]),
        .S(self_sf7[64]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[650]),
        .S(self_sf7[650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[651]),
        .S(self_sf7[651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[652]),
        .S(self_sf7[652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[653]),
        .S(self_sf7[653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[654]),
        .S(self_sf7[654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[655]),
        .S(self_sf7[655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[656]),
        .S(self_sf7[656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[657]),
        .S(self_sf7[657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[658]),
        .S(self_sf7[658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[659]),
        .S(self_sf7[659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[65].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[65]),
        .S(self_sf7[65]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[660]),
        .S(self_sf7[660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[661]),
        .S(self_sf7[661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[662]),
        .S(self_sf7[662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[663]),
        .S(self_sf7[663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[664]),
        .S(self_sf7[664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[665]),
        .S(self_sf7[665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[666]),
        .S(self_sf7[666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[667]),
        .S(self_sf7[667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[668]),
        .S(self_sf7[668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[669]),
        .S(self_sf7[669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[66].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[66]),
        .S(self_sf7[66]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[670]),
        .S(self_sf7[670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[671]),
        .S(self_sf7[671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[672]),
        .S(self_sf7[672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[673]),
        .S(self_sf7[673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[674]),
        .S(self_sf7[674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[675]),
        .S(self_sf7[675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[676]),
        .S(self_sf7[676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[677]),
        .S(self_sf7[677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[678]),
        .S(self_sf7[678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[679]),
        .S(self_sf7[679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[67].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[67]),
        .S(self_sf7[67]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[680]),
        .S(self_sf7[680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[681]),
        .S(self_sf7[681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[682]),
        .S(self_sf7[682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[683]),
        .S(self_sf7[683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[684]),
        .S(self_sf7[684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[685]),
        .S(self_sf7[685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[686]),
        .S(self_sf7[686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[687]),
        .S(self_sf7[687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[688]),
        .S(self_sf7[688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[689]),
        .S(self_sf7[689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[68].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[68]),
        .S(self_sf7[68]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[690]),
        .S(self_sf7[690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[691]),
        .S(self_sf7[691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[692]),
        .S(self_sf7[692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[693]),
        .S(self_sf7[693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[694]),
        .S(self_sf7[694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[695]),
        .S(self_sf7[695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[696]),
        .S(self_sf7[696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[697]),
        .S(self_sf7[697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[698]),
        .S(self_sf7[698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[699]),
        .S(self_sf7[699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[69].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[69]),
        .S(self_sf7[69]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[6].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[6]),
        .S(info_sf7[6]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[700]),
        .S(self_sf7[700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[701]),
        .S(self_sf7[701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[702]),
        .S(self_sf7[702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[703]),
        .S(self_sf7[703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[704]),
        .S(self_sf7[704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[705]),
        .S(self_sf7[705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[706]),
        .S(self_sf7[706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[707]),
        .S(self_sf7[707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[708]),
        .S(self_sf7[708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[709]),
        .S(self_sf7[709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[70].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[70]),
        .S(self_sf7[70]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[710]),
        .S(self_sf7[710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[711]),
        .S(self_sf7[711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[712]),
        .S(self_sf7[712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[713]),
        .S(self_sf7[713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[714]),
        .S(self_sf7[714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[715]),
        .S(self_sf7[715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[716]),
        .S(self_sf7[716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[717]),
        .S(self_sf7[717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[718]),
        .S(self_sf7[718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[719]),
        .S(self_sf7[719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[71].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[71]),
        .S(self_sf7[71]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[720]),
        .S(self_sf7[720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[721]),
        .S(self_sf7[721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[722]),
        .S(self_sf7[722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[723]),
        .S(self_sf7[723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[724]),
        .S(self_sf7[724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[725]),
        .S(self_sf7[725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[726]),
        .S(self_sf7[726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[727]),
        .S(self_sf7[727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[728]),
        .S(self_sf7[728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[729]),
        .S(self_sf7[729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[72].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[72]),
        .S(self_sf7[72]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[730]),
        .S(self_sf7[730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[731]),
        .S(self_sf7[731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[732]),
        .S(self_sf7[732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[733]),
        .S(self_sf7[733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[734]),
        .S(self_sf7[734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[735]),
        .S(self_sf7[735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[736]),
        .S(self_sf7[736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[737]),
        .S(self_sf7[737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[738]),
        .S(self_sf7[738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[739]),
        .S(self_sf7[739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[73].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[73]),
        .S(self_sf7[73]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[740]),
        .S(self_sf7[740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[741]),
        .S(self_sf7[741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[742]),
        .S(self_sf7[742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[743]),
        .S(self_sf7[743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[744]),
        .S(self_sf7[744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[745]),
        .S(self_sf7[745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[746]),
        .S(self_sf7[746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[747]),
        .S(self_sf7[747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[748]),
        .S(self_sf7[748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[749]),
        .S(self_sf7[749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[74].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[74]),
        .S(self_sf7[74]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[750]),
        .S(self_sf7[750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[751]),
        .S(self_sf7[751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[752]),
        .S(self_sf7[752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[753]),
        .S(self_sf7[753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[754]),
        .S(self_sf7[754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[755]),
        .S(self_sf7[755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[756]),
        .S(self_sf7[756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[757]),
        .S(self_sf7[757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[758]),
        .S(self_sf7[758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[759]),
        .S(self_sf7[759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[75].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[75]),
        .S(self_sf7[75]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[760]),
        .S(self_sf7[760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[761]),
        .S(self_sf7[761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[762]),
        .S(self_sf7[762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[763]),
        .S(self_sf7[763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[764]),
        .S(self_sf7[764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[765]),
        .S(self_sf7[765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[766]),
        .S(self_sf7[766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[767]),
        .S(self_sf7[767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[768]),
        .S(self_sf7[768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[769]),
        .S(self_sf7[769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[76].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[76]),
        .S(self_sf7[76]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[770]),
        .S(self_sf7[770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[771]),
        .S(self_sf7[771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[772]),
        .S(self_sf7[772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[773]),
        .S(self_sf7[773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[774]),
        .S(self_sf7[774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[775]),
        .S(self_sf7[775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[776]),
        .S(self_sf7[776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[777]),
        .S(self_sf7[777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[778]),
        .S(self_sf7[778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[779]),
        .S(self_sf7[779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[77].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[77]),
        .S(self_sf7[77]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[780]),
        .S(self_sf7[780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[781]),
        .S(self_sf7[781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[782]),
        .S(self_sf7[782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[783]),
        .S(self_sf7[783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[784]),
        .S(self_sf7[784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[785]),
        .S(self_sf7[785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[786]),
        .S(self_sf7[786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[787]),
        .S(self_sf7[787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[788]),
        .S(self_sf7[788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[789]),
        .S(self_sf7[789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[78].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[78]),
        .S(self_sf7[78]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[790]),
        .S(self_sf7[790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[791]),
        .S(self_sf7[791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[792]),
        .S(self_sf7[792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[793]),
        .S(self_sf7[793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[794]),
        .S(self_sf7[794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[795]),
        .S(self_sf7[795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[796]),
        .S(self_sf7[796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[797]),
        .S(self_sf7[797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[798]),
        .S(self_sf7[798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[799]),
        .S(self_sf7[799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[79].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[79]),
        .S(self_sf7[79]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[7].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[7]),
        .S(info_sf7[7]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[800].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[800]),
        .S(self_sf7[800]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[801].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[801]),
        .S(self_sf7[801]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[802].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[802]),
        .S(self_sf7[802]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[803].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[803]),
        .S(self_sf7[803]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[804].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[804]),
        .S(self_sf7[804]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[805].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[805]),
        .S(self_sf7[805]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[806].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[806]),
        .S(self_sf7[806]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[807].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[807]),
        .S(self_sf7[807]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[808].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[808]),
        .S(self_sf7[808]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[809].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[809]),
        .S(self_sf7[809]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[80].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[80]),
        .S(self_sf7[80]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[810].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[810]),
        .S(self_sf7[810]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[811].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[811]),
        .S(self_sf7[811]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[812].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[812]),
        .S(self_sf7[812]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[813].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[813]),
        .S(self_sf7[813]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[814].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[814]),
        .S(self_sf7[814]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[815].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[815]),
        .S(self_sf7[815]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[816].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[816]),
        .S(self_sf7[816]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[817].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[817]),
        .S(self_sf7[817]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[818].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[818]),
        .S(self_sf7[818]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[819].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[819]),
        .S(self_sf7[819]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[81].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[81]),
        .S(self_sf7[81]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[820].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[820]),
        .S(self_sf7[820]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[821].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[821]),
        .S(self_sf7[821]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[822].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[822]),
        .S(self_sf7[822]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[823].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[823]),
        .S(self_sf7[823]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[824].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[824]),
        .S(self_sf7[824]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[825].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[825]),
        .S(self_sf7[825]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[826].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[826]),
        .S(self_sf7[826]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[827].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[827]),
        .S(self_sf7[827]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[828].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[828]),
        .S(self_sf7[828]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[829].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[829]),
        .S(self_sf7[829]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[82].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[82]),
        .S(self_sf7[82]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[830].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[830]),
        .S(self_sf7[830]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[831].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[831]),
        .S(self_sf7[831]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[832].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[832]),
        .S(self_sf7[832]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[833].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[833]),
        .S(self_sf7[833]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[834].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[834]),
        .S(self_sf7[834]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[835].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[835]),
        .S(self_sf7[835]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[836].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[836]),
        .S(self_sf7[836]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[837].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[837]),
        .S(self_sf7[837]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[838].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[838]),
        .S(self_sf7[838]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[839].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[839]),
        .S(self_sf7[839]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[83].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[83]),
        .S(self_sf7[83]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[840].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[840]),
        .S(self_sf7[840]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[841].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[841]),
        .S(self_sf7[841]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[842].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[842]),
        .S(self_sf7[842]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[843].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[843]),
        .S(self_sf7[843]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[844].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[844]),
        .S(self_sf7[844]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[845].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[845]),
        .S(self_sf7[845]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[846].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[846]),
        .S(self_sf7[846]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[847].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[847]),
        .S(self_sf7[847]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[848].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[848]),
        .S(self_sf7[848]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[849].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[849]),
        .S(self_sf7[849]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[84].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[84]),
        .S(self_sf7[84]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[850].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[850]),
        .S(self_sf7[850]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[851].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[851]),
        .S(self_sf7[851]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[852].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[852]),
        .S(self_sf7[852]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[853].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[853]),
        .S(self_sf7[853]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[854].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[854]),
        .S(self_sf7[854]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[855].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[855]),
        .S(self_sf7[855]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[856].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[856]),
        .S(self_sf7[856]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[857].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[857]),
        .S(self_sf7[857]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[858].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[858]),
        .S(self_sf7[858]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[859].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[859]),
        .S(self_sf7[859]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[85].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[85]),
        .S(self_sf7[85]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[860].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[860]),
        .S(self_sf7[860]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[861].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[861]),
        .S(self_sf7[861]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[862].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[862]),
        .S(self_sf7[862]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[863].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[863]),
        .S(self_sf7[863]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[864].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[864]),
        .S(self_sf7[864]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[865].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[865]),
        .S(self_sf7[865]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[866].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[866]),
        .S(self_sf7[866]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[867].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[867]),
        .S(self_sf7[867]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[868].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[868]),
        .S(self_sf7[868]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[869].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[869]),
        .S(self_sf7[869]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[86].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[86]),
        .S(self_sf7[86]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[870].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[870]),
        .S(self_sf7[870]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[871].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[871]),
        .S(self_sf7[871]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[872].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[872]),
        .S(self_sf7[872]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[873].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[873]),
        .S(self_sf7[873]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[874].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[874]),
        .S(self_sf7[874]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[875].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[875]),
        .S(self_sf7[875]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[876].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[876]),
        .S(self_sf7[876]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[877].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[877]),
        .S(self_sf7[877]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[878].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[878]),
        .S(self_sf7[878]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[879].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[879]),
        .S(self_sf7[879]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[87].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[87]),
        .S(self_sf7[87]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[880].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[880]),
        .S(self_sf7[880]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[881].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[881]),
        .S(self_sf7[881]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[882].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[882]),
        .S(self_sf7[882]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[883].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[883]),
        .S(self_sf7[883]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[884].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[884]),
        .S(self_sf7[884]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[885].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[885]),
        .S(self_sf7[885]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[886].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[886]),
        .S(self_sf7[886]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[887].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[887]),
        .S(self_sf7[887]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[888].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[888]),
        .S(self_sf7[888]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[889].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[889]),
        .S(self_sf7[889]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[88].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[88]),
        .S(self_sf7[88]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[890].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[890]),
        .S(self_sf7[890]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[891].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[891]),
        .S(self_sf7[891]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[892].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[892]),
        .S(self_sf7[892]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[893].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[893]),
        .S(self_sf7[893]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[894].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[894]),
        .S(self_sf7[894]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[895].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[895]),
        .S(self_sf7[895]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[896].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[896]),
        .S(self_sf7[896]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[897].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[897]),
        .S(self_sf7[897]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[898].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[898]),
        .S(self_sf7[898]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[899].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[899]),
        .S(self_sf7[899]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[89].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[89]),
        .S(self_sf7[89]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[8].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[8]),
        .S(self_sf7[8]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[900].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[900]),
        .S(self_sf7[900]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[901].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[901]),
        .S(self_sf7[901]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[902].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[902]),
        .S(self_sf7[902]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[903].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[903]),
        .S(self_sf7[903]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[904].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[904]),
        .S(self_sf7[904]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[905].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[905]),
        .S(self_sf7[905]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[906].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[906]),
        .S(self_sf7[906]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[907].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[907]),
        .S(self_sf7[907]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[908].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[908]),
        .S(self_sf7[908]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[909].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[909]),
        .S(self_sf7[909]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[90].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[90]),
        .S(self_sf7[90]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[910].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[910]),
        .S(self_sf7[910]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[911].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[911]),
        .S(self_sf7[911]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[912].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[912]),
        .S(self_sf7[912]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[913].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[913]),
        .S(self_sf7[913]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[914].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[914]),
        .S(self_sf7[914]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[915].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[915]),
        .S(self_sf7[915]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[916].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[916]),
        .S(self_sf7[916]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[917].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[917]),
        .S(self_sf7[917]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[918].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[918]),
        .S(self_sf7[918]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[919].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[919]),
        .S(self_sf7[919]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[91].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[91]),
        .S(self_sf7[91]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[920].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[920]),
        .S(self_sf7[920]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[921].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[921]),
        .S(self_sf7[921]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[922].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[922]),
        .S(self_sf7[922]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[923].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[923]),
        .S(self_sf7[923]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[924].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[924]),
        .S(self_sf7[924]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[925].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[925]),
        .S(self_sf7[925]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[926].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[926]),
        .S(self_sf7[926]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[927].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[927]),
        .S(self_sf7[927]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[928].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[928]),
        .S(self_sf7[928]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[929].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[929]),
        .S(self_sf7[929]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[92].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[92]),
        .S(self_sf7[92]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[930].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[930]),
        .S(self_sf7[930]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[931].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[931]),
        .S(self_sf7[931]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[932].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[932]),
        .S(self_sf7[932]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[933].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[933]),
        .S(self_sf7[933]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[934].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[934]),
        .S(self_sf7[934]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[935].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[935]),
        .S(self_sf7[935]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[936].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[936]),
        .S(self_sf7[936]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[937].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[937]),
        .S(self_sf7[937]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[938].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[938]),
        .S(self_sf7[938]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[939].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[939]),
        .S(self_sf7[939]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[93].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[93]),
        .S(self_sf7[93]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[940].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[940]),
        .S(self_sf7[940]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[941].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[941]),
        .S(self_sf7[941]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[942].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[942]),
        .S(self_sf7[942]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[943].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[943]),
        .S(self_sf7[943]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[944].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[944]),
        .S(self_sf7[944]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[945].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[945]),
        .S(self_sf7[945]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[946].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[946]),
        .S(self_sf7[946]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[947].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[947]),
        .S(self_sf7[947]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[948].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[948]),
        .S(self_sf7[948]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[949].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[949]),
        .S(self_sf7[949]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[94].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[94]),
        .S(self_sf7[94]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[950].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[950]),
        .S(self_sf7[950]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[951].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[951]),
        .S(self_sf7[951]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[952].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[952]),
        .S(self_sf7[952]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[953].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[953]),
        .S(self_sf7[953]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[954].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[954]),
        .S(self_sf7[954]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[955].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[955]),
        .S(self_sf7[955]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[956].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[956]),
        .S(self_sf7[956]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[957].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[957]),
        .S(self_sf7[957]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[958].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[958]),
        .S(self_sf7[958]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[959].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[959]),
        .S(self_sf7[959]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[95].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[95]),
        .S(self_sf7[95]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[960].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[960]),
        .S(self_sf7[960]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[961].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[961]),
        .S(self_sf7[961]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[962].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[962]),
        .S(self_sf7[962]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[963].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[963]),
        .S(self_sf7[963]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[964].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[964]),
        .S(self_sf7[964]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[965].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[965]),
        .S(self_sf7[965]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[966].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[966]),
        .S(self_sf7[966]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[967].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[967]),
        .S(self_sf7[967]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[968].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[968]),
        .S(self_sf7[968]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[969].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[969]),
        .S(self_sf7[969]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[96].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[96]),
        .S(self_sf7[96]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[970].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[970]),
        .S(self_sf7[970]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[971].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[971]),
        .S(self_sf7[971]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[972].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[972]),
        .S(self_sf7[972]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[973].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[973]),
        .S(self_sf7[973]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[974].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[974]),
        .S(self_sf7[974]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[975].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[975]),
        .S(self_sf7[975]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[976].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[976]),
        .S(self_sf7[976]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[977].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[977]),
        .S(self_sf7[977]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[978].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[978]),
        .S(self_sf7[978]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[979].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[979]),
        .S(self_sf7[979]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[97].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[97]),
        .S(self_sf7[97]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[980].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[980]),
        .S(self_sf7[980]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[981].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[981]),
        .S(self_sf7[981]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[982].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[982]),
        .S(self_sf7[982]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[983].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[983]),
        .S(self_sf7[983]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[984].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[984]),
        .S(self_sf7[984]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[985].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[985]),
        .S(self_sf7[985]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[986].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[986]),
        .S(self_sf7[986]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[987].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[987]),
        .S(self_sf7[987]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[988].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[988]),
        .S(self_sf7[988]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[989].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[989]),
        .S(self_sf7[989]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[98].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[98]),
        .S(self_sf7[98]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[990].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[990]),
        .S(self_sf7[990]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[991].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[991]),
        .S(self_sf7[991]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[992].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[992]),
        .S(self_sf7[992]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[993].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[993]),
        .S(self_sf7[993]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[994].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[994]),
        .S(self_sf7[994]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[995].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[995]),
        .S(self_sf7[995]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[996].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[996]),
        .S(self_sf7[996]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[997].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[997]),
        .S(self_sf7[997]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[998].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[998]),
        .S(self_sf7[998]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[999].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[999]),
        .S(self_sf7[999]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[99].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[99]),
        .S(self_sf7[99]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[9].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[9]),
        .S(self_sf7[9]));
  (* BOX_TYPE = "black_box" *) 
  MUXF8 \activity_ROsf8[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf8[0]),
        .S(self_sf8[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF9 \activity_ROsf9[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf9[0]),
        .S(self_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_0
       (.I0(1'b0),
        .O(self_sf7[1802]));
  LUT1 #(
    .INIT(2'h2)) 
    i_1
       (.I0(1'b0),
        .O(self_sf7[1801]));
  LUT1 #(
    .INIT(2'h2)) 
    i_10
       (.I0(1'b0),
        .O(info_sf8[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_11
       (.I0(1'b0),
        .O(info_sf8[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_12
       (.I0(1'b0),
        .O(info_sf8[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_13
       (.I0(1'b0),
        .O(info_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_14
       (.I0(1'b0),
        .O(info_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_15
       (.I0(1'b0),
        .O(info_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_16
       (.I0(1'b0),
        .O(info_sf8[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_17
       (.I0(1'b0),
        .O(info_sf9[7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_18
       (.I0(1'b0),
        .O(info_sf9[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_19
       (.I0(1'b0),
        .O(info_sf9[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_2
       (.I0(1'b0),
        .O(self_sf7[1800]));
  LUT1 #(
    .INIT(2'h2)) 
    i_20
       (.I0(1'b0),
        .O(info_sf9[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_21
       (.I0(1'b0),
        .O(info_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_22
       (.I0(1'b0),
        .O(info_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_23
       (.I0(1'b0),
        .O(info_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_24
       (.I0(1'b0),
        .O(info_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_3
       (.I0(1'b0),
        .O(self_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_4
       (.I0(1'b0),
        .O(self_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_5
       (.I0(1'b0),
        .O(self_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_6
       (.I0(1'b0),
        .O(self_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_7
       (.I0(1'b0),
        .O(self_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_8
       (.I0(1'b0),
        .O(self_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_9
       (.I0(1'b0),
        .O(info_sf8[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst
       (.I0(self_sf7[7]),
        .O(info_sf7[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__0
       (.I0(self_sf7[6]),
        .O(info_sf7[6]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__1
       (.I0(self_sf7[5]),
        .O(info_sf7[5]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__2
       (.I0(self_sf7[4]),
        .O(info_sf7[4]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__3
       (.I0(self_sf7[3]),
        .O(info_sf7[3]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__4
       (.I0(self_sf7[2]),
        .O(info_sf7[2]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__5
       (.I0(self_sf7[1]),
        .O(info_sf7[1]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__6
       (.I0(self_sf7[0]),
        .O(info_sf7[0]));
endmodule

(* ORIG_REF_NAME = "muxer" *) (* box_type = "black_box" *) (* dont_touch = "true" *) 
module switch_elements_muxer__4
   (enable_i,
    info_o);
  input enable_i;
  output info_o;

  wire enable_i;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf7;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf8;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf9;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [1802:0]self_sf7;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf8;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf9;

  assign info_o = info_sf7[1];
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[0]),
        .S(info_sf7[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1000].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1000]),
        .S(self_sf7[1000]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1001].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1001]),
        .S(self_sf7[1001]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1002].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1002]),
        .S(self_sf7[1002]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1003].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1003]),
        .S(self_sf7[1003]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1004].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1004]),
        .S(self_sf7[1004]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1005].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1005]),
        .S(self_sf7[1005]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1006].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1006]),
        .S(self_sf7[1006]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1007].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1007]),
        .S(self_sf7[1007]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1008].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1008]),
        .S(self_sf7[1008]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1009].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1009]),
        .S(self_sf7[1009]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[100]),
        .S(self_sf7[100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1010].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1010]),
        .S(self_sf7[1010]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1011].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1011]),
        .S(self_sf7[1011]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1012].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1012]),
        .S(self_sf7[1012]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1013].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1013]),
        .S(self_sf7[1013]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1014].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1014]),
        .S(self_sf7[1014]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1015].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1015]),
        .S(self_sf7[1015]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1016].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1016]),
        .S(self_sf7[1016]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1017].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1017]),
        .S(self_sf7[1017]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1018].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1018]),
        .S(self_sf7[1018]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1019].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1019]),
        .S(self_sf7[1019]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[101]),
        .S(self_sf7[101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1020].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1020]),
        .S(self_sf7[1020]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1021].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1021]),
        .S(self_sf7[1021]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1022].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1022]),
        .S(self_sf7[1022]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1023].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1023]),
        .S(self_sf7[1023]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1024].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1024]),
        .S(self_sf7[1024]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1025].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1025]),
        .S(self_sf7[1025]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1026].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1026]),
        .S(self_sf7[1026]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1027].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1027]),
        .S(self_sf7[1027]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1028].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1028]),
        .S(self_sf7[1028]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1029].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1029]),
        .S(self_sf7[1029]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[102]),
        .S(self_sf7[102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1030].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1030]),
        .S(self_sf7[1030]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1031].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1031]),
        .S(self_sf7[1031]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1032].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1032]),
        .S(self_sf7[1032]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1033].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1033]),
        .S(self_sf7[1033]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1034].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1034]),
        .S(self_sf7[1034]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1035].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1035]),
        .S(self_sf7[1035]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1036].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1036]),
        .S(self_sf7[1036]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1037].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1037]),
        .S(self_sf7[1037]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1038].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1038]),
        .S(self_sf7[1038]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1039].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1039]),
        .S(self_sf7[1039]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[103]),
        .S(self_sf7[103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1040].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1040]),
        .S(self_sf7[1040]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1041].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1041]),
        .S(self_sf7[1041]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1042].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1042]),
        .S(self_sf7[1042]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1043].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1043]),
        .S(self_sf7[1043]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1044].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1044]),
        .S(self_sf7[1044]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1045].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1045]),
        .S(self_sf7[1045]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1046].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1046]),
        .S(self_sf7[1046]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1047].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1047]),
        .S(self_sf7[1047]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1048].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1048]),
        .S(self_sf7[1048]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1049].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1049]),
        .S(self_sf7[1049]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[104]),
        .S(self_sf7[104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1050].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1050]),
        .S(self_sf7[1050]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1051].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1051]),
        .S(self_sf7[1051]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1052].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1052]),
        .S(self_sf7[1052]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1053].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1053]),
        .S(self_sf7[1053]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1054].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1054]),
        .S(self_sf7[1054]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1055].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1055]),
        .S(self_sf7[1055]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1056].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1056]),
        .S(self_sf7[1056]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1057].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1057]),
        .S(self_sf7[1057]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1058].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1058]),
        .S(self_sf7[1058]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1059].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1059]),
        .S(self_sf7[1059]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[105]),
        .S(self_sf7[105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1060].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1060]),
        .S(self_sf7[1060]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1061].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1061]),
        .S(self_sf7[1061]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1062].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1062]),
        .S(self_sf7[1062]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1063].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1063]),
        .S(self_sf7[1063]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1064].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1064]),
        .S(self_sf7[1064]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1065].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1065]),
        .S(self_sf7[1065]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1066].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1066]),
        .S(self_sf7[1066]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1067].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1067]),
        .S(self_sf7[1067]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1068].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1068]),
        .S(self_sf7[1068]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1069].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1069]),
        .S(self_sf7[1069]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[106]),
        .S(self_sf7[106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1070].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1070]),
        .S(self_sf7[1070]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1071].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1071]),
        .S(self_sf7[1071]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1072].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1072]),
        .S(self_sf7[1072]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1073].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1073]),
        .S(self_sf7[1073]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1074].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1074]),
        .S(self_sf7[1074]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1075].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1075]),
        .S(self_sf7[1075]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1076].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1076]),
        .S(self_sf7[1076]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1077].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1077]),
        .S(self_sf7[1077]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1078].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1078]),
        .S(self_sf7[1078]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1079].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1079]),
        .S(self_sf7[1079]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[107]),
        .S(self_sf7[107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1080].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1080]),
        .S(self_sf7[1080]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1081].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1081]),
        .S(self_sf7[1081]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1082].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1082]),
        .S(self_sf7[1082]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1083].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1083]),
        .S(self_sf7[1083]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1084].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1084]),
        .S(self_sf7[1084]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1085].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1085]),
        .S(self_sf7[1085]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1086].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1086]),
        .S(self_sf7[1086]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1087].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1087]),
        .S(self_sf7[1087]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1088].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1088]),
        .S(self_sf7[1088]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1089].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1089]),
        .S(self_sf7[1089]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[108]),
        .S(self_sf7[108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1090].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1090]),
        .S(self_sf7[1090]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1091].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1091]),
        .S(self_sf7[1091]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1092].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1092]),
        .S(self_sf7[1092]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1093].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1093]),
        .S(self_sf7[1093]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1094].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1094]),
        .S(self_sf7[1094]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1095].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1095]),
        .S(self_sf7[1095]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1096].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1096]),
        .S(self_sf7[1096]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1097].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1097]),
        .S(self_sf7[1097]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1098].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1098]),
        .S(self_sf7[1098]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1099].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1099]),
        .S(self_sf7[1099]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[109]),
        .S(self_sf7[109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[10].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[10]),
        .S(self_sf7[10]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1100]),
        .S(self_sf7[1100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1101]),
        .S(self_sf7[1101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1102]),
        .S(self_sf7[1102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1103]),
        .S(self_sf7[1103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1104]),
        .S(self_sf7[1104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1105]),
        .S(self_sf7[1105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1106]),
        .S(self_sf7[1106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1107]),
        .S(self_sf7[1107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1108]),
        .S(self_sf7[1108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1109]),
        .S(self_sf7[1109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[110]),
        .S(self_sf7[110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1110]),
        .S(self_sf7[1110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1111]),
        .S(self_sf7[1111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1112]),
        .S(self_sf7[1112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1113]),
        .S(self_sf7[1113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1114]),
        .S(self_sf7[1114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1115]),
        .S(self_sf7[1115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1116]),
        .S(self_sf7[1116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1117]),
        .S(self_sf7[1117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1118]),
        .S(self_sf7[1118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1119]),
        .S(self_sf7[1119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[111]),
        .S(self_sf7[111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1120]),
        .S(self_sf7[1120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1121]),
        .S(self_sf7[1121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1122]),
        .S(self_sf7[1122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1123]),
        .S(self_sf7[1123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1124]),
        .S(self_sf7[1124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1125]),
        .S(self_sf7[1125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1126]),
        .S(self_sf7[1126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1127]),
        .S(self_sf7[1127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1128]),
        .S(self_sf7[1128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1129]),
        .S(self_sf7[1129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[112]),
        .S(self_sf7[112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1130]),
        .S(self_sf7[1130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1131]),
        .S(self_sf7[1131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1132]),
        .S(self_sf7[1132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1133]),
        .S(self_sf7[1133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1134]),
        .S(self_sf7[1134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1135]),
        .S(self_sf7[1135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1136]),
        .S(self_sf7[1136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1137]),
        .S(self_sf7[1137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1138]),
        .S(self_sf7[1138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1139]),
        .S(self_sf7[1139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[113]),
        .S(self_sf7[113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1140]),
        .S(self_sf7[1140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1141]),
        .S(self_sf7[1141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1142]),
        .S(self_sf7[1142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1143]),
        .S(self_sf7[1143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1144]),
        .S(self_sf7[1144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1145]),
        .S(self_sf7[1145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1146]),
        .S(self_sf7[1146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1147]),
        .S(self_sf7[1147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1148]),
        .S(self_sf7[1148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1149]),
        .S(self_sf7[1149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[114]),
        .S(self_sf7[114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1150]),
        .S(self_sf7[1150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1151]),
        .S(self_sf7[1151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1152]),
        .S(self_sf7[1152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1153]),
        .S(self_sf7[1153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1154]),
        .S(self_sf7[1154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1155]),
        .S(self_sf7[1155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1156]),
        .S(self_sf7[1156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1157]),
        .S(self_sf7[1157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1158]),
        .S(self_sf7[1158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1159]),
        .S(self_sf7[1159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[115]),
        .S(self_sf7[115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1160]),
        .S(self_sf7[1160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1161]),
        .S(self_sf7[1161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1162]),
        .S(self_sf7[1162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1163]),
        .S(self_sf7[1163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1164]),
        .S(self_sf7[1164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1165]),
        .S(self_sf7[1165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1166]),
        .S(self_sf7[1166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1167]),
        .S(self_sf7[1167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1168]),
        .S(self_sf7[1168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1169]),
        .S(self_sf7[1169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[116]),
        .S(self_sf7[116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1170]),
        .S(self_sf7[1170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1171]),
        .S(self_sf7[1171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1172]),
        .S(self_sf7[1172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1173]),
        .S(self_sf7[1173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1174]),
        .S(self_sf7[1174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1175]),
        .S(self_sf7[1175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1176]),
        .S(self_sf7[1176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1177]),
        .S(self_sf7[1177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1178]),
        .S(self_sf7[1178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1179]),
        .S(self_sf7[1179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[117]),
        .S(self_sf7[117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1180]),
        .S(self_sf7[1180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1181]),
        .S(self_sf7[1181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1182]),
        .S(self_sf7[1182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1183]),
        .S(self_sf7[1183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1184]),
        .S(self_sf7[1184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1185]),
        .S(self_sf7[1185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1186]),
        .S(self_sf7[1186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1187]),
        .S(self_sf7[1187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1188]),
        .S(self_sf7[1188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1189]),
        .S(self_sf7[1189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[118]),
        .S(self_sf7[118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1190]),
        .S(self_sf7[1190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1191]),
        .S(self_sf7[1191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1192]),
        .S(self_sf7[1192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1193]),
        .S(self_sf7[1193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1194]),
        .S(self_sf7[1194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1195]),
        .S(self_sf7[1195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1196]),
        .S(self_sf7[1196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1197]),
        .S(self_sf7[1197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1198]),
        .S(self_sf7[1198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1199]),
        .S(self_sf7[1199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[119]),
        .S(self_sf7[119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[11].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[11]),
        .S(self_sf7[11]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1200]),
        .S(self_sf7[1200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1201]),
        .S(self_sf7[1201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1202]),
        .S(self_sf7[1202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1203]),
        .S(self_sf7[1203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1204]),
        .S(self_sf7[1204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1205]),
        .S(self_sf7[1205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1206]),
        .S(self_sf7[1206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1207]),
        .S(self_sf7[1207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1208]),
        .S(self_sf7[1208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1209]),
        .S(self_sf7[1209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[120]),
        .S(self_sf7[120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1210]),
        .S(self_sf7[1210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1211]),
        .S(self_sf7[1211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1212]),
        .S(self_sf7[1212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1213]),
        .S(self_sf7[1213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1214]),
        .S(self_sf7[1214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1215]),
        .S(self_sf7[1215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1216]),
        .S(self_sf7[1216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1217]),
        .S(self_sf7[1217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1218]),
        .S(self_sf7[1218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1219]),
        .S(self_sf7[1219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[121]),
        .S(self_sf7[121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1220]),
        .S(self_sf7[1220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1221]),
        .S(self_sf7[1221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1222]),
        .S(self_sf7[1222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1223]),
        .S(self_sf7[1223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1224]),
        .S(self_sf7[1224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1225]),
        .S(self_sf7[1225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1226]),
        .S(self_sf7[1226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1227]),
        .S(self_sf7[1227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1228]),
        .S(self_sf7[1228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1229]),
        .S(self_sf7[1229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[122]),
        .S(self_sf7[122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1230]),
        .S(self_sf7[1230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1231]),
        .S(self_sf7[1231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1232]),
        .S(self_sf7[1232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1233]),
        .S(self_sf7[1233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1234]),
        .S(self_sf7[1234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1235]),
        .S(self_sf7[1235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1236]),
        .S(self_sf7[1236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1237]),
        .S(self_sf7[1237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1238]),
        .S(self_sf7[1238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1239]),
        .S(self_sf7[1239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[123]),
        .S(self_sf7[123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1240]),
        .S(self_sf7[1240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1241]),
        .S(self_sf7[1241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1242]),
        .S(self_sf7[1242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1243]),
        .S(self_sf7[1243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1244]),
        .S(self_sf7[1244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1245]),
        .S(self_sf7[1245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1246]),
        .S(self_sf7[1246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1247]),
        .S(self_sf7[1247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1248]),
        .S(self_sf7[1248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1249]),
        .S(self_sf7[1249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[124]),
        .S(self_sf7[124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1250]),
        .S(self_sf7[1250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1251]),
        .S(self_sf7[1251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1252]),
        .S(self_sf7[1252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1253]),
        .S(self_sf7[1253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1254]),
        .S(self_sf7[1254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1255]),
        .S(self_sf7[1255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1256]),
        .S(self_sf7[1256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1257]),
        .S(self_sf7[1257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1258]),
        .S(self_sf7[1258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1259]),
        .S(self_sf7[1259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[125]),
        .S(self_sf7[125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1260]),
        .S(self_sf7[1260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1261]),
        .S(self_sf7[1261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1262]),
        .S(self_sf7[1262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1263]),
        .S(self_sf7[1263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1264]),
        .S(self_sf7[1264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1265]),
        .S(self_sf7[1265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1266]),
        .S(self_sf7[1266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1267]),
        .S(self_sf7[1267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1268]),
        .S(self_sf7[1268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1269]),
        .S(self_sf7[1269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[126]),
        .S(self_sf7[126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1270]),
        .S(self_sf7[1270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1271]),
        .S(self_sf7[1271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1272]),
        .S(self_sf7[1272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1273]),
        .S(self_sf7[1273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1274]),
        .S(self_sf7[1274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1275]),
        .S(self_sf7[1275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1276]),
        .S(self_sf7[1276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1277]),
        .S(self_sf7[1277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1278]),
        .S(self_sf7[1278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1279]),
        .S(self_sf7[1279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[127]),
        .S(self_sf7[127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1280]),
        .S(self_sf7[1280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1281]),
        .S(self_sf7[1281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1282]),
        .S(self_sf7[1282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1283]),
        .S(self_sf7[1283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1284]),
        .S(self_sf7[1284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1285]),
        .S(self_sf7[1285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1286]),
        .S(self_sf7[1286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1287]),
        .S(self_sf7[1287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1288]),
        .S(self_sf7[1288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1289]),
        .S(self_sf7[1289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[128]),
        .S(self_sf7[128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1290]),
        .S(self_sf7[1290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1291]),
        .S(self_sf7[1291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1292]),
        .S(self_sf7[1292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1293]),
        .S(self_sf7[1293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1294]),
        .S(self_sf7[1294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1295]),
        .S(self_sf7[1295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1296]),
        .S(self_sf7[1296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1297]),
        .S(self_sf7[1297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1298]),
        .S(self_sf7[1298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1299]),
        .S(self_sf7[1299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[129]),
        .S(self_sf7[129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[12].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[12]),
        .S(self_sf7[12]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1300]),
        .S(self_sf7[1300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1301]),
        .S(self_sf7[1301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1302]),
        .S(self_sf7[1302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1303]),
        .S(self_sf7[1303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1304]),
        .S(self_sf7[1304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1305]),
        .S(self_sf7[1305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1306]),
        .S(self_sf7[1306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1307]),
        .S(self_sf7[1307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1308]),
        .S(self_sf7[1308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1309]),
        .S(self_sf7[1309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[130]),
        .S(self_sf7[130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1310]),
        .S(self_sf7[1310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1311]),
        .S(self_sf7[1311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1312]),
        .S(self_sf7[1312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1313]),
        .S(self_sf7[1313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1314]),
        .S(self_sf7[1314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1315]),
        .S(self_sf7[1315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1316]),
        .S(self_sf7[1316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1317]),
        .S(self_sf7[1317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1318]),
        .S(self_sf7[1318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1319]),
        .S(self_sf7[1319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[131]),
        .S(self_sf7[131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1320]),
        .S(self_sf7[1320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1321]),
        .S(self_sf7[1321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1322]),
        .S(self_sf7[1322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1323]),
        .S(self_sf7[1323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1324]),
        .S(self_sf7[1324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1325]),
        .S(self_sf7[1325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1326]),
        .S(self_sf7[1326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1327]),
        .S(self_sf7[1327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1328]),
        .S(self_sf7[1328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1329]),
        .S(self_sf7[1329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[132]),
        .S(self_sf7[132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1330]),
        .S(self_sf7[1330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1331]),
        .S(self_sf7[1331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1332]),
        .S(self_sf7[1332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1333]),
        .S(self_sf7[1333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1334]),
        .S(self_sf7[1334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1335]),
        .S(self_sf7[1335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1336]),
        .S(self_sf7[1336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1337]),
        .S(self_sf7[1337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1338]),
        .S(self_sf7[1338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1339]),
        .S(self_sf7[1339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[133]),
        .S(self_sf7[133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1340]),
        .S(self_sf7[1340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1341]),
        .S(self_sf7[1341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1342]),
        .S(self_sf7[1342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1343]),
        .S(self_sf7[1343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1344]),
        .S(self_sf7[1344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1345]),
        .S(self_sf7[1345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1346]),
        .S(self_sf7[1346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1347]),
        .S(self_sf7[1347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1348]),
        .S(self_sf7[1348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1349]),
        .S(self_sf7[1349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[134]),
        .S(self_sf7[134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1350]),
        .S(self_sf7[1350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1351]),
        .S(self_sf7[1351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1352]),
        .S(self_sf7[1352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1353]),
        .S(self_sf7[1353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1354]),
        .S(self_sf7[1354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1355]),
        .S(self_sf7[1355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1356]),
        .S(self_sf7[1356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1357]),
        .S(self_sf7[1357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1358]),
        .S(self_sf7[1358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1359]),
        .S(self_sf7[1359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[135]),
        .S(self_sf7[135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1360]),
        .S(self_sf7[1360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1361]),
        .S(self_sf7[1361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1362]),
        .S(self_sf7[1362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1363]),
        .S(self_sf7[1363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1364]),
        .S(self_sf7[1364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1365]),
        .S(self_sf7[1365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1366]),
        .S(self_sf7[1366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1367]),
        .S(self_sf7[1367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1368]),
        .S(self_sf7[1368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1369]),
        .S(self_sf7[1369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[136]),
        .S(self_sf7[136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1370]),
        .S(self_sf7[1370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1371]),
        .S(self_sf7[1371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1372]),
        .S(self_sf7[1372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1373]),
        .S(self_sf7[1373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1374]),
        .S(self_sf7[1374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1375]),
        .S(self_sf7[1375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1376]),
        .S(self_sf7[1376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1377]),
        .S(self_sf7[1377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1378]),
        .S(self_sf7[1378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1379]),
        .S(self_sf7[1379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[137]),
        .S(self_sf7[137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1380]),
        .S(self_sf7[1380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1381]),
        .S(self_sf7[1381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1382]),
        .S(self_sf7[1382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1383]),
        .S(self_sf7[1383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1384]),
        .S(self_sf7[1384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1385]),
        .S(self_sf7[1385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1386]),
        .S(self_sf7[1386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1387]),
        .S(self_sf7[1387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1388]),
        .S(self_sf7[1388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1389]),
        .S(self_sf7[1389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[138]),
        .S(self_sf7[138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1390]),
        .S(self_sf7[1390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1391]),
        .S(self_sf7[1391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1392]),
        .S(self_sf7[1392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1393]),
        .S(self_sf7[1393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1394]),
        .S(self_sf7[1394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1395]),
        .S(self_sf7[1395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1396]),
        .S(self_sf7[1396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1397]),
        .S(self_sf7[1397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1398]),
        .S(self_sf7[1398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1399]),
        .S(self_sf7[1399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[139]),
        .S(self_sf7[139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[13].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[13]),
        .S(self_sf7[13]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1400]),
        .S(self_sf7[1400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1401]),
        .S(self_sf7[1401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1402]),
        .S(self_sf7[1402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1403]),
        .S(self_sf7[1403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1404]),
        .S(self_sf7[1404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1405]),
        .S(self_sf7[1405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1406]),
        .S(self_sf7[1406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1407]),
        .S(self_sf7[1407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1408]),
        .S(self_sf7[1408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1409]),
        .S(self_sf7[1409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[140]),
        .S(self_sf7[140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1410]),
        .S(self_sf7[1410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1411]),
        .S(self_sf7[1411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1412]),
        .S(self_sf7[1412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1413]),
        .S(self_sf7[1413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1414]),
        .S(self_sf7[1414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1415]),
        .S(self_sf7[1415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1416]),
        .S(self_sf7[1416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1417]),
        .S(self_sf7[1417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1418]),
        .S(self_sf7[1418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1419]),
        .S(self_sf7[1419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[141]),
        .S(self_sf7[141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1420]),
        .S(self_sf7[1420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1421]),
        .S(self_sf7[1421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1422]),
        .S(self_sf7[1422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1423]),
        .S(self_sf7[1423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1424]),
        .S(self_sf7[1424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1425]),
        .S(self_sf7[1425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1426]),
        .S(self_sf7[1426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1427]),
        .S(self_sf7[1427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1428]),
        .S(self_sf7[1428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1429]),
        .S(self_sf7[1429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[142]),
        .S(self_sf7[142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1430]),
        .S(self_sf7[1430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1431]),
        .S(self_sf7[1431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1432]),
        .S(self_sf7[1432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1433]),
        .S(self_sf7[1433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1434]),
        .S(self_sf7[1434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1435]),
        .S(self_sf7[1435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1436]),
        .S(self_sf7[1436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1437]),
        .S(self_sf7[1437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1438]),
        .S(self_sf7[1438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1439]),
        .S(self_sf7[1439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[143]),
        .S(self_sf7[143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1440]),
        .S(self_sf7[1440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1441]),
        .S(self_sf7[1441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1442]),
        .S(self_sf7[1442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1443]),
        .S(self_sf7[1443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1444]),
        .S(self_sf7[1444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1445]),
        .S(self_sf7[1445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1446]),
        .S(self_sf7[1446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1447]),
        .S(self_sf7[1447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1448]),
        .S(self_sf7[1448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1449]),
        .S(self_sf7[1449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[144]),
        .S(self_sf7[144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1450]),
        .S(self_sf7[1450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1451]),
        .S(self_sf7[1451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1452]),
        .S(self_sf7[1452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1453]),
        .S(self_sf7[1453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1454]),
        .S(self_sf7[1454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1455]),
        .S(self_sf7[1455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1456]),
        .S(self_sf7[1456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1457]),
        .S(self_sf7[1457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1458]),
        .S(self_sf7[1458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1459]),
        .S(self_sf7[1459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[145]),
        .S(self_sf7[145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1460]),
        .S(self_sf7[1460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1461]),
        .S(self_sf7[1461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1462]),
        .S(self_sf7[1462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1463]),
        .S(self_sf7[1463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1464]),
        .S(self_sf7[1464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1465]),
        .S(self_sf7[1465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1466]),
        .S(self_sf7[1466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1467]),
        .S(self_sf7[1467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1468]),
        .S(self_sf7[1468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1469]),
        .S(self_sf7[1469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[146]),
        .S(self_sf7[146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1470]),
        .S(self_sf7[1470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1471]),
        .S(self_sf7[1471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1472]),
        .S(self_sf7[1472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1473]),
        .S(self_sf7[1473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1474]),
        .S(self_sf7[1474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1475]),
        .S(self_sf7[1475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1476]),
        .S(self_sf7[1476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1477]),
        .S(self_sf7[1477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1478]),
        .S(self_sf7[1478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1479]),
        .S(self_sf7[1479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[147]),
        .S(self_sf7[147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1480]),
        .S(self_sf7[1480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1481]),
        .S(self_sf7[1481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1482]),
        .S(self_sf7[1482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1483]),
        .S(self_sf7[1483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1484]),
        .S(self_sf7[1484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1485]),
        .S(self_sf7[1485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1486]),
        .S(self_sf7[1486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1487]),
        .S(self_sf7[1487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1488]),
        .S(self_sf7[1488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1489]),
        .S(self_sf7[1489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[148]),
        .S(self_sf7[148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1490]),
        .S(self_sf7[1490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1491]),
        .S(self_sf7[1491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1492]),
        .S(self_sf7[1492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1493]),
        .S(self_sf7[1493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1494]),
        .S(self_sf7[1494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1495]),
        .S(self_sf7[1495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1496]),
        .S(self_sf7[1496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1497]),
        .S(self_sf7[1497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1498]),
        .S(self_sf7[1498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1499]),
        .S(self_sf7[1499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[149]),
        .S(self_sf7[149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[14].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[14]),
        .S(self_sf7[14]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1500]),
        .S(self_sf7[1500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1501]),
        .S(self_sf7[1501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1502]),
        .S(self_sf7[1502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1503]),
        .S(self_sf7[1503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1504]),
        .S(self_sf7[1504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1505]),
        .S(self_sf7[1505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1506]),
        .S(self_sf7[1506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1507]),
        .S(self_sf7[1507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1508]),
        .S(self_sf7[1508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1509]),
        .S(self_sf7[1509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[150]),
        .S(self_sf7[150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1510]),
        .S(self_sf7[1510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1511]),
        .S(self_sf7[1511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1512]),
        .S(self_sf7[1512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1513]),
        .S(self_sf7[1513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1514]),
        .S(self_sf7[1514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1515]),
        .S(self_sf7[1515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1516]),
        .S(self_sf7[1516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1517]),
        .S(self_sf7[1517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1518]),
        .S(self_sf7[1518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1519]),
        .S(self_sf7[1519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[151]),
        .S(self_sf7[151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1520]),
        .S(self_sf7[1520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1521]),
        .S(self_sf7[1521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1522]),
        .S(self_sf7[1522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1523]),
        .S(self_sf7[1523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1524]),
        .S(self_sf7[1524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1525]),
        .S(self_sf7[1525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1526]),
        .S(self_sf7[1526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1527]),
        .S(self_sf7[1527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1528]),
        .S(self_sf7[1528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1529]),
        .S(self_sf7[1529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[152]),
        .S(self_sf7[152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1530]),
        .S(self_sf7[1530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1531]),
        .S(self_sf7[1531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1532]),
        .S(self_sf7[1532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1533]),
        .S(self_sf7[1533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1534]),
        .S(self_sf7[1534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1535]),
        .S(self_sf7[1535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1536]),
        .S(self_sf7[1536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1537]),
        .S(self_sf7[1537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1538]),
        .S(self_sf7[1538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1539]),
        .S(self_sf7[1539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[153]),
        .S(self_sf7[153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1540]),
        .S(self_sf7[1540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1541]),
        .S(self_sf7[1541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1542]),
        .S(self_sf7[1542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1543]),
        .S(self_sf7[1543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1544]),
        .S(self_sf7[1544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1545]),
        .S(self_sf7[1545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1546]),
        .S(self_sf7[1546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1547]),
        .S(self_sf7[1547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1548]),
        .S(self_sf7[1548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1549]),
        .S(self_sf7[1549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[154]),
        .S(self_sf7[154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1550]),
        .S(self_sf7[1550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1551]),
        .S(self_sf7[1551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1552]),
        .S(self_sf7[1552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1553]),
        .S(self_sf7[1553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1554]),
        .S(self_sf7[1554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1555]),
        .S(self_sf7[1555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1556]),
        .S(self_sf7[1556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1557]),
        .S(self_sf7[1557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1558]),
        .S(self_sf7[1558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1559]),
        .S(self_sf7[1559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[155]),
        .S(self_sf7[155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1560]),
        .S(self_sf7[1560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1561]),
        .S(self_sf7[1561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1562]),
        .S(self_sf7[1562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1563]),
        .S(self_sf7[1563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1564]),
        .S(self_sf7[1564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1565]),
        .S(self_sf7[1565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1566]),
        .S(self_sf7[1566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1567]),
        .S(self_sf7[1567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1568]),
        .S(self_sf7[1568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1569]),
        .S(self_sf7[1569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[156]),
        .S(self_sf7[156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1570]),
        .S(self_sf7[1570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1571]),
        .S(self_sf7[1571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1572]),
        .S(self_sf7[1572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1573]),
        .S(self_sf7[1573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1574]),
        .S(self_sf7[1574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1575]),
        .S(self_sf7[1575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1576]),
        .S(self_sf7[1576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1577]),
        .S(self_sf7[1577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1578]),
        .S(self_sf7[1578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1579]),
        .S(self_sf7[1579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[157]),
        .S(self_sf7[157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1580]),
        .S(self_sf7[1580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1581]),
        .S(self_sf7[1581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1582]),
        .S(self_sf7[1582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1583]),
        .S(self_sf7[1583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1584]),
        .S(self_sf7[1584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1585]),
        .S(self_sf7[1585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1586]),
        .S(self_sf7[1586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1587]),
        .S(self_sf7[1587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1588]),
        .S(self_sf7[1588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1589]),
        .S(self_sf7[1589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[158]),
        .S(self_sf7[158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1590]),
        .S(self_sf7[1590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1591]),
        .S(self_sf7[1591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1592]),
        .S(self_sf7[1592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1593]),
        .S(self_sf7[1593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1594]),
        .S(self_sf7[1594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1595]),
        .S(self_sf7[1595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1596]),
        .S(self_sf7[1596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1597]),
        .S(self_sf7[1597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1598]),
        .S(self_sf7[1598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1599]),
        .S(self_sf7[1599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[159]),
        .S(self_sf7[159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[15].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[15]),
        .S(self_sf7[15]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1600]),
        .S(self_sf7[1600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1601]),
        .S(self_sf7[1601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1602]),
        .S(self_sf7[1602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1603]),
        .S(self_sf7[1603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1604]),
        .S(self_sf7[1604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1605]),
        .S(self_sf7[1605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1606]),
        .S(self_sf7[1606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1607]),
        .S(self_sf7[1607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1608]),
        .S(self_sf7[1608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1609]),
        .S(self_sf7[1609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[160]),
        .S(self_sf7[160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1610]),
        .S(self_sf7[1610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1611]),
        .S(self_sf7[1611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1612]),
        .S(self_sf7[1612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1613]),
        .S(self_sf7[1613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1614]),
        .S(self_sf7[1614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1615]),
        .S(self_sf7[1615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1616]),
        .S(self_sf7[1616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1617]),
        .S(self_sf7[1617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1618]),
        .S(self_sf7[1618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1619]),
        .S(self_sf7[1619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[161]),
        .S(self_sf7[161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1620]),
        .S(self_sf7[1620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1621]),
        .S(self_sf7[1621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1622]),
        .S(self_sf7[1622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1623]),
        .S(self_sf7[1623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1624]),
        .S(self_sf7[1624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1625]),
        .S(self_sf7[1625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1626]),
        .S(self_sf7[1626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1627]),
        .S(self_sf7[1627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1628]),
        .S(self_sf7[1628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1629]),
        .S(self_sf7[1629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[162]),
        .S(self_sf7[162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1630]),
        .S(self_sf7[1630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1631]),
        .S(self_sf7[1631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1632]),
        .S(self_sf7[1632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1633]),
        .S(self_sf7[1633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1634]),
        .S(self_sf7[1634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1635]),
        .S(self_sf7[1635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1636]),
        .S(self_sf7[1636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1637]),
        .S(self_sf7[1637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1638]),
        .S(self_sf7[1638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1639]),
        .S(self_sf7[1639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[163]),
        .S(self_sf7[163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1640]),
        .S(self_sf7[1640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1641]),
        .S(self_sf7[1641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1642]),
        .S(self_sf7[1642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1643]),
        .S(self_sf7[1643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1644]),
        .S(self_sf7[1644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1645]),
        .S(self_sf7[1645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1646]),
        .S(self_sf7[1646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1647]),
        .S(self_sf7[1647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1648]),
        .S(self_sf7[1648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1649]),
        .S(self_sf7[1649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[164]),
        .S(self_sf7[164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1650]),
        .S(self_sf7[1650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1651]),
        .S(self_sf7[1651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1652]),
        .S(self_sf7[1652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1653]),
        .S(self_sf7[1653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1654]),
        .S(self_sf7[1654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1655]),
        .S(self_sf7[1655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1656]),
        .S(self_sf7[1656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1657]),
        .S(self_sf7[1657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1658]),
        .S(self_sf7[1658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1659]),
        .S(self_sf7[1659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[165]),
        .S(self_sf7[165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1660]),
        .S(self_sf7[1660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1661]),
        .S(self_sf7[1661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1662]),
        .S(self_sf7[1662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1663]),
        .S(self_sf7[1663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1664]),
        .S(self_sf7[1664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1665]),
        .S(self_sf7[1665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1666]),
        .S(self_sf7[1666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1667]),
        .S(self_sf7[1667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1668]),
        .S(self_sf7[1668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1669]),
        .S(self_sf7[1669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[166]),
        .S(self_sf7[166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1670]),
        .S(self_sf7[1670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1671]),
        .S(self_sf7[1671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1672]),
        .S(self_sf7[1672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1673]),
        .S(self_sf7[1673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1674]),
        .S(self_sf7[1674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1675]),
        .S(self_sf7[1675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1676]),
        .S(self_sf7[1676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1677]),
        .S(self_sf7[1677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1678]),
        .S(self_sf7[1678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1679]),
        .S(self_sf7[1679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[167]),
        .S(self_sf7[167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1680]),
        .S(self_sf7[1680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1681]),
        .S(self_sf7[1681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1682]),
        .S(self_sf7[1682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1683]),
        .S(self_sf7[1683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1684]),
        .S(self_sf7[1684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1685]),
        .S(self_sf7[1685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1686]),
        .S(self_sf7[1686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1687]),
        .S(self_sf7[1687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1688]),
        .S(self_sf7[1688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1689]),
        .S(self_sf7[1689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[168]),
        .S(self_sf7[168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1690]),
        .S(self_sf7[1690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1691]),
        .S(self_sf7[1691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1692]),
        .S(self_sf7[1692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1693]),
        .S(self_sf7[1693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1694]),
        .S(self_sf7[1694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1695]),
        .S(self_sf7[1695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1696]),
        .S(self_sf7[1696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1697]),
        .S(self_sf7[1697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1698]),
        .S(self_sf7[1698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1699]),
        .S(self_sf7[1699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[169]),
        .S(self_sf7[169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[16].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[16]),
        .S(self_sf7[16]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1700]),
        .S(self_sf7[1700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1701]),
        .S(self_sf7[1701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1702]),
        .S(self_sf7[1702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1703]),
        .S(self_sf7[1703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1704]),
        .S(self_sf7[1704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1705]),
        .S(self_sf7[1705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1706]),
        .S(self_sf7[1706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1707]),
        .S(self_sf7[1707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1708]),
        .S(self_sf7[1708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1709]),
        .S(self_sf7[1709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[170]),
        .S(self_sf7[170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1710]),
        .S(self_sf7[1710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1711]),
        .S(self_sf7[1711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1712]),
        .S(self_sf7[1712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1713]),
        .S(self_sf7[1713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1714]),
        .S(self_sf7[1714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1715]),
        .S(self_sf7[1715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1716]),
        .S(self_sf7[1716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1717]),
        .S(self_sf7[1717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1718]),
        .S(self_sf7[1718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1719]),
        .S(self_sf7[1719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[171]),
        .S(self_sf7[171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1720]),
        .S(self_sf7[1720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1721]),
        .S(self_sf7[1721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1722]),
        .S(self_sf7[1722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1723]),
        .S(self_sf7[1723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1724]),
        .S(self_sf7[1724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1725]),
        .S(self_sf7[1725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1726]),
        .S(self_sf7[1726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1727]),
        .S(self_sf7[1727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1728]),
        .S(self_sf7[1728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1729]),
        .S(self_sf7[1729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[172]),
        .S(self_sf7[172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1730]),
        .S(self_sf7[1730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1731]),
        .S(self_sf7[1731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1732]),
        .S(self_sf7[1732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1733]),
        .S(self_sf7[1733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1734]),
        .S(self_sf7[1734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1735]),
        .S(self_sf7[1735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1736]),
        .S(self_sf7[1736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1737]),
        .S(self_sf7[1737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1738]),
        .S(self_sf7[1738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1739]),
        .S(self_sf7[1739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[173]),
        .S(self_sf7[173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1740]),
        .S(self_sf7[1740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1741]),
        .S(self_sf7[1741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1742]),
        .S(self_sf7[1742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1743]),
        .S(self_sf7[1743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1744]),
        .S(self_sf7[1744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1745]),
        .S(self_sf7[1745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1746]),
        .S(self_sf7[1746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1747]),
        .S(self_sf7[1747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1748]),
        .S(self_sf7[1748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1749]),
        .S(self_sf7[1749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[174]),
        .S(self_sf7[174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1750]),
        .S(self_sf7[1750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1751]),
        .S(self_sf7[1751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1752]),
        .S(self_sf7[1752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1753]),
        .S(self_sf7[1753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1754]),
        .S(self_sf7[1754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1755]),
        .S(self_sf7[1755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1756]),
        .S(self_sf7[1756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1757]),
        .S(self_sf7[1757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1758]),
        .S(self_sf7[1758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1759]),
        .S(self_sf7[1759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[175]),
        .S(self_sf7[175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1760]),
        .S(self_sf7[1760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1761]),
        .S(self_sf7[1761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1762]),
        .S(self_sf7[1762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1763]),
        .S(self_sf7[1763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1764]),
        .S(self_sf7[1764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1765]),
        .S(self_sf7[1765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1766]),
        .S(self_sf7[1766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1767]),
        .S(self_sf7[1767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1768]),
        .S(self_sf7[1768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1769]),
        .S(self_sf7[1769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[176]),
        .S(self_sf7[176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1770]),
        .S(self_sf7[1770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1771]),
        .S(self_sf7[1771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1772]),
        .S(self_sf7[1772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1773]),
        .S(self_sf7[1773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1774]),
        .S(self_sf7[1774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1775]),
        .S(self_sf7[1775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1776]),
        .S(self_sf7[1776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1777]),
        .S(self_sf7[1777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1778]),
        .S(self_sf7[1778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1779]),
        .S(self_sf7[1779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[177]),
        .S(self_sf7[177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1780]),
        .S(self_sf7[1780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1781]),
        .S(self_sf7[1781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1782]),
        .S(self_sf7[1782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1783]),
        .S(self_sf7[1783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1784]),
        .S(self_sf7[1784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1785]),
        .S(self_sf7[1785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1786]),
        .S(self_sf7[1786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1787]),
        .S(self_sf7[1787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1788]),
        .S(self_sf7[1788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1789]),
        .S(self_sf7[1789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[178]),
        .S(self_sf7[178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1790]),
        .S(self_sf7[1790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1791]),
        .S(self_sf7[1791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1792]),
        .S(self_sf7[1792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1793]),
        .S(self_sf7[1793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1794]),
        .S(self_sf7[1794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1795]),
        .S(self_sf7[1795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1796]),
        .S(self_sf7[1796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1797]),
        .S(self_sf7[1797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1798]),
        .S(self_sf7[1798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1799]),
        .S(self_sf7[1799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[179]),
        .S(self_sf7[179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[17].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[17]),
        .S(self_sf7[17]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[180]),
        .S(self_sf7[180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[181]),
        .S(self_sf7[181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[182]),
        .S(self_sf7[182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[183]),
        .S(self_sf7[183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[184]),
        .S(self_sf7[184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[185]),
        .S(self_sf7[185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[186]),
        .S(self_sf7[186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[187]),
        .S(self_sf7[187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[188]),
        .S(self_sf7[188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[189]),
        .S(self_sf7[189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[18].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[18]),
        .S(self_sf7[18]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[190]),
        .S(self_sf7[190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[191]),
        .S(self_sf7[191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[192]),
        .S(self_sf7[192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[193]),
        .S(self_sf7[193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[194]),
        .S(self_sf7[194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[195]),
        .S(self_sf7[195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[196]),
        .S(self_sf7[196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[197]),
        .S(self_sf7[197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[198]),
        .S(self_sf7[198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[199]),
        .S(self_sf7[199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[19].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[19]),
        .S(self_sf7[19]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1]),
        .S(info_sf7[1]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[200]),
        .S(self_sf7[200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[201]),
        .S(self_sf7[201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[202]),
        .S(self_sf7[202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[203]),
        .S(self_sf7[203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[204]),
        .S(self_sf7[204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[205]),
        .S(self_sf7[205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[206]),
        .S(self_sf7[206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[207]),
        .S(self_sf7[207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[208]),
        .S(self_sf7[208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[209]),
        .S(self_sf7[209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[20].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[20]),
        .S(self_sf7[20]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[210]),
        .S(self_sf7[210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[211]),
        .S(self_sf7[211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[212]),
        .S(self_sf7[212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[213]),
        .S(self_sf7[213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[214]),
        .S(self_sf7[214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[215]),
        .S(self_sf7[215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[216]),
        .S(self_sf7[216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[217]),
        .S(self_sf7[217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[218]),
        .S(self_sf7[218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[219]),
        .S(self_sf7[219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[21].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[21]),
        .S(self_sf7[21]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[220]),
        .S(self_sf7[220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[221]),
        .S(self_sf7[221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[222]),
        .S(self_sf7[222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[223]),
        .S(self_sf7[223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[224]),
        .S(self_sf7[224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[225]),
        .S(self_sf7[225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[226]),
        .S(self_sf7[226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[227]),
        .S(self_sf7[227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[228]),
        .S(self_sf7[228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[229]),
        .S(self_sf7[229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[22].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[22]),
        .S(self_sf7[22]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[230]),
        .S(self_sf7[230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[231]),
        .S(self_sf7[231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[232]),
        .S(self_sf7[232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[233]),
        .S(self_sf7[233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[234]),
        .S(self_sf7[234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[235]),
        .S(self_sf7[235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[236]),
        .S(self_sf7[236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[237]),
        .S(self_sf7[237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[238]),
        .S(self_sf7[238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[239]),
        .S(self_sf7[239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[23].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[23]),
        .S(self_sf7[23]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[240]),
        .S(self_sf7[240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[241]),
        .S(self_sf7[241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[242]),
        .S(self_sf7[242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[243]),
        .S(self_sf7[243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[244]),
        .S(self_sf7[244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[245]),
        .S(self_sf7[245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[246]),
        .S(self_sf7[246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[247]),
        .S(self_sf7[247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[248]),
        .S(self_sf7[248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[249]),
        .S(self_sf7[249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[24].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[24]),
        .S(self_sf7[24]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[250]),
        .S(self_sf7[250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[251]),
        .S(self_sf7[251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[252]),
        .S(self_sf7[252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[253]),
        .S(self_sf7[253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[254]),
        .S(self_sf7[254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[255]),
        .S(self_sf7[255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[256]),
        .S(self_sf7[256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[257]),
        .S(self_sf7[257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[258]),
        .S(self_sf7[258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[259]),
        .S(self_sf7[259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[25].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[25]),
        .S(self_sf7[25]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[260]),
        .S(self_sf7[260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[261]),
        .S(self_sf7[261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[262]),
        .S(self_sf7[262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[263]),
        .S(self_sf7[263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[264]),
        .S(self_sf7[264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[265]),
        .S(self_sf7[265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[266]),
        .S(self_sf7[266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[267]),
        .S(self_sf7[267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[268]),
        .S(self_sf7[268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[269]),
        .S(self_sf7[269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[26].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[26]),
        .S(self_sf7[26]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[270]),
        .S(self_sf7[270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[271]),
        .S(self_sf7[271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[272]),
        .S(self_sf7[272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[273]),
        .S(self_sf7[273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[274]),
        .S(self_sf7[274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[275]),
        .S(self_sf7[275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[276]),
        .S(self_sf7[276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[277]),
        .S(self_sf7[277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[278]),
        .S(self_sf7[278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[279]),
        .S(self_sf7[279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[27].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[27]),
        .S(self_sf7[27]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[280]),
        .S(self_sf7[280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[281]),
        .S(self_sf7[281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[282]),
        .S(self_sf7[282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[283]),
        .S(self_sf7[283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[284]),
        .S(self_sf7[284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[285]),
        .S(self_sf7[285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[286]),
        .S(self_sf7[286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[287]),
        .S(self_sf7[287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[288]),
        .S(self_sf7[288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[289]),
        .S(self_sf7[289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[28].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[28]),
        .S(self_sf7[28]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[290]),
        .S(self_sf7[290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[291]),
        .S(self_sf7[291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[292]),
        .S(self_sf7[292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[293]),
        .S(self_sf7[293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[294]),
        .S(self_sf7[294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[295]),
        .S(self_sf7[295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[296]),
        .S(self_sf7[296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[297]),
        .S(self_sf7[297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[298]),
        .S(self_sf7[298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[299]),
        .S(self_sf7[299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[29].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[29]),
        .S(self_sf7[29]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[2].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[2]),
        .S(info_sf7[2]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[300]),
        .S(self_sf7[300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[301]),
        .S(self_sf7[301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[302]),
        .S(self_sf7[302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[303]),
        .S(self_sf7[303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[304]),
        .S(self_sf7[304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[305]),
        .S(self_sf7[305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[306]),
        .S(self_sf7[306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[307]),
        .S(self_sf7[307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[308]),
        .S(self_sf7[308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[309]),
        .S(self_sf7[309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[30].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[30]),
        .S(self_sf7[30]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[310]),
        .S(self_sf7[310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[311]),
        .S(self_sf7[311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[312]),
        .S(self_sf7[312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[313]),
        .S(self_sf7[313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[314]),
        .S(self_sf7[314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[315]),
        .S(self_sf7[315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[316]),
        .S(self_sf7[316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[317]),
        .S(self_sf7[317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[318]),
        .S(self_sf7[318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[319]),
        .S(self_sf7[319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[31].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[31]),
        .S(self_sf7[31]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[320]),
        .S(self_sf7[320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[321]),
        .S(self_sf7[321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[322]),
        .S(self_sf7[322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[323]),
        .S(self_sf7[323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[324]),
        .S(self_sf7[324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[325]),
        .S(self_sf7[325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[326]),
        .S(self_sf7[326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[327]),
        .S(self_sf7[327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[328]),
        .S(self_sf7[328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[329]),
        .S(self_sf7[329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[32].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[32]),
        .S(self_sf7[32]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[330]),
        .S(self_sf7[330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[331]),
        .S(self_sf7[331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[332]),
        .S(self_sf7[332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[333]),
        .S(self_sf7[333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[334]),
        .S(self_sf7[334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[335]),
        .S(self_sf7[335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[336]),
        .S(self_sf7[336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[337]),
        .S(self_sf7[337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[338]),
        .S(self_sf7[338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[339]),
        .S(self_sf7[339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[33].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[33]),
        .S(self_sf7[33]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[340]),
        .S(self_sf7[340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[341]),
        .S(self_sf7[341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[342]),
        .S(self_sf7[342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[343]),
        .S(self_sf7[343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[344]),
        .S(self_sf7[344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[345]),
        .S(self_sf7[345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[346]),
        .S(self_sf7[346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[347]),
        .S(self_sf7[347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[348]),
        .S(self_sf7[348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[349]),
        .S(self_sf7[349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[34].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[34]),
        .S(self_sf7[34]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[350]),
        .S(self_sf7[350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[351]),
        .S(self_sf7[351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[352]),
        .S(self_sf7[352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[353]),
        .S(self_sf7[353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[354]),
        .S(self_sf7[354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[355]),
        .S(self_sf7[355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[356]),
        .S(self_sf7[356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[357]),
        .S(self_sf7[357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[358]),
        .S(self_sf7[358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[359]),
        .S(self_sf7[359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[35].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[35]),
        .S(self_sf7[35]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[360]),
        .S(self_sf7[360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[361]),
        .S(self_sf7[361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[362]),
        .S(self_sf7[362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[363]),
        .S(self_sf7[363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[364]),
        .S(self_sf7[364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[365]),
        .S(self_sf7[365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[366]),
        .S(self_sf7[366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[367]),
        .S(self_sf7[367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[368]),
        .S(self_sf7[368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[369]),
        .S(self_sf7[369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[36].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[36]),
        .S(self_sf7[36]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[370]),
        .S(self_sf7[370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[371]),
        .S(self_sf7[371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[372]),
        .S(self_sf7[372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[373]),
        .S(self_sf7[373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[374]),
        .S(self_sf7[374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[375]),
        .S(self_sf7[375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[376]),
        .S(self_sf7[376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[377]),
        .S(self_sf7[377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[378]),
        .S(self_sf7[378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[379]),
        .S(self_sf7[379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[37].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[37]),
        .S(self_sf7[37]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[380]),
        .S(self_sf7[380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[381]),
        .S(self_sf7[381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[382]),
        .S(self_sf7[382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[383]),
        .S(self_sf7[383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[384]),
        .S(self_sf7[384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[385]),
        .S(self_sf7[385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[386]),
        .S(self_sf7[386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[387]),
        .S(self_sf7[387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[388]),
        .S(self_sf7[388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[389]),
        .S(self_sf7[389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[38].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[38]),
        .S(self_sf7[38]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[390]),
        .S(self_sf7[390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[391]),
        .S(self_sf7[391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[392]),
        .S(self_sf7[392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[393]),
        .S(self_sf7[393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[394]),
        .S(self_sf7[394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[395]),
        .S(self_sf7[395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[396]),
        .S(self_sf7[396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[397]),
        .S(self_sf7[397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[398]),
        .S(self_sf7[398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[399]),
        .S(self_sf7[399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[39].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[39]),
        .S(self_sf7[39]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[3].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[3]),
        .S(info_sf7[3]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[400]),
        .S(self_sf7[400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[401]),
        .S(self_sf7[401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[402]),
        .S(self_sf7[402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[403]),
        .S(self_sf7[403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[404]),
        .S(self_sf7[404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[405]),
        .S(self_sf7[405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[406]),
        .S(self_sf7[406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[407]),
        .S(self_sf7[407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[408]),
        .S(self_sf7[408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[409]),
        .S(self_sf7[409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[40].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[40]),
        .S(self_sf7[40]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[410]),
        .S(self_sf7[410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[411]),
        .S(self_sf7[411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[412]),
        .S(self_sf7[412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[413]),
        .S(self_sf7[413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[414]),
        .S(self_sf7[414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[415]),
        .S(self_sf7[415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[416]),
        .S(self_sf7[416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[417]),
        .S(self_sf7[417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[418]),
        .S(self_sf7[418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[419]),
        .S(self_sf7[419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[41].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[41]),
        .S(self_sf7[41]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[420]),
        .S(self_sf7[420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[421]),
        .S(self_sf7[421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[422]),
        .S(self_sf7[422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[423]),
        .S(self_sf7[423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[424]),
        .S(self_sf7[424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[425]),
        .S(self_sf7[425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[426]),
        .S(self_sf7[426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[427]),
        .S(self_sf7[427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[428]),
        .S(self_sf7[428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[429]),
        .S(self_sf7[429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[42].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[42]),
        .S(self_sf7[42]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[430]),
        .S(self_sf7[430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[431]),
        .S(self_sf7[431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[432]),
        .S(self_sf7[432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[433]),
        .S(self_sf7[433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[434]),
        .S(self_sf7[434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[435]),
        .S(self_sf7[435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[436]),
        .S(self_sf7[436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[437]),
        .S(self_sf7[437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[438]),
        .S(self_sf7[438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[439]),
        .S(self_sf7[439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[43].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[43]),
        .S(self_sf7[43]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[440]),
        .S(self_sf7[440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[441]),
        .S(self_sf7[441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[442]),
        .S(self_sf7[442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[443]),
        .S(self_sf7[443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[444]),
        .S(self_sf7[444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[445]),
        .S(self_sf7[445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[446]),
        .S(self_sf7[446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[447]),
        .S(self_sf7[447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[448]),
        .S(self_sf7[448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[449]),
        .S(self_sf7[449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[44].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[44]),
        .S(self_sf7[44]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[450]),
        .S(self_sf7[450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[451]),
        .S(self_sf7[451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[452]),
        .S(self_sf7[452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[453]),
        .S(self_sf7[453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[454]),
        .S(self_sf7[454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[455]),
        .S(self_sf7[455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[456]),
        .S(self_sf7[456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[457]),
        .S(self_sf7[457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[458]),
        .S(self_sf7[458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[459]),
        .S(self_sf7[459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[45].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[45]),
        .S(self_sf7[45]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[460]),
        .S(self_sf7[460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[461]),
        .S(self_sf7[461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[462]),
        .S(self_sf7[462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[463]),
        .S(self_sf7[463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[464]),
        .S(self_sf7[464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[465]),
        .S(self_sf7[465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[466]),
        .S(self_sf7[466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[467]),
        .S(self_sf7[467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[468]),
        .S(self_sf7[468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[469]),
        .S(self_sf7[469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[46].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[46]),
        .S(self_sf7[46]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[470]),
        .S(self_sf7[470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[471]),
        .S(self_sf7[471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[472]),
        .S(self_sf7[472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[473]),
        .S(self_sf7[473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[474]),
        .S(self_sf7[474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[475]),
        .S(self_sf7[475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[476]),
        .S(self_sf7[476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[477]),
        .S(self_sf7[477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[478]),
        .S(self_sf7[478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[479]),
        .S(self_sf7[479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[47].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[47]),
        .S(self_sf7[47]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[480]),
        .S(self_sf7[480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[481]),
        .S(self_sf7[481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[482]),
        .S(self_sf7[482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[483]),
        .S(self_sf7[483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[484]),
        .S(self_sf7[484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[485]),
        .S(self_sf7[485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[486]),
        .S(self_sf7[486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[487]),
        .S(self_sf7[487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[488]),
        .S(self_sf7[488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[489]),
        .S(self_sf7[489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[48].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[48]),
        .S(self_sf7[48]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[490]),
        .S(self_sf7[490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[491]),
        .S(self_sf7[491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[492]),
        .S(self_sf7[492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[493]),
        .S(self_sf7[493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[494]),
        .S(self_sf7[494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[495]),
        .S(self_sf7[495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[496]),
        .S(self_sf7[496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[497]),
        .S(self_sf7[497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[498]),
        .S(self_sf7[498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[499]),
        .S(self_sf7[499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[49].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[49]),
        .S(self_sf7[49]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[4].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[4]),
        .S(info_sf7[4]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[500]),
        .S(self_sf7[500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[501]),
        .S(self_sf7[501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[502]),
        .S(self_sf7[502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[503]),
        .S(self_sf7[503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[504]),
        .S(self_sf7[504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[505]),
        .S(self_sf7[505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[506]),
        .S(self_sf7[506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[507]),
        .S(self_sf7[507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[508]),
        .S(self_sf7[508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[509]),
        .S(self_sf7[509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[50].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[50]),
        .S(self_sf7[50]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[510]),
        .S(self_sf7[510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[511]),
        .S(self_sf7[511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[512]),
        .S(self_sf7[512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[513]),
        .S(self_sf7[513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[514]),
        .S(self_sf7[514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[515]),
        .S(self_sf7[515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[516]),
        .S(self_sf7[516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[517]),
        .S(self_sf7[517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[518]),
        .S(self_sf7[518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[519]),
        .S(self_sf7[519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[51].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[51]),
        .S(self_sf7[51]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[520]),
        .S(self_sf7[520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[521]),
        .S(self_sf7[521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[522]),
        .S(self_sf7[522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[523]),
        .S(self_sf7[523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[524]),
        .S(self_sf7[524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[525]),
        .S(self_sf7[525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[526]),
        .S(self_sf7[526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[527]),
        .S(self_sf7[527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[528]),
        .S(self_sf7[528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[529]),
        .S(self_sf7[529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[52].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[52]),
        .S(self_sf7[52]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[530]),
        .S(self_sf7[530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[531]),
        .S(self_sf7[531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[532]),
        .S(self_sf7[532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[533]),
        .S(self_sf7[533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[534]),
        .S(self_sf7[534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[535]),
        .S(self_sf7[535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[536]),
        .S(self_sf7[536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[537]),
        .S(self_sf7[537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[538]),
        .S(self_sf7[538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[539]),
        .S(self_sf7[539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[53].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[53]),
        .S(self_sf7[53]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[540]),
        .S(self_sf7[540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[541]),
        .S(self_sf7[541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[542]),
        .S(self_sf7[542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[543]),
        .S(self_sf7[543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[544]),
        .S(self_sf7[544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[545]),
        .S(self_sf7[545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[546]),
        .S(self_sf7[546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[547]),
        .S(self_sf7[547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[548]),
        .S(self_sf7[548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[549]),
        .S(self_sf7[549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[54].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[54]),
        .S(self_sf7[54]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[550]),
        .S(self_sf7[550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[551]),
        .S(self_sf7[551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[552]),
        .S(self_sf7[552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[553]),
        .S(self_sf7[553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[554]),
        .S(self_sf7[554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[555]),
        .S(self_sf7[555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[556]),
        .S(self_sf7[556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[557]),
        .S(self_sf7[557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[558]),
        .S(self_sf7[558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[559]),
        .S(self_sf7[559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[55].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[55]),
        .S(self_sf7[55]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[560]),
        .S(self_sf7[560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[561]),
        .S(self_sf7[561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[562]),
        .S(self_sf7[562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[563]),
        .S(self_sf7[563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[564]),
        .S(self_sf7[564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[565]),
        .S(self_sf7[565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[566]),
        .S(self_sf7[566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[567]),
        .S(self_sf7[567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[568]),
        .S(self_sf7[568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[569]),
        .S(self_sf7[569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[56].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[56]),
        .S(self_sf7[56]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[570]),
        .S(self_sf7[570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[571]),
        .S(self_sf7[571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[572]),
        .S(self_sf7[572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[573]),
        .S(self_sf7[573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[574]),
        .S(self_sf7[574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[575]),
        .S(self_sf7[575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[576]),
        .S(self_sf7[576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[577]),
        .S(self_sf7[577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[578]),
        .S(self_sf7[578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[579]),
        .S(self_sf7[579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[57].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[57]),
        .S(self_sf7[57]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[580]),
        .S(self_sf7[580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[581]),
        .S(self_sf7[581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[582]),
        .S(self_sf7[582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[583]),
        .S(self_sf7[583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[584]),
        .S(self_sf7[584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[585]),
        .S(self_sf7[585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[586]),
        .S(self_sf7[586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[587]),
        .S(self_sf7[587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[588]),
        .S(self_sf7[588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[589]),
        .S(self_sf7[589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[58].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[58]),
        .S(self_sf7[58]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[590]),
        .S(self_sf7[590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[591]),
        .S(self_sf7[591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[592]),
        .S(self_sf7[592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[593]),
        .S(self_sf7[593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[594]),
        .S(self_sf7[594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[595]),
        .S(self_sf7[595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[596]),
        .S(self_sf7[596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[597]),
        .S(self_sf7[597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[598]),
        .S(self_sf7[598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[599]),
        .S(self_sf7[599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[59].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[59]),
        .S(self_sf7[59]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[5].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[5]),
        .S(info_sf7[5]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[600]),
        .S(self_sf7[600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[601]),
        .S(self_sf7[601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[602]),
        .S(self_sf7[602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[603]),
        .S(self_sf7[603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[604]),
        .S(self_sf7[604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[605]),
        .S(self_sf7[605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[606]),
        .S(self_sf7[606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[607]),
        .S(self_sf7[607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[608]),
        .S(self_sf7[608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[609]),
        .S(self_sf7[609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[60].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[60]),
        .S(self_sf7[60]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[610]),
        .S(self_sf7[610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[611]),
        .S(self_sf7[611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[612]),
        .S(self_sf7[612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[613]),
        .S(self_sf7[613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[614]),
        .S(self_sf7[614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[615]),
        .S(self_sf7[615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[616]),
        .S(self_sf7[616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[617]),
        .S(self_sf7[617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[618]),
        .S(self_sf7[618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[619]),
        .S(self_sf7[619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[61].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[61]),
        .S(self_sf7[61]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[620]),
        .S(self_sf7[620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[621]),
        .S(self_sf7[621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[622]),
        .S(self_sf7[622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[623]),
        .S(self_sf7[623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[624]),
        .S(self_sf7[624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[625]),
        .S(self_sf7[625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[626]),
        .S(self_sf7[626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[627]),
        .S(self_sf7[627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[628]),
        .S(self_sf7[628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[629]),
        .S(self_sf7[629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[62].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[62]),
        .S(self_sf7[62]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[630]),
        .S(self_sf7[630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[631]),
        .S(self_sf7[631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[632]),
        .S(self_sf7[632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[633]),
        .S(self_sf7[633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[634]),
        .S(self_sf7[634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[635]),
        .S(self_sf7[635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[636]),
        .S(self_sf7[636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[637]),
        .S(self_sf7[637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[638]),
        .S(self_sf7[638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[639]),
        .S(self_sf7[639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[63].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[63]),
        .S(self_sf7[63]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[640]),
        .S(self_sf7[640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[641]),
        .S(self_sf7[641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[642]),
        .S(self_sf7[642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[643]),
        .S(self_sf7[643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[644]),
        .S(self_sf7[644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[645]),
        .S(self_sf7[645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[646]),
        .S(self_sf7[646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[647]),
        .S(self_sf7[647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[648]),
        .S(self_sf7[648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[649]),
        .S(self_sf7[649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[64].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[64]),
        .S(self_sf7[64]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[650]),
        .S(self_sf7[650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[651]),
        .S(self_sf7[651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[652]),
        .S(self_sf7[652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[653]),
        .S(self_sf7[653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[654]),
        .S(self_sf7[654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[655]),
        .S(self_sf7[655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[656]),
        .S(self_sf7[656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[657]),
        .S(self_sf7[657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[658]),
        .S(self_sf7[658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[659]),
        .S(self_sf7[659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[65].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[65]),
        .S(self_sf7[65]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[660]),
        .S(self_sf7[660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[661]),
        .S(self_sf7[661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[662]),
        .S(self_sf7[662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[663]),
        .S(self_sf7[663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[664]),
        .S(self_sf7[664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[665]),
        .S(self_sf7[665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[666]),
        .S(self_sf7[666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[667]),
        .S(self_sf7[667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[668]),
        .S(self_sf7[668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[669]),
        .S(self_sf7[669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[66].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[66]),
        .S(self_sf7[66]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[670]),
        .S(self_sf7[670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[671]),
        .S(self_sf7[671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[672]),
        .S(self_sf7[672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[673]),
        .S(self_sf7[673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[674]),
        .S(self_sf7[674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[675]),
        .S(self_sf7[675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[676]),
        .S(self_sf7[676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[677]),
        .S(self_sf7[677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[678]),
        .S(self_sf7[678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[679]),
        .S(self_sf7[679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[67].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[67]),
        .S(self_sf7[67]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[680]),
        .S(self_sf7[680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[681]),
        .S(self_sf7[681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[682]),
        .S(self_sf7[682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[683]),
        .S(self_sf7[683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[684]),
        .S(self_sf7[684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[685]),
        .S(self_sf7[685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[686]),
        .S(self_sf7[686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[687]),
        .S(self_sf7[687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[688]),
        .S(self_sf7[688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[689]),
        .S(self_sf7[689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[68].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[68]),
        .S(self_sf7[68]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[690]),
        .S(self_sf7[690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[691]),
        .S(self_sf7[691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[692]),
        .S(self_sf7[692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[693]),
        .S(self_sf7[693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[694]),
        .S(self_sf7[694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[695]),
        .S(self_sf7[695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[696]),
        .S(self_sf7[696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[697]),
        .S(self_sf7[697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[698]),
        .S(self_sf7[698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[699]),
        .S(self_sf7[699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[69].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[69]),
        .S(self_sf7[69]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[6].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[6]),
        .S(info_sf7[6]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[700]),
        .S(self_sf7[700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[701]),
        .S(self_sf7[701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[702]),
        .S(self_sf7[702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[703]),
        .S(self_sf7[703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[704]),
        .S(self_sf7[704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[705]),
        .S(self_sf7[705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[706]),
        .S(self_sf7[706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[707]),
        .S(self_sf7[707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[708]),
        .S(self_sf7[708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[709]),
        .S(self_sf7[709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[70].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[70]),
        .S(self_sf7[70]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[710]),
        .S(self_sf7[710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[711]),
        .S(self_sf7[711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[712]),
        .S(self_sf7[712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[713]),
        .S(self_sf7[713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[714]),
        .S(self_sf7[714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[715]),
        .S(self_sf7[715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[716]),
        .S(self_sf7[716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[717]),
        .S(self_sf7[717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[718]),
        .S(self_sf7[718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[719]),
        .S(self_sf7[719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[71].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[71]),
        .S(self_sf7[71]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[720]),
        .S(self_sf7[720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[721]),
        .S(self_sf7[721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[722]),
        .S(self_sf7[722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[723]),
        .S(self_sf7[723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[724]),
        .S(self_sf7[724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[725]),
        .S(self_sf7[725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[726]),
        .S(self_sf7[726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[727]),
        .S(self_sf7[727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[728]),
        .S(self_sf7[728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[729]),
        .S(self_sf7[729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[72].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[72]),
        .S(self_sf7[72]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[730]),
        .S(self_sf7[730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[731]),
        .S(self_sf7[731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[732]),
        .S(self_sf7[732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[733]),
        .S(self_sf7[733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[734]),
        .S(self_sf7[734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[735]),
        .S(self_sf7[735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[736]),
        .S(self_sf7[736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[737]),
        .S(self_sf7[737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[738]),
        .S(self_sf7[738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[739]),
        .S(self_sf7[739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[73].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[73]),
        .S(self_sf7[73]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[740]),
        .S(self_sf7[740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[741]),
        .S(self_sf7[741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[742]),
        .S(self_sf7[742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[743]),
        .S(self_sf7[743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[744]),
        .S(self_sf7[744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[745]),
        .S(self_sf7[745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[746]),
        .S(self_sf7[746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[747]),
        .S(self_sf7[747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[748]),
        .S(self_sf7[748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[749]),
        .S(self_sf7[749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[74].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[74]),
        .S(self_sf7[74]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[750]),
        .S(self_sf7[750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[751]),
        .S(self_sf7[751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[752]),
        .S(self_sf7[752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[753]),
        .S(self_sf7[753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[754]),
        .S(self_sf7[754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[755]),
        .S(self_sf7[755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[756]),
        .S(self_sf7[756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[757]),
        .S(self_sf7[757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[758]),
        .S(self_sf7[758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[759]),
        .S(self_sf7[759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[75].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[75]),
        .S(self_sf7[75]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[760]),
        .S(self_sf7[760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[761]),
        .S(self_sf7[761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[762]),
        .S(self_sf7[762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[763]),
        .S(self_sf7[763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[764]),
        .S(self_sf7[764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[765]),
        .S(self_sf7[765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[766]),
        .S(self_sf7[766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[767]),
        .S(self_sf7[767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[768]),
        .S(self_sf7[768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[769]),
        .S(self_sf7[769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[76].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[76]),
        .S(self_sf7[76]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[770]),
        .S(self_sf7[770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[771]),
        .S(self_sf7[771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[772]),
        .S(self_sf7[772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[773]),
        .S(self_sf7[773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[774]),
        .S(self_sf7[774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[775]),
        .S(self_sf7[775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[776]),
        .S(self_sf7[776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[777]),
        .S(self_sf7[777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[778]),
        .S(self_sf7[778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[779]),
        .S(self_sf7[779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[77].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[77]),
        .S(self_sf7[77]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[780]),
        .S(self_sf7[780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[781]),
        .S(self_sf7[781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[782]),
        .S(self_sf7[782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[783]),
        .S(self_sf7[783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[784]),
        .S(self_sf7[784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[785]),
        .S(self_sf7[785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[786]),
        .S(self_sf7[786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[787]),
        .S(self_sf7[787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[788]),
        .S(self_sf7[788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[789]),
        .S(self_sf7[789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[78].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[78]),
        .S(self_sf7[78]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[790]),
        .S(self_sf7[790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[791]),
        .S(self_sf7[791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[792]),
        .S(self_sf7[792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[793]),
        .S(self_sf7[793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[794]),
        .S(self_sf7[794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[795]),
        .S(self_sf7[795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[796]),
        .S(self_sf7[796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[797]),
        .S(self_sf7[797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[798]),
        .S(self_sf7[798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[799]),
        .S(self_sf7[799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[79].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[79]),
        .S(self_sf7[79]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[7].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[7]),
        .S(info_sf7[7]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[800].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[800]),
        .S(self_sf7[800]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[801].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[801]),
        .S(self_sf7[801]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[802].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[802]),
        .S(self_sf7[802]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[803].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[803]),
        .S(self_sf7[803]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[804].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[804]),
        .S(self_sf7[804]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[805].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[805]),
        .S(self_sf7[805]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[806].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[806]),
        .S(self_sf7[806]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[807].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[807]),
        .S(self_sf7[807]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[808].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[808]),
        .S(self_sf7[808]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[809].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[809]),
        .S(self_sf7[809]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[80].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[80]),
        .S(self_sf7[80]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[810].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[810]),
        .S(self_sf7[810]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[811].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[811]),
        .S(self_sf7[811]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[812].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[812]),
        .S(self_sf7[812]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[813].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[813]),
        .S(self_sf7[813]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[814].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[814]),
        .S(self_sf7[814]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[815].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[815]),
        .S(self_sf7[815]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[816].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[816]),
        .S(self_sf7[816]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[817].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[817]),
        .S(self_sf7[817]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[818].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[818]),
        .S(self_sf7[818]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[819].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[819]),
        .S(self_sf7[819]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[81].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[81]),
        .S(self_sf7[81]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[820].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[820]),
        .S(self_sf7[820]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[821].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[821]),
        .S(self_sf7[821]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[822].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[822]),
        .S(self_sf7[822]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[823].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[823]),
        .S(self_sf7[823]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[824].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[824]),
        .S(self_sf7[824]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[825].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[825]),
        .S(self_sf7[825]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[826].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[826]),
        .S(self_sf7[826]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[827].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[827]),
        .S(self_sf7[827]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[828].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[828]),
        .S(self_sf7[828]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[829].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[829]),
        .S(self_sf7[829]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[82].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[82]),
        .S(self_sf7[82]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[830].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[830]),
        .S(self_sf7[830]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[831].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[831]),
        .S(self_sf7[831]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[832].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[832]),
        .S(self_sf7[832]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[833].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[833]),
        .S(self_sf7[833]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[834].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[834]),
        .S(self_sf7[834]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[835].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[835]),
        .S(self_sf7[835]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[836].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[836]),
        .S(self_sf7[836]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[837].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[837]),
        .S(self_sf7[837]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[838].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[838]),
        .S(self_sf7[838]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[839].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[839]),
        .S(self_sf7[839]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[83].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[83]),
        .S(self_sf7[83]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[840].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[840]),
        .S(self_sf7[840]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[841].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[841]),
        .S(self_sf7[841]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[842].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[842]),
        .S(self_sf7[842]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[843].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[843]),
        .S(self_sf7[843]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[844].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[844]),
        .S(self_sf7[844]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[845].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[845]),
        .S(self_sf7[845]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[846].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[846]),
        .S(self_sf7[846]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[847].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[847]),
        .S(self_sf7[847]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[848].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[848]),
        .S(self_sf7[848]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[849].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[849]),
        .S(self_sf7[849]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[84].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[84]),
        .S(self_sf7[84]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[850].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[850]),
        .S(self_sf7[850]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[851].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[851]),
        .S(self_sf7[851]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[852].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[852]),
        .S(self_sf7[852]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[853].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[853]),
        .S(self_sf7[853]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[854].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[854]),
        .S(self_sf7[854]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[855].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[855]),
        .S(self_sf7[855]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[856].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[856]),
        .S(self_sf7[856]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[857].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[857]),
        .S(self_sf7[857]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[858].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[858]),
        .S(self_sf7[858]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[859].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[859]),
        .S(self_sf7[859]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[85].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[85]),
        .S(self_sf7[85]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[860].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[860]),
        .S(self_sf7[860]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[861].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[861]),
        .S(self_sf7[861]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[862].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[862]),
        .S(self_sf7[862]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[863].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[863]),
        .S(self_sf7[863]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[864].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[864]),
        .S(self_sf7[864]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[865].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[865]),
        .S(self_sf7[865]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[866].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[866]),
        .S(self_sf7[866]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[867].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[867]),
        .S(self_sf7[867]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[868].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[868]),
        .S(self_sf7[868]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[869].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[869]),
        .S(self_sf7[869]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[86].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[86]),
        .S(self_sf7[86]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[870].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[870]),
        .S(self_sf7[870]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[871].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[871]),
        .S(self_sf7[871]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[872].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[872]),
        .S(self_sf7[872]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[873].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[873]),
        .S(self_sf7[873]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[874].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[874]),
        .S(self_sf7[874]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[875].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[875]),
        .S(self_sf7[875]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[876].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[876]),
        .S(self_sf7[876]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[877].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[877]),
        .S(self_sf7[877]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[878].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[878]),
        .S(self_sf7[878]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[879].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[879]),
        .S(self_sf7[879]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[87].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[87]),
        .S(self_sf7[87]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[880].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[880]),
        .S(self_sf7[880]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[881].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[881]),
        .S(self_sf7[881]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[882].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[882]),
        .S(self_sf7[882]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[883].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[883]),
        .S(self_sf7[883]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[884].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[884]),
        .S(self_sf7[884]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[885].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[885]),
        .S(self_sf7[885]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[886].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[886]),
        .S(self_sf7[886]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[887].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[887]),
        .S(self_sf7[887]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[888].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[888]),
        .S(self_sf7[888]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[889].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[889]),
        .S(self_sf7[889]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[88].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[88]),
        .S(self_sf7[88]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[890].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[890]),
        .S(self_sf7[890]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[891].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[891]),
        .S(self_sf7[891]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[892].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[892]),
        .S(self_sf7[892]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[893].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[893]),
        .S(self_sf7[893]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[894].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[894]),
        .S(self_sf7[894]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[895].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[895]),
        .S(self_sf7[895]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[896].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[896]),
        .S(self_sf7[896]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[897].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[897]),
        .S(self_sf7[897]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[898].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[898]),
        .S(self_sf7[898]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[899].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[899]),
        .S(self_sf7[899]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[89].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[89]),
        .S(self_sf7[89]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[8].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[8]),
        .S(self_sf7[8]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[900].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[900]),
        .S(self_sf7[900]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[901].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[901]),
        .S(self_sf7[901]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[902].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[902]),
        .S(self_sf7[902]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[903].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[903]),
        .S(self_sf7[903]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[904].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[904]),
        .S(self_sf7[904]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[905].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[905]),
        .S(self_sf7[905]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[906].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[906]),
        .S(self_sf7[906]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[907].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[907]),
        .S(self_sf7[907]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[908].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[908]),
        .S(self_sf7[908]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[909].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[909]),
        .S(self_sf7[909]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[90].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[90]),
        .S(self_sf7[90]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[910].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[910]),
        .S(self_sf7[910]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[911].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[911]),
        .S(self_sf7[911]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[912].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[912]),
        .S(self_sf7[912]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[913].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[913]),
        .S(self_sf7[913]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[914].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[914]),
        .S(self_sf7[914]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[915].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[915]),
        .S(self_sf7[915]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[916].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[916]),
        .S(self_sf7[916]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[917].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[917]),
        .S(self_sf7[917]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[918].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[918]),
        .S(self_sf7[918]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[919].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[919]),
        .S(self_sf7[919]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[91].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[91]),
        .S(self_sf7[91]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[920].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[920]),
        .S(self_sf7[920]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[921].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[921]),
        .S(self_sf7[921]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[922].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[922]),
        .S(self_sf7[922]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[923].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[923]),
        .S(self_sf7[923]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[924].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[924]),
        .S(self_sf7[924]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[925].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[925]),
        .S(self_sf7[925]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[926].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[926]),
        .S(self_sf7[926]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[927].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[927]),
        .S(self_sf7[927]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[928].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[928]),
        .S(self_sf7[928]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[929].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[929]),
        .S(self_sf7[929]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[92].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[92]),
        .S(self_sf7[92]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[930].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[930]),
        .S(self_sf7[930]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[931].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[931]),
        .S(self_sf7[931]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[932].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[932]),
        .S(self_sf7[932]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[933].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[933]),
        .S(self_sf7[933]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[934].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[934]),
        .S(self_sf7[934]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[935].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[935]),
        .S(self_sf7[935]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[936].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[936]),
        .S(self_sf7[936]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[937].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[937]),
        .S(self_sf7[937]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[938].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[938]),
        .S(self_sf7[938]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[939].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[939]),
        .S(self_sf7[939]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[93].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[93]),
        .S(self_sf7[93]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[940].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[940]),
        .S(self_sf7[940]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[941].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[941]),
        .S(self_sf7[941]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[942].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[942]),
        .S(self_sf7[942]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[943].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[943]),
        .S(self_sf7[943]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[944].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[944]),
        .S(self_sf7[944]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[945].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[945]),
        .S(self_sf7[945]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[946].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[946]),
        .S(self_sf7[946]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[947].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[947]),
        .S(self_sf7[947]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[948].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[948]),
        .S(self_sf7[948]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[949].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[949]),
        .S(self_sf7[949]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[94].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[94]),
        .S(self_sf7[94]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[950].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[950]),
        .S(self_sf7[950]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[951].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[951]),
        .S(self_sf7[951]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[952].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[952]),
        .S(self_sf7[952]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[953].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[953]),
        .S(self_sf7[953]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[954].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[954]),
        .S(self_sf7[954]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[955].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[955]),
        .S(self_sf7[955]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[956].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[956]),
        .S(self_sf7[956]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[957].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[957]),
        .S(self_sf7[957]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[958].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[958]),
        .S(self_sf7[958]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[959].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[959]),
        .S(self_sf7[959]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[95].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[95]),
        .S(self_sf7[95]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[960].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[960]),
        .S(self_sf7[960]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[961].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[961]),
        .S(self_sf7[961]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[962].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[962]),
        .S(self_sf7[962]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[963].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[963]),
        .S(self_sf7[963]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[964].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[964]),
        .S(self_sf7[964]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[965].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[965]),
        .S(self_sf7[965]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[966].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[966]),
        .S(self_sf7[966]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[967].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[967]),
        .S(self_sf7[967]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[968].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[968]),
        .S(self_sf7[968]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[969].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[969]),
        .S(self_sf7[969]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[96].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[96]),
        .S(self_sf7[96]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[970].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[970]),
        .S(self_sf7[970]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[971].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[971]),
        .S(self_sf7[971]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[972].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[972]),
        .S(self_sf7[972]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[973].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[973]),
        .S(self_sf7[973]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[974].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[974]),
        .S(self_sf7[974]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[975].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[975]),
        .S(self_sf7[975]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[976].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[976]),
        .S(self_sf7[976]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[977].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[977]),
        .S(self_sf7[977]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[978].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[978]),
        .S(self_sf7[978]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[979].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[979]),
        .S(self_sf7[979]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[97].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[97]),
        .S(self_sf7[97]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[980].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[980]),
        .S(self_sf7[980]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[981].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[981]),
        .S(self_sf7[981]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[982].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[982]),
        .S(self_sf7[982]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[983].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[983]),
        .S(self_sf7[983]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[984].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[984]),
        .S(self_sf7[984]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[985].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[985]),
        .S(self_sf7[985]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[986].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[986]),
        .S(self_sf7[986]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[987].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[987]),
        .S(self_sf7[987]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[988].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[988]),
        .S(self_sf7[988]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[989].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[989]),
        .S(self_sf7[989]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[98].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[98]),
        .S(self_sf7[98]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[990].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[990]),
        .S(self_sf7[990]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[991].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[991]),
        .S(self_sf7[991]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[992].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[992]),
        .S(self_sf7[992]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[993].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[993]),
        .S(self_sf7[993]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[994].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[994]),
        .S(self_sf7[994]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[995].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[995]),
        .S(self_sf7[995]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[996].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[996]),
        .S(self_sf7[996]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[997].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[997]),
        .S(self_sf7[997]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[998].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[998]),
        .S(self_sf7[998]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[999].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[999]),
        .S(self_sf7[999]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[99].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[99]),
        .S(self_sf7[99]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[9].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[9]),
        .S(self_sf7[9]));
  (* BOX_TYPE = "black_box" *) 
  MUXF8 \activity_ROsf8[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf8[0]),
        .S(self_sf8[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF9 \activity_ROsf9[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf9[0]),
        .S(self_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_0
       (.I0(1'b0),
        .O(self_sf7[1802]));
  LUT1 #(
    .INIT(2'h2)) 
    i_1
       (.I0(1'b0),
        .O(self_sf7[1801]));
  LUT1 #(
    .INIT(2'h2)) 
    i_10
       (.I0(1'b0),
        .O(info_sf8[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_11
       (.I0(1'b0),
        .O(info_sf8[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_12
       (.I0(1'b0),
        .O(info_sf8[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_13
       (.I0(1'b0),
        .O(info_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_14
       (.I0(1'b0),
        .O(info_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_15
       (.I0(1'b0),
        .O(info_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_16
       (.I0(1'b0),
        .O(info_sf8[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_17
       (.I0(1'b0),
        .O(info_sf9[7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_18
       (.I0(1'b0),
        .O(info_sf9[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_19
       (.I0(1'b0),
        .O(info_sf9[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_2
       (.I0(1'b0),
        .O(self_sf7[1800]));
  LUT1 #(
    .INIT(2'h2)) 
    i_20
       (.I0(1'b0),
        .O(info_sf9[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_21
       (.I0(1'b0),
        .O(info_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_22
       (.I0(1'b0),
        .O(info_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_23
       (.I0(1'b0),
        .O(info_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_24
       (.I0(1'b0),
        .O(info_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_3
       (.I0(1'b0),
        .O(self_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_4
       (.I0(1'b0),
        .O(self_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_5
       (.I0(1'b0),
        .O(self_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_6
       (.I0(1'b0),
        .O(self_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_7
       (.I0(1'b0),
        .O(self_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_8
       (.I0(1'b0),
        .O(self_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_9
       (.I0(1'b0),
        .O(info_sf8[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst
       (.I0(self_sf7[7]),
        .O(info_sf7[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__0
       (.I0(self_sf7[6]),
        .O(info_sf7[6]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__1
       (.I0(self_sf7[5]),
        .O(info_sf7[5]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__2
       (.I0(self_sf7[4]),
        .O(info_sf7[4]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__3
       (.I0(self_sf7[3]),
        .O(info_sf7[3]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__4
       (.I0(self_sf7[2]),
        .O(info_sf7[2]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__5
       (.I0(self_sf7[1]),
        .O(info_sf7[1]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__6
       (.I0(self_sf7[0]),
        .O(info_sf7[0]));
endmodule

(* ORIG_REF_NAME = "muxer" *) (* box_type = "black_box" *) (* dont_touch = "true" *) 
module switch_elements_muxer__5
   (enable_i,
    info_o);
  input enable_i;
  output info_o;

  wire enable_i;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf7;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf8;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf9;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [1802:0]self_sf7;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf8;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf9;

  assign info_o = info_sf7[1];
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[0]),
        .S(info_sf7[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1000].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1000]),
        .S(self_sf7[1000]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1001].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1001]),
        .S(self_sf7[1001]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1002].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1002]),
        .S(self_sf7[1002]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1003].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1003]),
        .S(self_sf7[1003]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1004].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1004]),
        .S(self_sf7[1004]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1005].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1005]),
        .S(self_sf7[1005]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1006].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1006]),
        .S(self_sf7[1006]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1007].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1007]),
        .S(self_sf7[1007]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1008].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1008]),
        .S(self_sf7[1008]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1009].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1009]),
        .S(self_sf7[1009]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[100]),
        .S(self_sf7[100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1010].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1010]),
        .S(self_sf7[1010]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1011].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1011]),
        .S(self_sf7[1011]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1012].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1012]),
        .S(self_sf7[1012]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1013].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1013]),
        .S(self_sf7[1013]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1014].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1014]),
        .S(self_sf7[1014]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1015].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1015]),
        .S(self_sf7[1015]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1016].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1016]),
        .S(self_sf7[1016]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1017].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1017]),
        .S(self_sf7[1017]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1018].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1018]),
        .S(self_sf7[1018]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1019].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1019]),
        .S(self_sf7[1019]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[101]),
        .S(self_sf7[101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1020].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1020]),
        .S(self_sf7[1020]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1021].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1021]),
        .S(self_sf7[1021]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1022].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1022]),
        .S(self_sf7[1022]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1023].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1023]),
        .S(self_sf7[1023]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1024].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1024]),
        .S(self_sf7[1024]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1025].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1025]),
        .S(self_sf7[1025]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1026].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1026]),
        .S(self_sf7[1026]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1027].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1027]),
        .S(self_sf7[1027]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1028].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1028]),
        .S(self_sf7[1028]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1029].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1029]),
        .S(self_sf7[1029]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[102]),
        .S(self_sf7[102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1030].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1030]),
        .S(self_sf7[1030]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1031].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1031]),
        .S(self_sf7[1031]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1032].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1032]),
        .S(self_sf7[1032]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1033].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1033]),
        .S(self_sf7[1033]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1034].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1034]),
        .S(self_sf7[1034]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1035].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1035]),
        .S(self_sf7[1035]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1036].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1036]),
        .S(self_sf7[1036]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1037].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1037]),
        .S(self_sf7[1037]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1038].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1038]),
        .S(self_sf7[1038]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1039].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1039]),
        .S(self_sf7[1039]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[103]),
        .S(self_sf7[103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1040].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1040]),
        .S(self_sf7[1040]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1041].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1041]),
        .S(self_sf7[1041]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1042].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1042]),
        .S(self_sf7[1042]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1043].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1043]),
        .S(self_sf7[1043]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1044].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1044]),
        .S(self_sf7[1044]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1045].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1045]),
        .S(self_sf7[1045]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1046].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1046]),
        .S(self_sf7[1046]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1047].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1047]),
        .S(self_sf7[1047]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1048].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1048]),
        .S(self_sf7[1048]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1049].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1049]),
        .S(self_sf7[1049]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[104]),
        .S(self_sf7[104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1050].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1050]),
        .S(self_sf7[1050]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1051].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1051]),
        .S(self_sf7[1051]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1052].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1052]),
        .S(self_sf7[1052]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1053].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1053]),
        .S(self_sf7[1053]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1054].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1054]),
        .S(self_sf7[1054]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1055].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1055]),
        .S(self_sf7[1055]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1056].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1056]),
        .S(self_sf7[1056]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1057].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1057]),
        .S(self_sf7[1057]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1058].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1058]),
        .S(self_sf7[1058]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1059].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1059]),
        .S(self_sf7[1059]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[105]),
        .S(self_sf7[105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1060].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1060]),
        .S(self_sf7[1060]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1061].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1061]),
        .S(self_sf7[1061]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1062].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1062]),
        .S(self_sf7[1062]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1063].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1063]),
        .S(self_sf7[1063]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1064].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1064]),
        .S(self_sf7[1064]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1065].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1065]),
        .S(self_sf7[1065]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1066].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1066]),
        .S(self_sf7[1066]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1067].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1067]),
        .S(self_sf7[1067]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1068].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1068]),
        .S(self_sf7[1068]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1069].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1069]),
        .S(self_sf7[1069]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[106]),
        .S(self_sf7[106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1070].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1070]),
        .S(self_sf7[1070]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1071].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1071]),
        .S(self_sf7[1071]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1072].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1072]),
        .S(self_sf7[1072]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1073].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1073]),
        .S(self_sf7[1073]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1074].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1074]),
        .S(self_sf7[1074]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1075].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1075]),
        .S(self_sf7[1075]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1076].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1076]),
        .S(self_sf7[1076]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1077].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1077]),
        .S(self_sf7[1077]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1078].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1078]),
        .S(self_sf7[1078]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1079].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1079]),
        .S(self_sf7[1079]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[107]),
        .S(self_sf7[107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1080].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1080]),
        .S(self_sf7[1080]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1081].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1081]),
        .S(self_sf7[1081]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1082].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1082]),
        .S(self_sf7[1082]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1083].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1083]),
        .S(self_sf7[1083]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1084].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1084]),
        .S(self_sf7[1084]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1085].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1085]),
        .S(self_sf7[1085]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1086].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1086]),
        .S(self_sf7[1086]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1087].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1087]),
        .S(self_sf7[1087]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1088].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1088]),
        .S(self_sf7[1088]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1089].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1089]),
        .S(self_sf7[1089]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[108]),
        .S(self_sf7[108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1090].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1090]),
        .S(self_sf7[1090]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1091].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1091]),
        .S(self_sf7[1091]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1092].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1092]),
        .S(self_sf7[1092]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1093].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1093]),
        .S(self_sf7[1093]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1094].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1094]),
        .S(self_sf7[1094]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1095].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1095]),
        .S(self_sf7[1095]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1096].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1096]),
        .S(self_sf7[1096]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1097].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1097]),
        .S(self_sf7[1097]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1098].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1098]),
        .S(self_sf7[1098]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1099].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1099]),
        .S(self_sf7[1099]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[109]),
        .S(self_sf7[109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[10].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[10]),
        .S(self_sf7[10]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1100]),
        .S(self_sf7[1100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1101]),
        .S(self_sf7[1101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1102]),
        .S(self_sf7[1102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1103]),
        .S(self_sf7[1103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1104]),
        .S(self_sf7[1104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1105]),
        .S(self_sf7[1105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1106]),
        .S(self_sf7[1106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1107]),
        .S(self_sf7[1107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1108]),
        .S(self_sf7[1108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1109]),
        .S(self_sf7[1109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[110]),
        .S(self_sf7[110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1110]),
        .S(self_sf7[1110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1111]),
        .S(self_sf7[1111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1112]),
        .S(self_sf7[1112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1113]),
        .S(self_sf7[1113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1114]),
        .S(self_sf7[1114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1115]),
        .S(self_sf7[1115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1116]),
        .S(self_sf7[1116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1117]),
        .S(self_sf7[1117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1118]),
        .S(self_sf7[1118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1119]),
        .S(self_sf7[1119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[111]),
        .S(self_sf7[111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1120]),
        .S(self_sf7[1120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1121]),
        .S(self_sf7[1121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1122]),
        .S(self_sf7[1122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1123]),
        .S(self_sf7[1123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1124]),
        .S(self_sf7[1124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1125]),
        .S(self_sf7[1125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1126]),
        .S(self_sf7[1126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1127]),
        .S(self_sf7[1127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1128]),
        .S(self_sf7[1128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1129]),
        .S(self_sf7[1129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[112]),
        .S(self_sf7[112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1130]),
        .S(self_sf7[1130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1131]),
        .S(self_sf7[1131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1132]),
        .S(self_sf7[1132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1133]),
        .S(self_sf7[1133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1134]),
        .S(self_sf7[1134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1135]),
        .S(self_sf7[1135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1136]),
        .S(self_sf7[1136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1137]),
        .S(self_sf7[1137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1138]),
        .S(self_sf7[1138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1139]),
        .S(self_sf7[1139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[113]),
        .S(self_sf7[113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1140]),
        .S(self_sf7[1140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1141]),
        .S(self_sf7[1141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1142]),
        .S(self_sf7[1142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1143]),
        .S(self_sf7[1143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1144]),
        .S(self_sf7[1144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1145]),
        .S(self_sf7[1145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1146]),
        .S(self_sf7[1146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1147]),
        .S(self_sf7[1147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1148]),
        .S(self_sf7[1148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1149]),
        .S(self_sf7[1149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[114]),
        .S(self_sf7[114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1150]),
        .S(self_sf7[1150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1151]),
        .S(self_sf7[1151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1152]),
        .S(self_sf7[1152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1153]),
        .S(self_sf7[1153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1154]),
        .S(self_sf7[1154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1155]),
        .S(self_sf7[1155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1156]),
        .S(self_sf7[1156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1157]),
        .S(self_sf7[1157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1158]),
        .S(self_sf7[1158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1159]),
        .S(self_sf7[1159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[115]),
        .S(self_sf7[115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1160]),
        .S(self_sf7[1160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1161]),
        .S(self_sf7[1161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1162]),
        .S(self_sf7[1162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1163]),
        .S(self_sf7[1163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1164]),
        .S(self_sf7[1164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1165]),
        .S(self_sf7[1165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1166]),
        .S(self_sf7[1166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1167]),
        .S(self_sf7[1167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1168]),
        .S(self_sf7[1168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1169]),
        .S(self_sf7[1169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[116]),
        .S(self_sf7[116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1170]),
        .S(self_sf7[1170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1171]),
        .S(self_sf7[1171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1172]),
        .S(self_sf7[1172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1173]),
        .S(self_sf7[1173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1174]),
        .S(self_sf7[1174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1175]),
        .S(self_sf7[1175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1176]),
        .S(self_sf7[1176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1177]),
        .S(self_sf7[1177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1178]),
        .S(self_sf7[1178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1179]),
        .S(self_sf7[1179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[117]),
        .S(self_sf7[117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1180]),
        .S(self_sf7[1180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1181]),
        .S(self_sf7[1181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1182]),
        .S(self_sf7[1182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1183]),
        .S(self_sf7[1183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1184]),
        .S(self_sf7[1184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1185]),
        .S(self_sf7[1185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1186]),
        .S(self_sf7[1186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1187]),
        .S(self_sf7[1187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1188]),
        .S(self_sf7[1188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1189]),
        .S(self_sf7[1189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[118]),
        .S(self_sf7[118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1190]),
        .S(self_sf7[1190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1191]),
        .S(self_sf7[1191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1192]),
        .S(self_sf7[1192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1193]),
        .S(self_sf7[1193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1194]),
        .S(self_sf7[1194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1195]),
        .S(self_sf7[1195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1196]),
        .S(self_sf7[1196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1197]),
        .S(self_sf7[1197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1198]),
        .S(self_sf7[1198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1199]),
        .S(self_sf7[1199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[119]),
        .S(self_sf7[119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[11].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[11]),
        .S(self_sf7[11]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1200]),
        .S(self_sf7[1200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1201]),
        .S(self_sf7[1201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1202]),
        .S(self_sf7[1202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1203]),
        .S(self_sf7[1203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1204]),
        .S(self_sf7[1204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1205]),
        .S(self_sf7[1205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1206]),
        .S(self_sf7[1206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1207]),
        .S(self_sf7[1207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1208]),
        .S(self_sf7[1208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1209]),
        .S(self_sf7[1209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[120]),
        .S(self_sf7[120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1210]),
        .S(self_sf7[1210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1211]),
        .S(self_sf7[1211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1212]),
        .S(self_sf7[1212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1213]),
        .S(self_sf7[1213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1214]),
        .S(self_sf7[1214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1215]),
        .S(self_sf7[1215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1216]),
        .S(self_sf7[1216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1217]),
        .S(self_sf7[1217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1218]),
        .S(self_sf7[1218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1219]),
        .S(self_sf7[1219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[121]),
        .S(self_sf7[121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1220]),
        .S(self_sf7[1220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1221]),
        .S(self_sf7[1221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1222]),
        .S(self_sf7[1222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1223]),
        .S(self_sf7[1223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1224]),
        .S(self_sf7[1224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1225]),
        .S(self_sf7[1225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1226]),
        .S(self_sf7[1226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1227]),
        .S(self_sf7[1227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1228]),
        .S(self_sf7[1228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1229]),
        .S(self_sf7[1229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[122]),
        .S(self_sf7[122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1230]),
        .S(self_sf7[1230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1231]),
        .S(self_sf7[1231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1232]),
        .S(self_sf7[1232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1233]),
        .S(self_sf7[1233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1234]),
        .S(self_sf7[1234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1235]),
        .S(self_sf7[1235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1236]),
        .S(self_sf7[1236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1237]),
        .S(self_sf7[1237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1238]),
        .S(self_sf7[1238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1239]),
        .S(self_sf7[1239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[123]),
        .S(self_sf7[123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1240]),
        .S(self_sf7[1240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1241]),
        .S(self_sf7[1241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1242]),
        .S(self_sf7[1242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1243]),
        .S(self_sf7[1243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1244]),
        .S(self_sf7[1244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1245]),
        .S(self_sf7[1245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1246]),
        .S(self_sf7[1246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1247]),
        .S(self_sf7[1247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1248]),
        .S(self_sf7[1248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1249]),
        .S(self_sf7[1249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[124]),
        .S(self_sf7[124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1250]),
        .S(self_sf7[1250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1251]),
        .S(self_sf7[1251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1252]),
        .S(self_sf7[1252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1253]),
        .S(self_sf7[1253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1254]),
        .S(self_sf7[1254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1255]),
        .S(self_sf7[1255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1256]),
        .S(self_sf7[1256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1257]),
        .S(self_sf7[1257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1258]),
        .S(self_sf7[1258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1259]),
        .S(self_sf7[1259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[125]),
        .S(self_sf7[125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1260]),
        .S(self_sf7[1260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1261]),
        .S(self_sf7[1261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1262]),
        .S(self_sf7[1262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1263]),
        .S(self_sf7[1263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1264]),
        .S(self_sf7[1264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1265]),
        .S(self_sf7[1265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1266]),
        .S(self_sf7[1266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1267]),
        .S(self_sf7[1267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1268]),
        .S(self_sf7[1268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1269]),
        .S(self_sf7[1269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[126]),
        .S(self_sf7[126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1270]),
        .S(self_sf7[1270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1271]),
        .S(self_sf7[1271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1272]),
        .S(self_sf7[1272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1273]),
        .S(self_sf7[1273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1274]),
        .S(self_sf7[1274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1275]),
        .S(self_sf7[1275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1276]),
        .S(self_sf7[1276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1277]),
        .S(self_sf7[1277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1278]),
        .S(self_sf7[1278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1279]),
        .S(self_sf7[1279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[127]),
        .S(self_sf7[127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1280]),
        .S(self_sf7[1280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1281]),
        .S(self_sf7[1281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1282]),
        .S(self_sf7[1282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1283]),
        .S(self_sf7[1283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1284]),
        .S(self_sf7[1284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1285]),
        .S(self_sf7[1285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1286]),
        .S(self_sf7[1286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1287]),
        .S(self_sf7[1287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1288]),
        .S(self_sf7[1288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1289]),
        .S(self_sf7[1289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[128]),
        .S(self_sf7[128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1290]),
        .S(self_sf7[1290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1291]),
        .S(self_sf7[1291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1292]),
        .S(self_sf7[1292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1293]),
        .S(self_sf7[1293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1294]),
        .S(self_sf7[1294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1295]),
        .S(self_sf7[1295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1296]),
        .S(self_sf7[1296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1297]),
        .S(self_sf7[1297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1298]),
        .S(self_sf7[1298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1299]),
        .S(self_sf7[1299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[129]),
        .S(self_sf7[129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[12].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[12]),
        .S(self_sf7[12]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1300]),
        .S(self_sf7[1300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1301]),
        .S(self_sf7[1301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1302]),
        .S(self_sf7[1302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1303]),
        .S(self_sf7[1303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1304]),
        .S(self_sf7[1304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1305]),
        .S(self_sf7[1305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1306]),
        .S(self_sf7[1306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1307]),
        .S(self_sf7[1307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1308]),
        .S(self_sf7[1308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1309]),
        .S(self_sf7[1309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[130]),
        .S(self_sf7[130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1310]),
        .S(self_sf7[1310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1311]),
        .S(self_sf7[1311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1312]),
        .S(self_sf7[1312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1313]),
        .S(self_sf7[1313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1314]),
        .S(self_sf7[1314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1315]),
        .S(self_sf7[1315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1316]),
        .S(self_sf7[1316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1317]),
        .S(self_sf7[1317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1318]),
        .S(self_sf7[1318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1319]),
        .S(self_sf7[1319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[131]),
        .S(self_sf7[131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1320]),
        .S(self_sf7[1320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1321]),
        .S(self_sf7[1321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1322]),
        .S(self_sf7[1322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1323]),
        .S(self_sf7[1323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1324]),
        .S(self_sf7[1324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1325]),
        .S(self_sf7[1325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1326]),
        .S(self_sf7[1326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1327]),
        .S(self_sf7[1327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1328]),
        .S(self_sf7[1328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1329]),
        .S(self_sf7[1329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[132]),
        .S(self_sf7[132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1330]),
        .S(self_sf7[1330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1331]),
        .S(self_sf7[1331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1332]),
        .S(self_sf7[1332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1333]),
        .S(self_sf7[1333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1334]),
        .S(self_sf7[1334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1335]),
        .S(self_sf7[1335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1336]),
        .S(self_sf7[1336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1337]),
        .S(self_sf7[1337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1338]),
        .S(self_sf7[1338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1339]),
        .S(self_sf7[1339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[133]),
        .S(self_sf7[133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1340]),
        .S(self_sf7[1340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1341]),
        .S(self_sf7[1341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1342]),
        .S(self_sf7[1342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1343]),
        .S(self_sf7[1343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1344]),
        .S(self_sf7[1344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1345]),
        .S(self_sf7[1345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1346]),
        .S(self_sf7[1346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1347]),
        .S(self_sf7[1347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1348]),
        .S(self_sf7[1348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1349]),
        .S(self_sf7[1349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[134]),
        .S(self_sf7[134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1350]),
        .S(self_sf7[1350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1351]),
        .S(self_sf7[1351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1352]),
        .S(self_sf7[1352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1353]),
        .S(self_sf7[1353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1354]),
        .S(self_sf7[1354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1355]),
        .S(self_sf7[1355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1356]),
        .S(self_sf7[1356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1357]),
        .S(self_sf7[1357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1358]),
        .S(self_sf7[1358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1359]),
        .S(self_sf7[1359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[135]),
        .S(self_sf7[135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1360]),
        .S(self_sf7[1360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1361]),
        .S(self_sf7[1361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1362]),
        .S(self_sf7[1362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1363]),
        .S(self_sf7[1363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1364]),
        .S(self_sf7[1364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1365]),
        .S(self_sf7[1365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1366]),
        .S(self_sf7[1366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1367]),
        .S(self_sf7[1367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1368]),
        .S(self_sf7[1368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1369]),
        .S(self_sf7[1369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[136]),
        .S(self_sf7[136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1370]),
        .S(self_sf7[1370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1371]),
        .S(self_sf7[1371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1372]),
        .S(self_sf7[1372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1373]),
        .S(self_sf7[1373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1374]),
        .S(self_sf7[1374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1375]),
        .S(self_sf7[1375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1376]),
        .S(self_sf7[1376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1377]),
        .S(self_sf7[1377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1378]),
        .S(self_sf7[1378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1379]),
        .S(self_sf7[1379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[137]),
        .S(self_sf7[137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1380]),
        .S(self_sf7[1380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1381]),
        .S(self_sf7[1381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1382]),
        .S(self_sf7[1382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1383]),
        .S(self_sf7[1383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1384]),
        .S(self_sf7[1384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1385]),
        .S(self_sf7[1385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1386]),
        .S(self_sf7[1386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1387]),
        .S(self_sf7[1387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1388]),
        .S(self_sf7[1388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1389]),
        .S(self_sf7[1389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[138]),
        .S(self_sf7[138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1390]),
        .S(self_sf7[1390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1391]),
        .S(self_sf7[1391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1392]),
        .S(self_sf7[1392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1393]),
        .S(self_sf7[1393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1394]),
        .S(self_sf7[1394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1395]),
        .S(self_sf7[1395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1396]),
        .S(self_sf7[1396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1397]),
        .S(self_sf7[1397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1398]),
        .S(self_sf7[1398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1399]),
        .S(self_sf7[1399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[139]),
        .S(self_sf7[139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[13].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[13]),
        .S(self_sf7[13]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1400]),
        .S(self_sf7[1400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1401]),
        .S(self_sf7[1401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1402]),
        .S(self_sf7[1402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1403]),
        .S(self_sf7[1403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1404]),
        .S(self_sf7[1404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1405]),
        .S(self_sf7[1405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1406]),
        .S(self_sf7[1406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1407]),
        .S(self_sf7[1407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1408]),
        .S(self_sf7[1408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1409]),
        .S(self_sf7[1409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[140]),
        .S(self_sf7[140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1410]),
        .S(self_sf7[1410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1411]),
        .S(self_sf7[1411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1412]),
        .S(self_sf7[1412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1413]),
        .S(self_sf7[1413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1414]),
        .S(self_sf7[1414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1415]),
        .S(self_sf7[1415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1416]),
        .S(self_sf7[1416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1417]),
        .S(self_sf7[1417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1418]),
        .S(self_sf7[1418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1419]),
        .S(self_sf7[1419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[141]),
        .S(self_sf7[141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1420]),
        .S(self_sf7[1420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1421]),
        .S(self_sf7[1421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1422]),
        .S(self_sf7[1422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1423]),
        .S(self_sf7[1423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1424]),
        .S(self_sf7[1424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1425]),
        .S(self_sf7[1425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1426]),
        .S(self_sf7[1426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1427]),
        .S(self_sf7[1427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1428]),
        .S(self_sf7[1428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1429]),
        .S(self_sf7[1429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[142]),
        .S(self_sf7[142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1430]),
        .S(self_sf7[1430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1431]),
        .S(self_sf7[1431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1432]),
        .S(self_sf7[1432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1433]),
        .S(self_sf7[1433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1434]),
        .S(self_sf7[1434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1435]),
        .S(self_sf7[1435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1436]),
        .S(self_sf7[1436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1437]),
        .S(self_sf7[1437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1438]),
        .S(self_sf7[1438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1439]),
        .S(self_sf7[1439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[143]),
        .S(self_sf7[143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1440]),
        .S(self_sf7[1440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1441]),
        .S(self_sf7[1441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1442]),
        .S(self_sf7[1442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1443]),
        .S(self_sf7[1443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1444]),
        .S(self_sf7[1444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1445]),
        .S(self_sf7[1445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1446]),
        .S(self_sf7[1446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1447]),
        .S(self_sf7[1447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1448]),
        .S(self_sf7[1448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1449]),
        .S(self_sf7[1449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[144]),
        .S(self_sf7[144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1450]),
        .S(self_sf7[1450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1451]),
        .S(self_sf7[1451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1452]),
        .S(self_sf7[1452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1453]),
        .S(self_sf7[1453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1454]),
        .S(self_sf7[1454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1455]),
        .S(self_sf7[1455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1456]),
        .S(self_sf7[1456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1457]),
        .S(self_sf7[1457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1458]),
        .S(self_sf7[1458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1459]),
        .S(self_sf7[1459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[145]),
        .S(self_sf7[145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1460]),
        .S(self_sf7[1460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1461]),
        .S(self_sf7[1461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1462]),
        .S(self_sf7[1462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1463]),
        .S(self_sf7[1463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1464]),
        .S(self_sf7[1464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1465]),
        .S(self_sf7[1465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1466]),
        .S(self_sf7[1466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1467]),
        .S(self_sf7[1467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1468]),
        .S(self_sf7[1468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1469]),
        .S(self_sf7[1469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[146]),
        .S(self_sf7[146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1470]),
        .S(self_sf7[1470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1471]),
        .S(self_sf7[1471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1472]),
        .S(self_sf7[1472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1473]),
        .S(self_sf7[1473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1474]),
        .S(self_sf7[1474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1475]),
        .S(self_sf7[1475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1476]),
        .S(self_sf7[1476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1477]),
        .S(self_sf7[1477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1478]),
        .S(self_sf7[1478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1479]),
        .S(self_sf7[1479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[147]),
        .S(self_sf7[147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1480]),
        .S(self_sf7[1480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1481]),
        .S(self_sf7[1481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1482]),
        .S(self_sf7[1482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1483]),
        .S(self_sf7[1483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1484]),
        .S(self_sf7[1484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1485]),
        .S(self_sf7[1485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1486]),
        .S(self_sf7[1486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1487]),
        .S(self_sf7[1487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1488]),
        .S(self_sf7[1488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1489]),
        .S(self_sf7[1489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[148]),
        .S(self_sf7[148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1490]),
        .S(self_sf7[1490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1491]),
        .S(self_sf7[1491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1492]),
        .S(self_sf7[1492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1493]),
        .S(self_sf7[1493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1494]),
        .S(self_sf7[1494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1495]),
        .S(self_sf7[1495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1496]),
        .S(self_sf7[1496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1497]),
        .S(self_sf7[1497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1498]),
        .S(self_sf7[1498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1499]),
        .S(self_sf7[1499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[149]),
        .S(self_sf7[149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[14].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[14]),
        .S(self_sf7[14]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1500]),
        .S(self_sf7[1500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1501]),
        .S(self_sf7[1501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1502]),
        .S(self_sf7[1502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1503]),
        .S(self_sf7[1503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1504]),
        .S(self_sf7[1504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1505]),
        .S(self_sf7[1505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1506]),
        .S(self_sf7[1506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1507]),
        .S(self_sf7[1507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1508]),
        .S(self_sf7[1508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1509]),
        .S(self_sf7[1509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[150]),
        .S(self_sf7[150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1510]),
        .S(self_sf7[1510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1511]),
        .S(self_sf7[1511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1512]),
        .S(self_sf7[1512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1513]),
        .S(self_sf7[1513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1514]),
        .S(self_sf7[1514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1515]),
        .S(self_sf7[1515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1516]),
        .S(self_sf7[1516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1517]),
        .S(self_sf7[1517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1518]),
        .S(self_sf7[1518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1519]),
        .S(self_sf7[1519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[151]),
        .S(self_sf7[151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1520]),
        .S(self_sf7[1520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1521]),
        .S(self_sf7[1521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1522]),
        .S(self_sf7[1522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1523]),
        .S(self_sf7[1523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1524]),
        .S(self_sf7[1524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1525]),
        .S(self_sf7[1525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1526]),
        .S(self_sf7[1526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1527]),
        .S(self_sf7[1527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1528]),
        .S(self_sf7[1528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1529]),
        .S(self_sf7[1529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[152]),
        .S(self_sf7[152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1530]),
        .S(self_sf7[1530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1531]),
        .S(self_sf7[1531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1532]),
        .S(self_sf7[1532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1533]),
        .S(self_sf7[1533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1534]),
        .S(self_sf7[1534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1535]),
        .S(self_sf7[1535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1536]),
        .S(self_sf7[1536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1537]),
        .S(self_sf7[1537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1538]),
        .S(self_sf7[1538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1539]),
        .S(self_sf7[1539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[153]),
        .S(self_sf7[153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1540]),
        .S(self_sf7[1540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1541]),
        .S(self_sf7[1541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1542]),
        .S(self_sf7[1542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1543]),
        .S(self_sf7[1543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1544]),
        .S(self_sf7[1544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1545]),
        .S(self_sf7[1545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1546]),
        .S(self_sf7[1546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1547]),
        .S(self_sf7[1547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1548]),
        .S(self_sf7[1548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1549]),
        .S(self_sf7[1549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[154]),
        .S(self_sf7[154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1550]),
        .S(self_sf7[1550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1551]),
        .S(self_sf7[1551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1552]),
        .S(self_sf7[1552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1553]),
        .S(self_sf7[1553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1554]),
        .S(self_sf7[1554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1555]),
        .S(self_sf7[1555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1556]),
        .S(self_sf7[1556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1557]),
        .S(self_sf7[1557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1558]),
        .S(self_sf7[1558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1559]),
        .S(self_sf7[1559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[155]),
        .S(self_sf7[155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1560]),
        .S(self_sf7[1560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1561]),
        .S(self_sf7[1561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1562]),
        .S(self_sf7[1562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1563]),
        .S(self_sf7[1563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1564]),
        .S(self_sf7[1564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1565]),
        .S(self_sf7[1565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1566]),
        .S(self_sf7[1566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1567]),
        .S(self_sf7[1567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1568]),
        .S(self_sf7[1568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1569]),
        .S(self_sf7[1569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[156]),
        .S(self_sf7[156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1570]),
        .S(self_sf7[1570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1571]),
        .S(self_sf7[1571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1572]),
        .S(self_sf7[1572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1573]),
        .S(self_sf7[1573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1574]),
        .S(self_sf7[1574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1575]),
        .S(self_sf7[1575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1576]),
        .S(self_sf7[1576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1577]),
        .S(self_sf7[1577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1578]),
        .S(self_sf7[1578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1579]),
        .S(self_sf7[1579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[157]),
        .S(self_sf7[157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1580]),
        .S(self_sf7[1580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1581]),
        .S(self_sf7[1581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1582]),
        .S(self_sf7[1582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1583]),
        .S(self_sf7[1583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1584]),
        .S(self_sf7[1584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1585]),
        .S(self_sf7[1585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1586]),
        .S(self_sf7[1586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1587]),
        .S(self_sf7[1587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1588]),
        .S(self_sf7[1588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1589]),
        .S(self_sf7[1589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[158]),
        .S(self_sf7[158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1590]),
        .S(self_sf7[1590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1591]),
        .S(self_sf7[1591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1592]),
        .S(self_sf7[1592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1593]),
        .S(self_sf7[1593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1594]),
        .S(self_sf7[1594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1595]),
        .S(self_sf7[1595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1596]),
        .S(self_sf7[1596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1597]),
        .S(self_sf7[1597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1598]),
        .S(self_sf7[1598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1599]),
        .S(self_sf7[1599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[159]),
        .S(self_sf7[159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[15].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[15]),
        .S(self_sf7[15]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1600]),
        .S(self_sf7[1600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1601]),
        .S(self_sf7[1601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1602]),
        .S(self_sf7[1602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1603]),
        .S(self_sf7[1603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1604]),
        .S(self_sf7[1604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1605]),
        .S(self_sf7[1605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1606]),
        .S(self_sf7[1606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1607]),
        .S(self_sf7[1607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1608]),
        .S(self_sf7[1608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1609]),
        .S(self_sf7[1609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[160]),
        .S(self_sf7[160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1610]),
        .S(self_sf7[1610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1611]),
        .S(self_sf7[1611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1612]),
        .S(self_sf7[1612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1613]),
        .S(self_sf7[1613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1614]),
        .S(self_sf7[1614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1615]),
        .S(self_sf7[1615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1616]),
        .S(self_sf7[1616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1617]),
        .S(self_sf7[1617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1618]),
        .S(self_sf7[1618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1619]),
        .S(self_sf7[1619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[161]),
        .S(self_sf7[161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1620]),
        .S(self_sf7[1620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1621]),
        .S(self_sf7[1621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1622]),
        .S(self_sf7[1622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1623]),
        .S(self_sf7[1623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1624]),
        .S(self_sf7[1624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1625]),
        .S(self_sf7[1625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1626]),
        .S(self_sf7[1626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1627]),
        .S(self_sf7[1627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1628]),
        .S(self_sf7[1628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1629]),
        .S(self_sf7[1629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[162]),
        .S(self_sf7[162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1630]),
        .S(self_sf7[1630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1631]),
        .S(self_sf7[1631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1632]),
        .S(self_sf7[1632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1633]),
        .S(self_sf7[1633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1634]),
        .S(self_sf7[1634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1635]),
        .S(self_sf7[1635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1636]),
        .S(self_sf7[1636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1637]),
        .S(self_sf7[1637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1638]),
        .S(self_sf7[1638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1639]),
        .S(self_sf7[1639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[163]),
        .S(self_sf7[163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1640]),
        .S(self_sf7[1640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1641]),
        .S(self_sf7[1641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1642]),
        .S(self_sf7[1642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1643]),
        .S(self_sf7[1643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1644]),
        .S(self_sf7[1644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1645]),
        .S(self_sf7[1645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1646]),
        .S(self_sf7[1646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1647]),
        .S(self_sf7[1647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1648]),
        .S(self_sf7[1648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1649]),
        .S(self_sf7[1649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[164]),
        .S(self_sf7[164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1650]),
        .S(self_sf7[1650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1651]),
        .S(self_sf7[1651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1652]),
        .S(self_sf7[1652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1653]),
        .S(self_sf7[1653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1654]),
        .S(self_sf7[1654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1655]),
        .S(self_sf7[1655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1656]),
        .S(self_sf7[1656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1657]),
        .S(self_sf7[1657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1658]),
        .S(self_sf7[1658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1659]),
        .S(self_sf7[1659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[165]),
        .S(self_sf7[165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1660]),
        .S(self_sf7[1660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1661]),
        .S(self_sf7[1661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1662]),
        .S(self_sf7[1662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1663]),
        .S(self_sf7[1663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1664]),
        .S(self_sf7[1664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1665]),
        .S(self_sf7[1665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1666]),
        .S(self_sf7[1666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1667]),
        .S(self_sf7[1667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1668]),
        .S(self_sf7[1668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1669]),
        .S(self_sf7[1669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[166]),
        .S(self_sf7[166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1670]),
        .S(self_sf7[1670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1671]),
        .S(self_sf7[1671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1672]),
        .S(self_sf7[1672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1673]),
        .S(self_sf7[1673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1674]),
        .S(self_sf7[1674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1675]),
        .S(self_sf7[1675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1676]),
        .S(self_sf7[1676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1677]),
        .S(self_sf7[1677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1678]),
        .S(self_sf7[1678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1679]),
        .S(self_sf7[1679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[167]),
        .S(self_sf7[167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1680]),
        .S(self_sf7[1680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1681]),
        .S(self_sf7[1681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1682]),
        .S(self_sf7[1682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1683]),
        .S(self_sf7[1683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1684]),
        .S(self_sf7[1684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1685]),
        .S(self_sf7[1685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1686]),
        .S(self_sf7[1686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1687]),
        .S(self_sf7[1687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1688]),
        .S(self_sf7[1688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1689]),
        .S(self_sf7[1689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[168]),
        .S(self_sf7[168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1690]),
        .S(self_sf7[1690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1691]),
        .S(self_sf7[1691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1692]),
        .S(self_sf7[1692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1693]),
        .S(self_sf7[1693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1694]),
        .S(self_sf7[1694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1695]),
        .S(self_sf7[1695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1696]),
        .S(self_sf7[1696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1697]),
        .S(self_sf7[1697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1698]),
        .S(self_sf7[1698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1699]),
        .S(self_sf7[1699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[169]),
        .S(self_sf7[169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[16].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[16]),
        .S(self_sf7[16]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1700]),
        .S(self_sf7[1700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1701]),
        .S(self_sf7[1701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1702]),
        .S(self_sf7[1702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1703]),
        .S(self_sf7[1703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1704]),
        .S(self_sf7[1704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1705]),
        .S(self_sf7[1705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1706]),
        .S(self_sf7[1706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1707]),
        .S(self_sf7[1707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1708]),
        .S(self_sf7[1708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1709]),
        .S(self_sf7[1709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[170]),
        .S(self_sf7[170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1710]),
        .S(self_sf7[1710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1711]),
        .S(self_sf7[1711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1712]),
        .S(self_sf7[1712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1713]),
        .S(self_sf7[1713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1714]),
        .S(self_sf7[1714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1715]),
        .S(self_sf7[1715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1716]),
        .S(self_sf7[1716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1717]),
        .S(self_sf7[1717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1718]),
        .S(self_sf7[1718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1719]),
        .S(self_sf7[1719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[171]),
        .S(self_sf7[171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1720]),
        .S(self_sf7[1720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1721]),
        .S(self_sf7[1721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1722]),
        .S(self_sf7[1722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1723]),
        .S(self_sf7[1723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1724]),
        .S(self_sf7[1724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1725]),
        .S(self_sf7[1725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1726]),
        .S(self_sf7[1726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1727]),
        .S(self_sf7[1727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1728]),
        .S(self_sf7[1728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1729]),
        .S(self_sf7[1729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[172]),
        .S(self_sf7[172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1730]),
        .S(self_sf7[1730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1731]),
        .S(self_sf7[1731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1732]),
        .S(self_sf7[1732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1733]),
        .S(self_sf7[1733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1734]),
        .S(self_sf7[1734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1735]),
        .S(self_sf7[1735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1736]),
        .S(self_sf7[1736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1737]),
        .S(self_sf7[1737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1738]),
        .S(self_sf7[1738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1739]),
        .S(self_sf7[1739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[173]),
        .S(self_sf7[173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1740]),
        .S(self_sf7[1740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1741]),
        .S(self_sf7[1741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1742]),
        .S(self_sf7[1742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1743]),
        .S(self_sf7[1743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1744]),
        .S(self_sf7[1744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1745]),
        .S(self_sf7[1745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1746]),
        .S(self_sf7[1746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1747]),
        .S(self_sf7[1747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1748]),
        .S(self_sf7[1748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1749]),
        .S(self_sf7[1749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[174]),
        .S(self_sf7[174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1750]),
        .S(self_sf7[1750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1751]),
        .S(self_sf7[1751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1752]),
        .S(self_sf7[1752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1753]),
        .S(self_sf7[1753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1754]),
        .S(self_sf7[1754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1755]),
        .S(self_sf7[1755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1756]),
        .S(self_sf7[1756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1757]),
        .S(self_sf7[1757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1758]),
        .S(self_sf7[1758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1759]),
        .S(self_sf7[1759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[175]),
        .S(self_sf7[175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1760]),
        .S(self_sf7[1760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1761]),
        .S(self_sf7[1761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1762]),
        .S(self_sf7[1762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1763]),
        .S(self_sf7[1763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1764]),
        .S(self_sf7[1764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1765]),
        .S(self_sf7[1765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1766]),
        .S(self_sf7[1766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1767]),
        .S(self_sf7[1767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1768]),
        .S(self_sf7[1768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1769]),
        .S(self_sf7[1769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[176]),
        .S(self_sf7[176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1770]),
        .S(self_sf7[1770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1771]),
        .S(self_sf7[1771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1772]),
        .S(self_sf7[1772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1773]),
        .S(self_sf7[1773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1774]),
        .S(self_sf7[1774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1775]),
        .S(self_sf7[1775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1776]),
        .S(self_sf7[1776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1777]),
        .S(self_sf7[1777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1778]),
        .S(self_sf7[1778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1779]),
        .S(self_sf7[1779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[177]),
        .S(self_sf7[177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1780]),
        .S(self_sf7[1780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1781]),
        .S(self_sf7[1781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1782]),
        .S(self_sf7[1782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1783]),
        .S(self_sf7[1783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1784]),
        .S(self_sf7[1784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1785]),
        .S(self_sf7[1785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1786]),
        .S(self_sf7[1786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1787]),
        .S(self_sf7[1787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1788]),
        .S(self_sf7[1788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1789]),
        .S(self_sf7[1789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[178]),
        .S(self_sf7[178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1790]),
        .S(self_sf7[1790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1791]),
        .S(self_sf7[1791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1792]),
        .S(self_sf7[1792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1793]),
        .S(self_sf7[1793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1794]),
        .S(self_sf7[1794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1795]),
        .S(self_sf7[1795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1796]),
        .S(self_sf7[1796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1797]),
        .S(self_sf7[1797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1798]),
        .S(self_sf7[1798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1799]),
        .S(self_sf7[1799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[179]),
        .S(self_sf7[179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[17].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[17]),
        .S(self_sf7[17]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[180]),
        .S(self_sf7[180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[181]),
        .S(self_sf7[181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[182]),
        .S(self_sf7[182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[183]),
        .S(self_sf7[183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[184]),
        .S(self_sf7[184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[185]),
        .S(self_sf7[185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[186]),
        .S(self_sf7[186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[187]),
        .S(self_sf7[187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[188]),
        .S(self_sf7[188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[189]),
        .S(self_sf7[189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[18].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[18]),
        .S(self_sf7[18]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[190]),
        .S(self_sf7[190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[191]),
        .S(self_sf7[191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[192]),
        .S(self_sf7[192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[193]),
        .S(self_sf7[193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[194]),
        .S(self_sf7[194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[195]),
        .S(self_sf7[195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[196]),
        .S(self_sf7[196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[197]),
        .S(self_sf7[197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[198]),
        .S(self_sf7[198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[199]),
        .S(self_sf7[199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[19].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[19]),
        .S(self_sf7[19]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1]),
        .S(info_sf7[1]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[200]),
        .S(self_sf7[200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[201]),
        .S(self_sf7[201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[202]),
        .S(self_sf7[202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[203]),
        .S(self_sf7[203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[204]),
        .S(self_sf7[204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[205]),
        .S(self_sf7[205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[206]),
        .S(self_sf7[206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[207]),
        .S(self_sf7[207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[208]),
        .S(self_sf7[208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[209]),
        .S(self_sf7[209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[20].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[20]),
        .S(self_sf7[20]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[210]),
        .S(self_sf7[210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[211]),
        .S(self_sf7[211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[212]),
        .S(self_sf7[212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[213]),
        .S(self_sf7[213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[214]),
        .S(self_sf7[214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[215]),
        .S(self_sf7[215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[216]),
        .S(self_sf7[216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[217]),
        .S(self_sf7[217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[218]),
        .S(self_sf7[218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[219]),
        .S(self_sf7[219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[21].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[21]),
        .S(self_sf7[21]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[220]),
        .S(self_sf7[220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[221]),
        .S(self_sf7[221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[222]),
        .S(self_sf7[222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[223]),
        .S(self_sf7[223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[224]),
        .S(self_sf7[224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[225]),
        .S(self_sf7[225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[226]),
        .S(self_sf7[226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[227]),
        .S(self_sf7[227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[228]),
        .S(self_sf7[228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[229]),
        .S(self_sf7[229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[22].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[22]),
        .S(self_sf7[22]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[230]),
        .S(self_sf7[230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[231]),
        .S(self_sf7[231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[232]),
        .S(self_sf7[232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[233]),
        .S(self_sf7[233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[234]),
        .S(self_sf7[234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[235]),
        .S(self_sf7[235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[236]),
        .S(self_sf7[236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[237]),
        .S(self_sf7[237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[238]),
        .S(self_sf7[238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[239]),
        .S(self_sf7[239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[23].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[23]),
        .S(self_sf7[23]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[240]),
        .S(self_sf7[240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[241]),
        .S(self_sf7[241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[242]),
        .S(self_sf7[242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[243]),
        .S(self_sf7[243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[244]),
        .S(self_sf7[244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[245]),
        .S(self_sf7[245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[246]),
        .S(self_sf7[246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[247]),
        .S(self_sf7[247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[248]),
        .S(self_sf7[248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[249]),
        .S(self_sf7[249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[24].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[24]),
        .S(self_sf7[24]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[250]),
        .S(self_sf7[250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[251]),
        .S(self_sf7[251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[252]),
        .S(self_sf7[252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[253]),
        .S(self_sf7[253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[254]),
        .S(self_sf7[254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[255]),
        .S(self_sf7[255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[256]),
        .S(self_sf7[256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[257]),
        .S(self_sf7[257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[258]),
        .S(self_sf7[258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[259]),
        .S(self_sf7[259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[25].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[25]),
        .S(self_sf7[25]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[260]),
        .S(self_sf7[260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[261]),
        .S(self_sf7[261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[262]),
        .S(self_sf7[262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[263]),
        .S(self_sf7[263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[264]),
        .S(self_sf7[264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[265]),
        .S(self_sf7[265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[266]),
        .S(self_sf7[266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[267]),
        .S(self_sf7[267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[268]),
        .S(self_sf7[268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[269]),
        .S(self_sf7[269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[26].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[26]),
        .S(self_sf7[26]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[270]),
        .S(self_sf7[270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[271]),
        .S(self_sf7[271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[272]),
        .S(self_sf7[272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[273]),
        .S(self_sf7[273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[274]),
        .S(self_sf7[274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[275]),
        .S(self_sf7[275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[276]),
        .S(self_sf7[276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[277]),
        .S(self_sf7[277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[278]),
        .S(self_sf7[278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[279]),
        .S(self_sf7[279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[27].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[27]),
        .S(self_sf7[27]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[280]),
        .S(self_sf7[280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[281]),
        .S(self_sf7[281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[282]),
        .S(self_sf7[282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[283]),
        .S(self_sf7[283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[284]),
        .S(self_sf7[284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[285]),
        .S(self_sf7[285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[286]),
        .S(self_sf7[286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[287]),
        .S(self_sf7[287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[288]),
        .S(self_sf7[288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[289]),
        .S(self_sf7[289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[28].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[28]),
        .S(self_sf7[28]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[290]),
        .S(self_sf7[290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[291]),
        .S(self_sf7[291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[292]),
        .S(self_sf7[292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[293]),
        .S(self_sf7[293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[294]),
        .S(self_sf7[294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[295]),
        .S(self_sf7[295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[296]),
        .S(self_sf7[296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[297]),
        .S(self_sf7[297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[298]),
        .S(self_sf7[298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[299]),
        .S(self_sf7[299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[29].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[29]),
        .S(self_sf7[29]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[2].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[2]),
        .S(info_sf7[2]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[300]),
        .S(self_sf7[300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[301]),
        .S(self_sf7[301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[302]),
        .S(self_sf7[302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[303]),
        .S(self_sf7[303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[304]),
        .S(self_sf7[304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[305]),
        .S(self_sf7[305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[306]),
        .S(self_sf7[306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[307]),
        .S(self_sf7[307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[308]),
        .S(self_sf7[308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[309]),
        .S(self_sf7[309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[30].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[30]),
        .S(self_sf7[30]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[310]),
        .S(self_sf7[310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[311]),
        .S(self_sf7[311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[312]),
        .S(self_sf7[312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[313]),
        .S(self_sf7[313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[314]),
        .S(self_sf7[314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[315]),
        .S(self_sf7[315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[316]),
        .S(self_sf7[316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[317]),
        .S(self_sf7[317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[318]),
        .S(self_sf7[318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[319]),
        .S(self_sf7[319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[31].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[31]),
        .S(self_sf7[31]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[320]),
        .S(self_sf7[320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[321]),
        .S(self_sf7[321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[322]),
        .S(self_sf7[322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[323]),
        .S(self_sf7[323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[324]),
        .S(self_sf7[324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[325]),
        .S(self_sf7[325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[326]),
        .S(self_sf7[326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[327]),
        .S(self_sf7[327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[328]),
        .S(self_sf7[328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[329]),
        .S(self_sf7[329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[32].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[32]),
        .S(self_sf7[32]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[330]),
        .S(self_sf7[330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[331]),
        .S(self_sf7[331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[332]),
        .S(self_sf7[332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[333]),
        .S(self_sf7[333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[334]),
        .S(self_sf7[334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[335]),
        .S(self_sf7[335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[336]),
        .S(self_sf7[336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[337]),
        .S(self_sf7[337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[338]),
        .S(self_sf7[338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[339]),
        .S(self_sf7[339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[33].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[33]),
        .S(self_sf7[33]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[340]),
        .S(self_sf7[340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[341]),
        .S(self_sf7[341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[342]),
        .S(self_sf7[342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[343]),
        .S(self_sf7[343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[344]),
        .S(self_sf7[344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[345]),
        .S(self_sf7[345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[346]),
        .S(self_sf7[346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[347]),
        .S(self_sf7[347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[348]),
        .S(self_sf7[348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[349]),
        .S(self_sf7[349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[34].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[34]),
        .S(self_sf7[34]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[350]),
        .S(self_sf7[350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[351]),
        .S(self_sf7[351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[352]),
        .S(self_sf7[352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[353]),
        .S(self_sf7[353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[354]),
        .S(self_sf7[354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[355]),
        .S(self_sf7[355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[356]),
        .S(self_sf7[356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[357]),
        .S(self_sf7[357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[358]),
        .S(self_sf7[358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[359]),
        .S(self_sf7[359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[35].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[35]),
        .S(self_sf7[35]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[360]),
        .S(self_sf7[360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[361]),
        .S(self_sf7[361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[362]),
        .S(self_sf7[362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[363]),
        .S(self_sf7[363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[364]),
        .S(self_sf7[364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[365]),
        .S(self_sf7[365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[366]),
        .S(self_sf7[366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[367]),
        .S(self_sf7[367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[368]),
        .S(self_sf7[368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[369]),
        .S(self_sf7[369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[36].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[36]),
        .S(self_sf7[36]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[370]),
        .S(self_sf7[370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[371]),
        .S(self_sf7[371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[372]),
        .S(self_sf7[372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[373]),
        .S(self_sf7[373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[374]),
        .S(self_sf7[374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[375]),
        .S(self_sf7[375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[376]),
        .S(self_sf7[376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[377]),
        .S(self_sf7[377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[378]),
        .S(self_sf7[378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[379]),
        .S(self_sf7[379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[37].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[37]),
        .S(self_sf7[37]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[380]),
        .S(self_sf7[380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[381]),
        .S(self_sf7[381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[382]),
        .S(self_sf7[382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[383]),
        .S(self_sf7[383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[384]),
        .S(self_sf7[384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[385]),
        .S(self_sf7[385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[386]),
        .S(self_sf7[386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[387]),
        .S(self_sf7[387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[388]),
        .S(self_sf7[388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[389]),
        .S(self_sf7[389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[38].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[38]),
        .S(self_sf7[38]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[390]),
        .S(self_sf7[390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[391]),
        .S(self_sf7[391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[392]),
        .S(self_sf7[392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[393]),
        .S(self_sf7[393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[394]),
        .S(self_sf7[394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[395]),
        .S(self_sf7[395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[396]),
        .S(self_sf7[396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[397]),
        .S(self_sf7[397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[398]),
        .S(self_sf7[398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[399]),
        .S(self_sf7[399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[39].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[39]),
        .S(self_sf7[39]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[3].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[3]),
        .S(info_sf7[3]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[400]),
        .S(self_sf7[400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[401]),
        .S(self_sf7[401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[402]),
        .S(self_sf7[402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[403]),
        .S(self_sf7[403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[404]),
        .S(self_sf7[404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[405]),
        .S(self_sf7[405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[406]),
        .S(self_sf7[406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[407]),
        .S(self_sf7[407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[408]),
        .S(self_sf7[408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[409]),
        .S(self_sf7[409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[40].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[40]),
        .S(self_sf7[40]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[410]),
        .S(self_sf7[410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[411]),
        .S(self_sf7[411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[412]),
        .S(self_sf7[412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[413]),
        .S(self_sf7[413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[414]),
        .S(self_sf7[414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[415]),
        .S(self_sf7[415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[416]),
        .S(self_sf7[416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[417]),
        .S(self_sf7[417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[418]),
        .S(self_sf7[418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[419]),
        .S(self_sf7[419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[41].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[41]),
        .S(self_sf7[41]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[420]),
        .S(self_sf7[420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[421]),
        .S(self_sf7[421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[422]),
        .S(self_sf7[422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[423]),
        .S(self_sf7[423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[424]),
        .S(self_sf7[424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[425]),
        .S(self_sf7[425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[426]),
        .S(self_sf7[426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[427]),
        .S(self_sf7[427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[428]),
        .S(self_sf7[428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[429]),
        .S(self_sf7[429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[42].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[42]),
        .S(self_sf7[42]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[430]),
        .S(self_sf7[430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[431]),
        .S(self_sf7[431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[432]),
        .S(self_sf7[432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[433]),
        .S(self_sf7[433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[434]),
        .S(self_sf7[434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[435]),
        .S(self_sf7[435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[436]),
        .S(self_sf7[436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[437]),
        .S(self_sf7[437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[438]),
        .S(self_sf7[438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[439]),
        .S(self_sf7[439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[43].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[43]),
        .S(self_sf7[43]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[440]),
        .S(self_sf7[440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[441]),
        .S(self_sf7[441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[442]),
        .S(self_sf7[442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[443]),
        .S(self_sf7[443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[444]),
        .S(self_sf7[444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[445]),
        .S(self_sf7[445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[446]),
        .S(self_sf7[446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[447]),
        .S(self_sf7[447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[448]),
        .S(self_sf7[448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[449]),
        .S(self_sf7[449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[44].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[44]),
        .S(self_sf7[44]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[450]),
        .S(self_sf7[450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[451]),
        .S(self_sf7[451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[452]),
        .S(self_sf7[452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[453]),
        .S(self_sf7[453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[454]),
        .S(self_sf7[454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[455]),
        .S(self_sf7[455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[456]),
        .S(self_sf7[456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[457]),
        .S(self_sf7[457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[458]),
        .S(self_sf7[458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[459]),
        .S(self_sf7[459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[45].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[45]),
        .S(self_sf7[45]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[460]),
        .S(self_sf7[460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[461]),
        .S(self_sf7[461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[462]),
        .S(self_sf7[462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[463]),
        .S(self_sf7[463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[464]),
        .S(self_sf7[464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[465]),
        .S(self_sf7[465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[466]),
        .S(self_sf7[466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[467]),
        .S(self_sf7[467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[468]),
        .S(self_sf7[468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[469]),
        .S(self_sf7[469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[46].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[46]),
        .S(self_sf7[46]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[470]),
        .S(self_sf7[470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[471]),
        .S(self_sf7[471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[472]),
        .S(self_sf7[472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[473]),
        .S(self_sf7[473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[474]),
        .S(self_sf7[474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[475]),
        .S(self_sf7[475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[476]),
        .S(self_sf7[476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[477]),
        .S(self_sf7[477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[478]),
        .S(self_sf7[478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[479]),
        .S(self_sf7[479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[47].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[47]),
        .S(self_sf7[47]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[480]),
        .S(self_sf7[480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[481]),
        .S(self_sf7[481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[482]),
        .S(self_sf7[482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[483]),
        .S(self_sf7[483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[484]),
        .S(self_sf7[484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[485]),
        .S(self_sf7[485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[486]),
        .S(self_sf7[486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[487]),
        .S(self_sf7[487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[488]),
        .S(self_sf7[488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[489]),
        .S(self_sf7[489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[48].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[48]),
        .S(self_sf7[48]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[490]),
        .S(self_sf7[490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[491]),
        .S(self_sf7[491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[492]),
        .S(self_sf7[492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[493]),
        .S(self_sf7[493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[494]),
        .S(self_sf7[494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[495]),
        .S(self_sf7[495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[496]),
        .S(self_sf7[496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[497]),
        .S(self_sf7[497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[498]),
        .S(self_sf7[498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[499]),
        .S(self_sf7[499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[49].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[49]),
        .S(self_sf7[49]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[4].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[4]),
        .S(info_sf7[4]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[500]),
        .S(self_sf7[500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[501]),
        .S(self_sf7[501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[502]),
        .S(self_sf7[502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[503]),
        .S(self_sf7[503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[504]),
        .S(self_sf7[504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[505]),
        .S(self_sf7[505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[506]),
        .S(self_sf7[506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[507]),
        .S(self_sf7[507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[508]),
        .S(self_sf7[508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[509]),
        .S(self_sf7[509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[50].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[50]),
        .S(self_sf7[50]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[510]),
        .S(self_sf7[510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[511]),
        .S(self_sf7[511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[512]),
        .S(self_sf7[512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[513]),
        .S(self_sf7[513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[514]),
        .S(self_sf7[514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[515]),
        .S(self_sf7[515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[516]),
        .S(self_sf7[516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[517]),
        .S(self_sf7[517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[518]),
        .S(self_sf7[518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[519]),
        .S(self_sf7[519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[51].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[51]),
        .S(self_sf7[51]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[520]),
        .S(self_sf7[520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[521]),
        .S(self_sf7[521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[522]),
        .S(self_sf7[522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[523]),
        .S(self_sf7[523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[524]),
        .S(self_sf7[524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[525]),
        .S(self_sf7[525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[526]),
        .S(self_sf7[526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[527]),
        .S(self_sf7[527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[528]),
        .S(self_sf7[528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[529]),
        .S(self_sf7[529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[52].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[52]),
        .S(self_sf7[52]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[530]),
        .S(self_sf7[530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[531]),
        .S(self_sf7[531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[532]),
        .S(self_sf7[532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[533]),
        .S(self_sf7[533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[534]),
        .S(self_sf7[534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[535]),
        .S(self_sf7[535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[536]),
        .S(self_sf7[536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[537]),
        .S(self_sf7[537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[538]),
        .S(self_sf7[538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[539]),
        .S(self_sf7[539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[53].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[53]),
        .S(self_sf7[53]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[540]),
        .S(self_sf7[540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[541]),
        .S(self_sf7[541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[542]),
        .S(self_sf7[542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[543]),
        .S(self_sf7[543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[544]),
        .S(self_sf7[544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[545]),
        .S(self_sf7[545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[546]),
        .S(self_sf7[546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[547]),
        .S(self_sf7[547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[548]),
        .S(self_sf7[548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[549]),
        .S(self_sf7[549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[54].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[54]),
        .S(self_sf7[54]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[550]),
        .S(self_sf7[550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[551]),
        .S(self_sf7[551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[552]),
        .S(self_sf7[552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[553]),
        .S(self_sf7[553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[554]),
        .S(self_sf7[554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[555]),
        .S(self_sf7[555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[556]),
        .S(self_sf7[556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[557]),
        .S(self_sf7[557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[558]),
        .S(self_sf7[558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[559]),
        .S(self_sf7[559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[55].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[55]),
        .S(self_sf7[55]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[560]),
        .S(self_sf7[560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[561]),
        .S(self_sf7[561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[562]),
        .S(self_sf7[562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[563]),
        .S(self_sf7[563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[564]),
        .S(self_sf7[564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[565]),
        .S(self_sf7[565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[566]),
        .S(self_sf7[566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[567]),
        .S(self_sf7[567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[568]),
        .S(self_sf7[568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[569]),
        .S(self_sf7[569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[56].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[56]),
        .S(self_sf7[56]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[570]),
        .S(self_sf7[570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[571]),
        .S(self_sf7[571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[572]),
        .S(self_sf7[572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[573]),
        .S(self_sf7[573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[574]),
        .S(self_sf7[574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[575]),
        .S(self_sf7[575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[576]),
        .S(self_sf7[576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[577]),
        .S(self_sf7[577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[578]),
        .S(self_sf7[578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[579]),
        .S(self_sf7[579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[57].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[57]),
        .S(self_sf7[57]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[580]),
        .S(self_sf7[580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[581]),
        .S(self_sf7[581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[582]),
        .S(self_sf7[582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[583]),
        .S(self_sf7[583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[584]),
        .S(self_sf7[584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[585]),
        .S(self_sf7[585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[586]),
        .S(self_sf7[586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[587]),
        .S(self_sf7[587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[588]),
        .S(self_sf7[588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[589]),
        .S(self_sf7[589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[58].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[58]),
        .S(self_sf7[58]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[590]),
        .S(self_sf7[590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[591]),
        .S(self_sf7[591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[592]),
        .S(self_sf7[592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[593]),
        .S(self_sf7[593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[594]),
        .S(self_sf7[594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[595]),
        .S(self_sf7[595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[596]),
        .S(self_sf7[596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[597]),
        .S(self_sf7[597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[598]),
        .S(self_sf7[598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[599]),
        .S(self_sf7[599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[59].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[59]),
        .S(self_sf7[59]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[5].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[5]),
        .S(info_sf7[5]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[600]),
        .S(self_sf7[600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[601]),
        .S(self_sf7[601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[602]),
        .S(self_sf7[602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[603]),
        .S(self_sf7[603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[604]),
        .S(self_sf7[604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[605]),
        .S(self_sf7[605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[606]),
        .S(self_sf7[606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[607]),
        .S(self_sf7[607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[608]),
        .S(self_sf7[608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[609]),
        .S(self_sf7[609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[60].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[60]),
        .S(self_sf7[60]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[610]),
        .S(self_sf7[610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[611]),
        .S(self_sf7[611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[612]),
        .S(self_sf7[612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[613]),
        .S(self_sf7[613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[614]),
        .S(self_sf7[614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[615]),
        .S(self_sf7[615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[616]),
        .S(self_sf7[616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[617]),
        .S(self_sf7[617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[618]),
        .S(self_sf7[618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[619]),
        .S(self_sf7[619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[61].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[61]),
        .S(self_sf7[61]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[620]),
        .S(self_sf7[620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[621]),
        .S(self_sf7[621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[622]),
        .S(self_sf7[622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[623]),
        .S(self_sf7[623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[624]),
        .S(self_sf7[624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[625]),
        .S(self_sf7[625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[626]),
        .S(self_sf7[626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[627]),
        .S(self_sf7[627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[628]),
        .S(self_sf7[628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[629]),
        .S(self_sf7[629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[62].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[62]),
        .S(self_sf7[62]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[630]),
        .S(self_sf7[630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[631]),
        .S(self_sf7[631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[632]),
        .S(self_sf7[632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[633]),
        .S(self_sf7[633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[634]),
        .S(self_sf7[634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[635]),
        .S(self_sf7[635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[636]),
        .S(self_sf7[636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[637]),
        .S(self_sf7[637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[638]),
        .S(self_sf7[638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[639]),
        .S(self_sf7[639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[63].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[63]),
        .S(self_sf7[63]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[640]),
        .S(self_sf7[640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[641]),
        .S(self_sf7[641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[642]),
        .S(self_sf7[642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[643]),
        .S(self_sf7[643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[644]),
        .S(self_sf7[644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[645]),
        .S(self_sf7[645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[646]),
        .S(self_sf7[646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[647]),
        .S(self_sf7[647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[648]),
        .S(self_sf7[648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[649]),
        .S(self_sf7[649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[64].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[64]),
        .S(self_sf7[64]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[650]),
        .S(self_sf7[650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[651]),
        .S(self_sf7[651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[652]),
        .S(self_sf7[652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[653]),
        .S(self_sf7[653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[654]),
        .S(self_sf7[654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[655]),
        .S(self_sf7[655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[656]),
        .S(self_sf7[656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[657]),
        .S(self_sf7[657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[658]),
        .S(self_sf7[658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[659]),
        .S(self_sf7[659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[65].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[65]),
        .S(self_sf7[65]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[660]),
        .S(self_sf7[660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[661]),
        .S(self_sf7[661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[662]),
        .S(self_sf7[662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[663]),
        .S(self_sf7[663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[664]),
        .S(self_sf7[664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[665]),
        .S(self_sf7[665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[666]),
        .S(self_sf7[666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[667]),
        .S(self_sf7[667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[668]),
        .S(self_sf7[668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[669]),
        .S(self_sf7[669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[66].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[66]),
        .S(self_sf7[66]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[670]),
        .S(self_sf7[670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[671]),
        .S(self_sf7[671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[672]),
        .S(self_sf7[672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[673]),
        .S(self_sf7[673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[674]),
        .S(self_sf7[674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[675]),
        .S(self_sf7[675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[676]),
        .S(self_sf7[676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[677]),
        .S(self_sf7[677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[678]),
        .S(self_sf7[678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[679]),
        .S(self_sf7[679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[67].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[67]),
        .S(self_sf7[67]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[680]),
        .S(self_sf7[680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[681]),
        .S(self_sf7[681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[682]),
        .S(self_sf7[682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[683]),
        .S(self_sf7[683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[684]),
        .S(self_sf7[684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[685]),
        .S(self_sf7[685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[686]),
        .S(self_sf7[686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[687]),
        .S(self_sf7[687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[688]),
        .S(self_sf7[688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[689]),
        .S(self_sf7[689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[68].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[68]),
        .S(self_sf7[68]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[690]),
        .S(self_sf7[690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[691]),
        .S(self_sf7[691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[692]),
        .S(self_sf7[692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[693]),
        .S(self_sf7[693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[694]),
        .S(self_sf7[694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[695]),
        .S(self_sf7[695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[696]),
        .S(self_sf7[696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[697]),
        .S(self_sf7[697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[698]),
        .S(self_sf7[698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[699]),
        .S(self_sf7[699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[69].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[69]),
        .S(self_sf7[69]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[6].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[6]),
        .S(info_sf7[6]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[700]),
        .S(self_sf7[700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[701]),
        .S(self_sf7[701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[702]),
        .S(self_sf7[702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[703]),
        .S(self_sf7[703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[704]),
        .S(self_sf7[704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[705]),
        .S(self_sf7[705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[706]),
        .S(self_sf7[706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[707]),
        .S(self_sf7[707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[708]),
        .S(self_sf7[708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[709]),
        .S(self_sf7[709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[70].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[70]),
        .S(self_sf7[70]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[710]),
        .S(self_sf7[710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[711]),
        .S(self_sf7[711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[712]),
        .S(self_sf7[712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[713]),
        .S(self_sf7[713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[714]),
        .S(self_sf7[714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[715]),
        .S(self_sf7[715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[716]),
        .S(self_sf7[716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[717]),
        .S(self_sf7[717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[718]),
        .S(self_sf7[718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[719]),
        .S(self_sf7[719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[71].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[71]),
        .S(self_sf7[71]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[720]),
        .S(self_sf7[720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[721]),
        .S(self_sf7[721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[722]),
        .S(self_sf7[722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[723]),
        .S(self_sf7[723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[724]),
        .S(self_sf7[724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[725]),
        .S(self_sf7[725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[726]),
        .S(self_sf7[726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[727]),
        .S(self_sf7[727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[728]),
        .S(self_sf7[728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[729]),
        .S(self_sf7[729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[72].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[72]),
        .S(self_sf7[72]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[730]),
        .S(self_sf7[730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[731]),
        .S(self_sf7[731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[732]),
        .S(self_sf7[732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[733]),
        .S(self_sf7[733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[734]),
        .S(self_sf7[734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[735]),
        .S(self_sf7[735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[736]),
        .S(self_sf7[736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[737]),
        .S(self_sf7[737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[738]),
        .S(self_sf7[738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[739]),
        .S(self_sf7[739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[73].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[73]),
        .S(self_sf7[73]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[740]),
        .S(self_sf7[740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[741]),
        .S(self_sf7[741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[742]),
        .S(self_sf7[742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[743]),
        .S(self_sf7[743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[744]),
        .S(self_sf7[744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[745]),
        .S(self_sf7[745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[746]),
        .S(self_sf7[746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[747]),
        .S(self_sf7[747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[748]),
        .S(self_sf7[748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[749]),
        .S(self_sf7[749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[74].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[74]),
        .S(self_sf7[74]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[750]),
        .S(self_sf7[750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[751]),
        .S(self_sf7[751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[752]),
        .S(self_sf7[752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[753]),
        .S(self_sf7[753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[754]),
        .S(self_sf7[754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[755]),
        .S(self_sf7[755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[756]),
        .S(self_sf7[756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[757]),
        .S(self_sf7[757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[758]),
        .S(self_sf7[758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[759]),
        .S(self_sf7[759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[75].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[75]),
        .S(self_sf7[75]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[760]),
        .S(self_sf7[760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[761]),
        .S(self_sf7[761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[762]),
        .S(self_sf7[762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[763]),
        .S(self_sf7[763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[764]),
        .S(self_sf7[764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[765]),
        .S(self_sf7[765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[766]),
        .S(self_sf7[766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[767]),
        .S(self_sf7[767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[768]),
        .S(self_sf7[768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[769]),
        .S(self_sf7[769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[76].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[76]),
        .S(self_sf7[76]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[770]),
        .S(self_sf7[770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[771]),
        .S(self_sf7[771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[772]),
        .S(self_sf7[772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[773]),
        .S(self_sf7[773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[774]),
        .S(self_sf7[774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[775]),
        .S(self_sf7[775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[776]),
        .S(self_sf7[776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[777]),
        .S(self_sf7[777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[778]),
        .S(self_sf7[778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[779]),
        .S(self_sf7[779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[77].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[77]),
        .S(self_sf7[77]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[780]),
        .S(self_sf7[780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[781]),
        .S(self_sf7[781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[782]),
        .S(self_sf7[782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[783]),
        .S(self_sf7[783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[784]),
        .S(self_sf7[784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[785]),
        .S(self_sf7[785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[786]),
        .S(self_sf7[786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[787]),
        .S(self_sf7[787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[788]),
        .S(self_sf7[788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[789]),
        .S(self_sf7[789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[78].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[78]),
        .S(self_sf7[78]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[790]),
        .S(self_sf7[790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[791]),
        .S(self_sf7[791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[792]),
        .S(self_sf7[792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[793]),
        .S(self_sf7[793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[794]),
        .S(self_sf7[794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[795]),
        .S(self_sf7[795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[796]),
        .S(self_sf7[796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[797]),
        .S(self_sf7[797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[798]),
        .S(self_sf7[798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[799]),
        .S(self_sf7[799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[79].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[79]),
        .S(self_sf7[79]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[7].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[7]),
        .S(info_sf7[7]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[800].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[800]),
        .S(self_sf7[800]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[801].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[801]),
        .S(self_sf7[801]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[802].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[802]),
        .S(self_sf7[802]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[803].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[803]),
        .S(self_sf7[803]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[804].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[804]),
        .S(self_sf7[804]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[805].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[805]),
        .S(self_sf7[805]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[806].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[806]),
        .S(self_sf7[806]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[807].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[807]),
        .S(self_sf7[807]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[808].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[808]),
        .S(self_sf7[808]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[809].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[809]),
        .S(self_sf7[809]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[80].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[80]),
        .S(self_sf7[80]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[810].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[810]),
        .S(self_sf7[810]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[811].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[811]),
        .S(self_sf7[811]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[812].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[812]),
        .S(self_sf7[812]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[813].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[813]),
        .S(self_sf7[813]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[814].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[814]),
        .S(self_sf7[814]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[815].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[815]),
        .S(self_sf7[815]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[816].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[816]),
        .S(self_sf7[816]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[817].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[817]),
        .S(self_sf7[817]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[818].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[818]),
        .S(self_sf7[818]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[819].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[819]),
        .S(self_sf7[819]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[81].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[81]),
        .S(self_sf7[81]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[820].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[820]),
        .S(self_sf7[820]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[821].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[821]),
        .S(self_sf7[821]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[822].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[822]),
        .S(self_sf7[822]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[823].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[823]),
        .S(self_sf7[823]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[824].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[824]),
        .S(self_sf7[824]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[825].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[825]),
        .S(self_sf7[825]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[826].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[826]),
        .S(self_sf7[826]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[827].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[827]),
        .S(self_sf7[827]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[828].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[828]),
        .S(self_sf7[828]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[829].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[829]),
        .S(self_sf7[829]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[82].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[82]),
        .S(self_sf7[82]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[830].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[830]),
        .S(self_sf7[830]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[831].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[831]),
        .S(self_sf7[831]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[832].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[832]),
        .S(self_sf7[832]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[833].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[833]),
        .S(self_sf7[833]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[834].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[834]),
        .S(self_sf7[834]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[835].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[835]),
        .S(self_sf7[835]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[836].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[836]),
        .S(self_sf7[836]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[837].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[837]),
        .S(self_sf7[837]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[838].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[838]),
        .S(self_sf7[838]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[839].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[839]),
        .S(self_sf7[839]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[83].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[83]),
        .S(self_sf7[83]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[840].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[840]),
        .S(self_sf7[840]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[841].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[841]),
        .S(self_sf7[841]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[842].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[842]),
        .S(self_sf7[842]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[843].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[843]),
        .S(self_sf7[843]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[844].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[844]),
        .S(self_sf7[844]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[845].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[845]),
        .S(self_sf7[845]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[846].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[846]),
        .S(self_sf7[846]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[847].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[847]),
        .S(self_sf7[847]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[848].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[848]),
        .S(self_sf7[848]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[849].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[849]),
        .S(self_sf7[849]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[84].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[84]),
        .S(self_sf7[84]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[850].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[850]),
        .S(self_sf7[850]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[851].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[851]),
        .S(self_sf7[851]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[852].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[852]),
        .S(self_sf7[852]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[853].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[853]),
        .S(self_sf7[853]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[854].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[854]),
        .S(self_sf7[854]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[855].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[855]),
        .S(self_sf7[855]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[856].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[856]),
        .S(self_sf7[856]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[857].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[857]),
        .S(self_sf7[857]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[858].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[858]),
        .S(self_sf7[858]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[859].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[859]),
        .S(self_sf7[859]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[85].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[85]),
        .S(self_sf7[85]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[860].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[860]),
        .S(self_sf7[860]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[861].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[861]),
        .S(self_sf7[861]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[862].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[862]),
        .S(self_sf7[862]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[863].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[863]),
        .S(self_sf7[863]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[864].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[864]),
        .S(self_sf7[864]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[865].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[865]),
        .S(self_sf7[865]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[866].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[866]),
        .S(self_sf7[866]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[867].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[867]),
        .S(self_sf7[867]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[868].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[868]),
        .S(self_sf7[868]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[869].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[869]),
        .S(self_sf7[869]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[86].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[86]),
        .S(self_sf7[86]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[870].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[870]),
        .S(self_sf7[870]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[871].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[871]),
        .S(self_sf7[871]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[872].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[872]),
        .S(self_sf7[872]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[873].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[873]),
        .S(self_sf7[873]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[874].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[874]),
        .S(self_sf7[874]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[875].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[875]),
        .S(self_sf7[875]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[876].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[876]),
        .S(self_sf7[876]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[877].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[877]),
        .S(self_sf7[877]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[878].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[878]),
        .S(self_sf7[878]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[879].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[879]),
        .S(self_sf7[879]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[87].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[87]),
        .S(self_sf7[87]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[880].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[880]),
        .S(self_sf7[880]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[881].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[881]),
        .S(self_sf7[881]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[882].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[882]),
        .S(self_sf7[882]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[883].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[883]),
        .S(self_sf7[883]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[884].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[884]),
        .S(self_sf7[884]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[885].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[885]),
        .S(self_sf7[885]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[886].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[886]),
        .S(self_sf7[886]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[887].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[887]),
        .S(self_sf7[887]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[888].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[888]),
        .S(self_sf7[888]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[889].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[889]),
        .S(self_sf7[889]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[88].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[88]),
        .S(self_sf7[88]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[890].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[890]),
        .S(self_sf7[890]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[891].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[891]),
        .S(self_sf7[891]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[892].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[892]),
        .S(self_sf7[892]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[893].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[893]),
        .S(self_sf7[893]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[894].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[894]),
        .S(self_sf7[894]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[895].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[895]),
        .S(self_sf7[895]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[896].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[896]),
        .S(self_sf7[896]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[897].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[897]),
        .S(self_sf7[897]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[898].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[898]),
        .S(self_sf7[898]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[899].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[899]),
        .S(self_sf7[899]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[89].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[89]),
        .S(self_sf7[89]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[8].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[8]),
        .S(self_sf7[8]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[900].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[900]),
        .S(self_sf7[900]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[901].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[901]),
        .S(self_sf7[901]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[902].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[902]),
        .S(self_sf7[902]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[903].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[903]),
        .S(self_sf7[903]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[904].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[904]),
        .S(self_sf7[904]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[905].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[905]),
        .S(self_sf7[905]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[906].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[906]),
        .S(self_sf7[906]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[907].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[907]),
        .S(self_sf7[907]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[908].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[908]),
        .S(self_sf7[908]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[909].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[909]),
        .S(self_sf7[909]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[90].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[90]),
        .S(self_sf7[90]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[910].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[910]),
        .S(self_sf7[910]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[911].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[911]),
        .S(self_sf7[911]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[912].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[912]),
        .S(self_sf7[912]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[913].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[913]),
        .S(self_sf7[913]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[914].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[914]),
        .S(self_sf7[914]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[915].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[915]),
        .S(self_sf7[915]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[916].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[916]),
        .S(self_sf7[916]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[917].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[917]),
        .S(self_sf7[917]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[918].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[918]),
        .S(self_sf7[918]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[919].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[919]),
        .S(self_sf7[919]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[91].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[91]),
        .S(self_sf7[91]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[920].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[920]),
        .S(self_sf7[920]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[921].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[921]),
        .S(self_sf7[921]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[922].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[922]),
        .S(self_sf7[922]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[923].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[923]),
        .S(self_sf7[923]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[924].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[924]),
        .S(self_sf7[924]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[925].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[925]),
        .S(self_sf7[925]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[926].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[926]),
        .S(self_sf7[926]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[927].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[927]),
        .S(self_sf7[927]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[928].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[928]),
        .S(self_sf7[928]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[929].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[929]),
        .S(self_sf7[929]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[92].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[92]),
        .S(self_sf7[92]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[930].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[930]),
        .S(self_sf7[930]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[931].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[931]),
        .S(self_sf7[931]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[932].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[932]),
        .S(self_sf7[932]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[933].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[933]),
        .S(self_sf7[933]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[934].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[934]),
        .S(self_sf7[934]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[935].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[935]),
        .S(self_sf7[935]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[936].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[936]),
        .S(self_sf7[936]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[937].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[937]),
        .S(self_sf7[937]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[938].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[938]),
        .S(self_sf7[938]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[939].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[939]),
        .S(self_sf7[939]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[93].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[93]),
        .S(self_sf7[93]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[940].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[940]),
        .S(self_sf7[940]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[941].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[941]),
        .S(self_sf7[941]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[942].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[942]),
        .S(self_sf7[942]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[943].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[943]),
        .S(self_sf7[943]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[944].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[944]),
        .S(self_sf7[944]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[945].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[945]),
        .S(self_sf7[945]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[946].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[946]),
        .S(self_sf7[946]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[947].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[947]),
        .S(self_sf7[947]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[948].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[948]),
        .S(self_sf7[948]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[949].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[949]),
        .S(self_sf7[949]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[94].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[94]),
        .S(self_sf7[94]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[950].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[950]),
        .S(self_sf7[950]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[951].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[951]),
        .S(self_sf7[951]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[952].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[952]),
        .S(self_sf7[952]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[953].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[953]),
        .S(self_sf7[953]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[954].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[954]),
        .S(self_sf7[954]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[955].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[955]),
        .S(self_sf7[955]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[956].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[956]),
        .S(self_sf7[956]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[957].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[957]),
        .S(self_sf7[957]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[958].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[958]),
        .S(self_sf7[958]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[959].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[959]),
        .S(self_sf7[959]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[95].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[95]),
        .S(self_sf7[95]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[960].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[960]),
        .S(self_sf7[960]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[961].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[961]),
        .S(self_sf7[961]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[962].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[962]),
        .S(self_sf7[962]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[963].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[963]),
        .S(self_sf7[963]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[964].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[964]),
        .S(self_sf7[964]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[965].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[965]),
        .S(self_sf7[965]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[966].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[966]),
        .S(self_sf7[966]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[967].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[967]),
        .S(self_sf7[967]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[968].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[968]),
        .S(self_sf7[968]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[969].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[969]),
        .S(self_sf7[969]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[96].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[96]),
        .S(self_sf7[96]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[970].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[970]),
        .S(self_sf7[970]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[971].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[971]),
        .S(self_sf7[971]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[972].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[972]),
        .S(self_sf7[972]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[973].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[973]),
        .S(self_sf7[973]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[974].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[974]),
        .S(self_sf7[974]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[975].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[975]),
        .S(self_sf7[975]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[976].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[976]),
        .S(self_sf7[976]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[977].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[977]),
        .S(self_sf7[977]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[978].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[978]),
        .S(self_sf7[978]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[979].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[979]),
        .S(self_sf7[979]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[97].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[97]),
        .S(self_sf7[97]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[980].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[980]),
        .S(self_sf7[980]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[981].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[981]),
        .S(self_sf7[981]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[982].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[982]),
        .S(self_sf7[982]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[983].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[983]),
        .S(self_sf7[983]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[984].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[984]),
        .S(self_sf7[984]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[985].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[985]),
        .S(self_sf7[985]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[986].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[986]),
        .S(self_sf7[986]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[987].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[987]),
        .S(self_sf7[987]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[988].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[988]),
        .S(self_sf7[988]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[989].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[989]),
        .S(self_sf7[989]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[98].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[98]),
        .S(self_sf7[98]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[990].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[990]),
        .S(self_sf7[990]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[991].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[991]),
        .S(self_sf7[991]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[992].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[992]),
        .S(self_sf7[992]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[993].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[993]),
        .S(self_sf7[993]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[994].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[994]),
        .S(self_sf7[994]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[995].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[995]),
        .S(self_sf7[995]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[996].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[996]),
        .S(self_sf7[996]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[997].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[997]),
        .S(self_sf7[997]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[998].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[998]),
        .S(self_sf7[998]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[999].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[999]),
        .S(self_sf7[999]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[99].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[99]),
        .S(self_sf7[99]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[9].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[9]),
        .S(self_sf7[9]));
  (* BOX_TYPE = "black_box" *) 
  MUXF8 \activity_ROsf8[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf8[0]),
        .S(self_sf8[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF9 \activity_ROsf9[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf9[0]),
        .S(self_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_0
       (.I0(1'b0),
        .O(self_sf7[1802]));
  LUT1 #(
    .INIT(2'h2)) 
    i_1
       (.I0(1'b0),
        .O(self_sf7[1801]));
  LUT1 #(
    .INIT(2'h2)) 
    i_10
       (.I0(1'b0),
        .O(info_sf8[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_11
       (.I0(1'b0),
        .O(info_sf8[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_12
       (.I0(1'b0),
        .O(info_sf8[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_13
       (.I0(1'b0),
        .O(info_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_14
       (.I0(1'b0),
        .O(info_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_15
       (.I0(1'b0),
        .O(info_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_16
       (.I0(1'b0),
        .O(info_sf8[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_17
       (.I0(1'b0),
        .O(info_sf9[7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_18
       (.I0(1'b0),
        .O(info_sf9[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_19
       (.I0(1'b0),
        .O(info_sf9[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_2
       (.I0(1'b0),
        .O(self_sf7[1800]));
  LUT1 #(
    .INIT(2'h2)) 
    i_20
       (.I0(1'b0),
        .O(info_sf9[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_21
       (.I0(1'b0),
        .O(info_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_22
       (.I0(1'b0),
        .O(info_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_23
       (.I0(1'b0),
        .O(info_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_24
       (.I0(1'b0),
        .O(info_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_3
       (.I0(1'b0),
        .O(self_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_4
       (.I0(1'b0),
        .O(self_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_5
       (.I0(1'b0),
        .O(self_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_6
       (.I0(1'b0),
        .O(self_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_7
       (.I0(1'b0),
        .O(self_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_8
       (.I0(1'b0),
        .O(self_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_9
       (.I0(1'b0),
        .O(info_sf8[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst
       (.I0(self_sf7[7]),
        .O(info_sf7[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__0
       (.I0(self_sf7[6]),
        .O(info_sf7[6]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__1
       (.I0(self_sf7[5]),
        .O(info_sf7[5]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__2
       (.I0(self_sf7[4]),
        .O(info_sf7[4]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__3
       (.I0(self_sf7[3]),
        .O(info_sf7[3]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__4
       (.I0(self_sf7[2]),
        .O(info_sf7[2]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__5
       (.I0(self_sf7[1]),
        .O(info_sf7[1]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__6
       (.I0(self_sf7[0]),
        .O(info_sf7[0]));
endmodule

(* ORIG_REF_NAME = "muxer" *) (* box_type = "black_box" *) (* dont_touch = "true" *) 
module switch_elements_muxer__6
   (enable_i,
    info_o);
  input enable_i;
  output info_o;

  wire enable_i;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf7;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf8;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf9;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [1802:0]self_sf7;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf8;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf9;

  assign info_o = info_sf7[1];
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[0]),
        .S(info_sf7[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1000].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1000]),
        .S(self_sf7[1000]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1001].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1001]),
        .S(self_sf7[1001]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1002].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1002]),
        .S(self_sf7[1002]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1003].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1003]),
        .S(self_sf7[1003]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1004].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1004]),
        .S(self_sf7[1004]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1005].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1005]),
        .S(self_sf7[1005]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1006].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1006]),
        .S(self_sf7[1006]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1007].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1007]),
        .S(self_sf7[1007]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1008].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1008]),
        .S(self_sf7[1008]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1009].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1009]),
        .S(self_sf7[1009]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[100]),
        .S(self_sf7[100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1010].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1010]),
        .S(self_sf7[1010]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1011].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1011]),
        .S(self_sf7[1011]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1012].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1012]),
        .S(self_sf7[1012]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1013].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1013]),
        .S(self_sf7[1013]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1014].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1014]),
        .S(self_sf7[1014]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1015].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1015]),
        .S(self_sf7[1015]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1016].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1016]),
        .S(self_sf7[1016]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1017].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1017]),
        .S(self_sf7[1017]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1018].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1018]),
        .S(self_sf7[1018]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1019].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1019]),
        .S(self_sf7[1019]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[101]),
        .S(self_sf7[101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1020].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1020]),
        .S(self_sf7[1020]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1021].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1021]),
        .S(self_sf7[1021]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1022].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1022]),
        .S(self_sf7[1022]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1023].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1023]),
        .S(self_sf7[1023]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1024].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1024]),
        .S(self_sf7[1024]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1025].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1025]),
        .S(self_sf7[1025]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1026].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1026]),
        .S(self_sf7[1026]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1027].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1027]),
        .S(self_sf7[1027]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1028].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1028]),
        .S(self_sf7[1028]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1029].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1029]),
        .S(self_sf7[1029]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[102]),
        .S(self_sf7[102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1030].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1030]),
        .S(self_sf7[1030]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1031].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1031]),
        .S(self_sf7[1031]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1032].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1032]),
        .S(self_sf7[1032]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1033].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1033]),
        .S(self_sf7[1033]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1034].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1034]),
        .S(self_sf7[1034]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1035].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1035]),
        .S(self_sf7[1035]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1036].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1036]),
        .S(self_sf7[1036]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1037].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1037]),
        .S(self_sf7[1037]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1038].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1038]),
        .S(self_sf7[1038]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1039].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1039]),
        .S(self_sf7[1039]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[103]),
        .S(self_sf7[103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1040].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1040]),
        .S(self_sf7[1040]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1041].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1041]),
        .S(self_sf7[1041]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1042].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1042]),
        .S(self_sf7[1042]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1043].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1043]),
        .S(self_sf7[1043]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1044].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1044]),
        .S(self_sf7[1044]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1045].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1045]),
        .S(self_sf7[1045]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1046].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1046]),
        .S(self_sf7[1046]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1047].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1047]),
        .S(self_sf7[1047]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1048].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1048]),
        .S(self_sf7[1048]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1049].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1049]),
        .S(self_sf7[1049]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[104]),
        .S(self_sf7[104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1050].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1050]),
        .S(self_sf7[1050]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1051].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1051]),
        .S(self_sf7[1051]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1052].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1052]),
        .S(self_sf7[1052]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1053].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1053]),
        .S(self_sf7[1053]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1054].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1054]),
        .S(self_sf7[1054]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1055].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1055]),
        .S(self_sf7[1055]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1056].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1056]),
        .S(self_sf7[1056]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1057].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1057]),
        .S(self_sf7[1057]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1058].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1058]),
        .S(self_sf7[1058]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1059].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1059]),
        .S(self_sf7[1059]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[105]),
        .S(self_sf7[105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1060].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1060]),
        .S(self_sf7[1060]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1061].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1061]),
        .S(self_sf7[1061]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1062].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1062]),
        .S(self_sf7[1062]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1063].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1063]),
        .S(self_sf7[1063]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1064].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1064]),
        .S(self_sf7[1064]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1065].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1065]),
        .S(self_sf7[1065]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1066].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1066]),
        .S(self_sf7[1066]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1067].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1067]),
        .S(self_sf7[1067]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1068].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1068]),
        .S(self_sf7[1068]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1069].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1069]),
        .S(self_sf7[1069]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[106]),
        .S(self_sf7[106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1070].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1070]),
        .S(self_sf7[1070]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1071].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1071]),
        .S(self_sf7[1071]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1072].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1072]),
        .S(self_sf7[1072]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1073].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1073]),
        .S(self_sf7[1073]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1074].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1074]),
        .S(self_sf7[1074]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1075].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1075]),
        .S(self_sf7[1075]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1076].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1076]),
        .S(self_sf7[1076]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1077].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1077]),
        .S(self_sf7[1077]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1078].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1078]),
        .S(self_sf7[1078]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1079].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1079]),
        .S(self_sf7[1079]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[107]),
        .S(self_sf7[107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1080].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1080]),
        .S(self_sf7[1080]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1081].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1081]),
        .S(self_sf7[1081]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1082].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1082]),
        .S(self_sf7[1082]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1083].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1083]),
        .S(self_sf7[1083]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1084].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1084]),
        .S(self_sf7[1084]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1085].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1085]),
        .S(self_sf7[1085]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1086].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1086]),
        .S(self_sf7[1086]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1087].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1087]),
        .S(self_sf7[1087]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1088].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1088]),
        .S(self_sf7[1088]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1089].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1089]),
        .S(self_sf7[1089]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[108]),
        .S(self_sf7[108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1090].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1090]),
        .S(self_sf7[1090]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1091].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1091]),
        .S(self_sf7[1091]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1092].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1092]),
        .S(self_sf7[1092]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1093].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1093]),
        .S(self_sf7[1093]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1094].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1094]),
        .S(self_sf7[1094]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1095].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1095]),
        .S(self_sf7[1095]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1096].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1096]),
        .S(self_sf7[1096]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1097].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1097]),
        .S(self_sf7[1097]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1098].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1098]),
        .S(self_sf7[1098]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1099].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1099]),
        .S(self_sf7[1099]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[109]),
        .S(self_sf7[109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[10].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[10]),
        .S(self_sf7[10]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1100]),
        .S(self_sf7[1100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1101]),
        .S(self_sf7[1101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1102]),
        .S(self_sf7[1102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1103]),
        .S(self_sf7[1103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1104]),
        .S(self_sf7[1104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1105]),
        .S(self_sf7[1105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1106]),
        .S(self_sf7[1106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1107]),
        .S(self_sf7[1107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1108]),
        .S(self_sf7[1108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1109]),
        .S(self_sf7[1109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[110]),
        .S(self_sf7[110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1110]),
        .S(self_sf7[1110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1111]),
        .S(self_sf7[1111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1112]),
        .S(self_sf7[1112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1113]),
        .S(self_sf7[1113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1114]),
        .S(self_sf7[1114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1115]),
        .S(self_sf7[1115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1116]),
        .S(self_sf7[1116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1117]),
        .S(self_sf7[1117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1118]),
        .S(self_sf7[1118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1119]),
        .S(self_sf7[1119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[111]),
        .S(self_sf7[111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1120]),
        .S(self_sf7[1120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1121]),
        .S(self_sf7[1121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1122]),
        .S(self_sf7[1122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1123]),
        .S(self_sf7[1123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1124]),
        .S(self_sf7[1124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1125]),
        .S(self_sf7[1125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1126]),
        .S(self_sf7[1126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1127]),
        .S(self_sf7[1127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1128]),
        .S(self_sf7[1128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1129]),
        .S(self_sf7[1129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[112]),
        .S(self_sf7[112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1130]),
        .S(self_sf7[1130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1131]),
        .S(self_sf7[1131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1132]),
        .S(self_sf7[1132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1133]),
        .S(self_sf7[1133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1134]),
        .S(self_sf7[1134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1135]),
        .S(self_sf7[1135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1136]),
        .S(self_sf7[1136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1137]),
        .S(self_sf7[1137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1138]),
        .S(self_sf7[1138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1139]),
        .S(self_sf7[1139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[113]),
        .S(self_sf7[113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1140]),
        .S(self_sf7[1140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1141]),
        .S(self_sf7[1141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1142]),
        .S(self_sf7[1142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1143]),
        .S(self_sf7[1143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1144]),
        .S(self_sf7[1144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1145]),
        .S(self_sf7[1145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1146]),
        .S(self_sf7[1146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1147]),
        .S(self_sf7[1147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1148]),
        .S(self_sf7[1148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1149]),
        .S(self_sf7[1149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[114]),
        .S(self_sf7[114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1150]),
        .S(self_sf7[1150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1151]),
        .S(self_sf7[1151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1152]),
        .S(self_sf7[1152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1153]),
        .S(self_sf7[1153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1154]),
        .S(self_sf7[1154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1155]),
        .S(self_sf7[1155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1156]),
        .S(self_sf7[1156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1157]),
        .S(self_sf7[1157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1158]),
        .S(self_sf7[1158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1159]),
        .S(self_sf7[1159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[115]),
        .S(self_sf7[115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1160]),
        .S(self_sf7[1160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1161]),
        .S(self_sf7[1161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1162]),
        .S(self_sf7[1162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1163]),
        .S(self_sf7[1163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1164]),
        .S(self_sf7[1164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1165]),
        .S(self_sf7[1165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1166]),
        .S(self_sf7[1166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1167]),
        .S(self_sf7[1167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1168]),
        .S(self_sf7[1168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1169]),
        .S(self_sf7[1169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[116]),
        .S(self_sf7[116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1170]),
        .S(self_sf7[1170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1171]),
        .S(self_sf7[1171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1172]),
        .S(self_sf7[1172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1173]),
        .S(self_sf7[1173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1174]),
        .S(self_sf7[1174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1175]),
        .S(self_sf7[1175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1176]),
        .S(self_sf7[1176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1177]),
        .S(self_sf7[1177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1178]),
        .S(self_sf7[1178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1179]),
        .S(self_sf7[1179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[117]),
        .S(self_sf7[117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1180]),
        .S(self_sf7[1180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1181]),
        .S(self_sf7[1181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1182]),
        .S(self_sf7[1182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1183]),
        .S(self_sf7[1183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1184]),
        .S(self_sf7[1184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1185]),
        .S(self_sf7[1185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1186]),
        .S(self_sf7[1186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1187]),
        .S(self_sf7[1187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1188]),
        .S(self_sf7[1188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1189]),
        .S(self_sf7[1189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[118]),
        .S(self_sf7[118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1190]),
        .S(self_sf7[1190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1191]),
        .S(self_sf7[1191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1192]),
        .S(self_sf7[1192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1193]),
        .S(self_sf7[1193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1194]),
        .S(self_sf7[1194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1195]),
        .S(self_sf7[1195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1196]),
        .S(self_sf7[1196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1197]),
        .S(self_sf7[1197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1198]),
        .S(self_sf7[1198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1199]),
        .S(self_sf7[1199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[119]),
        .S(self_sf7[119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[11].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[11]),
        .S(self_sf7[11]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1200]),
        .S(self_sf7[1200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1201]),
        .S(self_sf7[1201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1202]),
        .S(self_sf7[1202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1203]),
        .S(self_sf7[1203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1204]),
        .S(self_sf7[1204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1205]),
        .S(self_sf7[1205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1206]),
        .S(self_sf7[1206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1207]),
        .S(self_sf7[1207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1208]),
        .S(self_sf7[1208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1209]),
        .S(self_sf7[1209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[120]),
        .S(self_sf7[120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1210]),
        .S(self_sf7[1210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1211]),
        .S(self_sf7[1211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1212]),
        .S(self_sf7[1212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1213]),
        .S(self_sf7[1213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1214]),
        .S(self_sf7[1214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1215]),
        .S(self_sf7[1215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1216]),
        .S(self_sf7[1216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1217]),
        .S(self_sf7[1217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1218]),
        .S(self_sf7[1218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1219]),
        .S(self_sf7[1219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[121]),
        .S(self_sf7[121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1220]),
        .S(self_sf7[1220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1221]),
        .S(self_sf7[1221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1222]),
        .S(self_sf7[1222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1223]),
        .S(self_sf7[1223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1224]),
        .S(self_sf7[1224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1225]),
        .S(self_sf7[1225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1226]),
        .S(self_sf7[1226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1227]),
        .S(self_sf7[1227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1228]),
        .S(self_sf7[1228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1229]),
        .S(self_sf7[1229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[122]),
        .S(self_sf7[122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1230]),
        .S(self_sf7[1230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1231]),
        .S(self_sf7[1231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1232]),
        .S(self_sf7[1232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1233]),
        .S(self_sf7[1233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1234]),
        .S(self_sf7[1234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1235]),
        .S(self_sf7[1235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1236]),
        .S(self_sf7[1236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1237]),
        .S(self_sf7[1237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1238]),
        .S(self_sf7[1238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1239]),
        .S(self_sf7[1239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[123]),
        .S(self_sf7[123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1240]),
        .S(self_sf7[1240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1241]),
        .S(self_sf7[1241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1242]),
        .S(self_sf7[1242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1243]),
        .S(self_sf7[1243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1244]),
        .S(self_sf7[1244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1245]),
        .S(self_sf7[1245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1246]),
        .S(self_sf7[1246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1247]),
        .S(self_sf7[1247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1248]),
        .S(self_sf7[1248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1249]),
        .S(self_sf7[1249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[124]),
        .S(self_sf7[124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1250]),
        .S(self_sf7[1250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1251]),
        .S(self_sf7[1251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1252]),
        .S(self_sf7[1252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1253]),
        .S(self_sf7[1253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1254]),
        .S(self_sf7[1254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1255]),
        .S(self_sf7[1255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1256]),
        .S(self_sf7[1256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1257]),
        .S(self_sf7[1257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1258]),
        .S(self_sf7[1258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1259]),
        .S(self_sf7[1259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[125]),
        .S(self_sf7[125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1260]),
        .S(self_sf7[1260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1261]),
        .S(self_sf7[1261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1262]),
        .S(self_sf7[1262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1263]),
        .S(self_sf7[1263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1264]),
        .S(self_sf7[1264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1265]),
        .S(self_sf7[1265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1266]),
        .S(self_sf7[1266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1267]),
        .S(self_sf7[1267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1268]),
        .S(self_sf7[1268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1269]),
        .S(self_sf7[1269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[126]),
        .S(self_sf7[126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1270]),
        .S(self_sf7[1270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1271]),
        .S(self_sf7[1271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1272]),
        .S(self_sf7[1272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1273]),
        .S(self_sf7[1273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1274]),
        .S(self_sf7[1274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1275]),
        .S(self_sf7[1275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1276]),
        .S(self_sf7[1276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1277]),
        .S(self_sf7[1277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1278]),
        .S(self_sf7[1278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1279]),
        .S(self_sf7[1279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[127]),
        .S(self_sf7[127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1280]),
        .S(self_sf7[1280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1281]),
        .S(self_sf7[1281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1282]),
        .S(self_sf7[1282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1283]),
        .S(self_sf7[1283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1284]),
        .S(self_sf7[1284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1285]),
        .S(self_sf7[1285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1286]),
        .S(self_sf7[1286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1287]),
        .S(self_sf7[1287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1288]),
        .S(self_sf7[1288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1289]),
        .S(self_sf7[1289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[128]),
        .S(self_sf7[128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1290]),
        .S(self_sf7[1290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1291]),
        .S(self_sf7[1291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1292]),
        .S(self_sf7[1292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1293]),
        .S(self_sf7[1293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1294]),
        .S(self_sf7[1294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1295]),
        .S(self_sf7[1295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1296]),
        .S(self_sf7[1296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1297]),
        .S(self_sf7[1297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1298]),
        .S(self_sf7[1298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1299]),
        .S(self_sf7[1299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[129]),
        .S(self_sf7[129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[12].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[12]),
        .S(self_sf7[12]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1300]),
        .S(self_sf7[1300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1301]),
        .S(self_sf7[1301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1302]),
        .S(self_sf7[1302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1303]),
        .S(self_sf7[1303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1304]),
        .S(self_sf7[1304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1305]),
        .S(self_sf7[1305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1306]),
        .S(self_sf7[1306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1307]),
        .S(self_sf7[1307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1308]),
        .S(self_sf7[1308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1309]),
        .S(self_sf7[1309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[130]),
        .S(self_sf7[130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1310]),
        .S(self_sf7[1310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1311]),
        .S(self_sf7[1311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1312]),
        .S(self_sf7[1312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1313]),
        .S(self_sf7[1313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1314]),
        .S(self_sf7[1314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1315]),
        .S(self_sf7[1315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1316]),
        .S(self_sf7[1316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1317]),
        .S(self_sf7[1317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1318]),
        .S(self_sf7[1318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1319]),
        .S(self_sf7[1319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[131]),
        .S(self_sf7[131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1320]),
        .S(self_sf7[1320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1321]),
        .S(self_sf7[1321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1322]),
        .S(self_sf7[1322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1323]),
        .S(self_sf7[1323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1324]),
        .S(self_sf7[1324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1325]),
        .S(self_sf7[1325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1326]),
        .S(self_sf7[1326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1327]),
        .S(self_sf7[1327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1328]),
        .S(self_sf7[1328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1329]),
        .S(self_sf7[1329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[132]),
        .S(self_sf7[132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1330]),
        .S(self_sf7[1330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1331]),
        .S(self_sf7[1331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1332]),
        .S(self_sf7[1332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1333]),
        .S(self_sf7[1333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1334]),
        .S(self_sf7[1334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1335]),
        .S(self_sf7[1335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1336]),
        .S(self_sf7[1336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1337]),
        .S(self_sf7[1337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1338]),
        .S(self_sf7[1338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1339]),
        .S(self_sf7[1339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[133]),
        .S(self_sf7[133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1340]),
        .S(self_sf7[1340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1341]),
        .S(self_sf7[1341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1342]),
        .S(self_sf7[1342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1343]),
        .S(self_sf7[1343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1344]),
        .S(self_sf7[1344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1345]),
        .S(self_sf7[1345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1346]),
        .S(self_sf7[1346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1347]),
        .S(self_sf7[1347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1348]),
        .S(self_sf7[1348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1349]),
        .S(self_sf7[1349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[134]),
        .S(self_sf7[134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1350]),
        .S(self_sf7[1350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1351]),
        .S(self_sf7[1351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1352]),
        .S(self_sf7[1352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1353]),
        .S(self_sf7[1353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1354]),
        .S(self_sf7[1354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1355]),
        .S(self_sf7[1355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1356]),
        .S(self_sf7[1356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1357]),
        .S(self_sf7[1357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1358]),
        .S(self_sf7[1358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1359]),
        .S(self_sf7[1359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[135]),
        .S(self_sf7[135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1360]),
        .S(self_sf7[1360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1361]),
        .S(self_sf7[1361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1362]),
        .S(self_sf7[1362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1363]),
        .S(self_sf7[1363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1364]),
        .S(self_sf7[1364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1365]),
        .S(self_sf7[1365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1366]),
        .S(self_sf7[1366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1367]),
        .S(self_sf7[1367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1368]),
        .S(self_sf7[1368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1369]),
        .S(self_sf7[1369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[136]),
        .S(self_sf7[136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1370]),
        .S(self_sf7[1370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1371]),
        .S(self_sf7[1371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1372]),
        .S(self_sf7[1372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1373]),
        .S(self_sf7[1373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1374]),
        .S(self_sf7[1374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1375]),
        .S(self_sf7[1375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1376]),
        .S(self_sf7[1376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1377]),
        .S(self_sf7[1377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1378]),
        .S(self_sf7[1378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1379]),
        .S(self_sf7[1379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[137]),
        .S(self_sf7[137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1380]),
        .S(self_sf7[1380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1381]),
        .S(self_sf7[1381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1382]),
        .S(self_sf7[1382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1383]),
        .S(self_sf7[1383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1384]),
        .S(self_sf7[1384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1385]),
        .S(self_sf7[1385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1386]),
        .S(self_sf7[1386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1387]),
        .S(self_sf7[1387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1388]),
        .S(self_sf7[1388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1389]),
        .S(self_sf7[1389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[138]),
        .S(self_sf7[138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1390]),
        .S(self_sf7[1390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1391]),
        .S(self_sf7[1391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1392]),
        .S(self_sf7[1392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1393]),
        .S(self_sf7[1393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1394]),
        .S(self_sf7[1394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1395]),
        .S(self_sf7[1395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1396]),
        .S(self_sf7[1396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1397]),
        .S(self_sf7[1397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1398]),
        .S(self_sf7[1398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1399]),
        .S(self_sf7[1399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[139]),
        .S(self_sf7[139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[13].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[13]),
        .S(self_sf7[13]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1400]),
        .S(self_sf7[1400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1401]),
        .S(self_sf7[1401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1402]),
        .S(self_sf7[1402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1403]),
        .S(self_sf7[1403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1404]),
        .S(self_sf7[1404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1405]),
        .S(self_sf7[1405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1406]),
        .S(self_sf7[1406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1407]),
        .S(self_sf7[1407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1408]),
        .S(self_sf7[1408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1409]),
        .S(self_sf7[1409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[140]),
        .S(self_sf7[140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1410]),
        .S(self_sf7[1410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1411]),
        .S(self_sf7[1411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1412]),
        .S(self_sf7[1412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1413]),
        .S(self_sf7[1413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1414]),
        .S(self_sf7[1414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1415]),
        .S(self_sf7[1415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1416]),
        .S(self_sf7[1416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1417]),
        .S(self_sf7[1417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1418]),
        .S(self_sf7[1418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1419]),
        .S(self_sf7[1419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[141]),
        .S(self_sf7[141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1420]),
        .S(self_sf7[1420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1421]),
        .S(self_sf7[1421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1422]),
        .S(self_sf7[1422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1423]),
        .S(self_sf7[1423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1424]),
        .S(self_sf7[1424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1425]),
        .S(self_sf7[1425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1426]),
        .S(self_sf7[1426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1427]),
        .S(self_sf7[1427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1428]),
        .S(self_sf7[1428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1429]),
        .S(self_sf7[1429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[142]),
        .S(self_sf7[142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1430]),
        .S(self_sf7[1430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1431]),
        .S(self_sf7[1431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1432]),
        .S(self_sf7[1432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1433]),
        .S(self_sf7[1433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1434]),
        .S(self_sf7[1434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1435]),
        .S(self_sf7[1435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1436]),
        .S(self_sf7[1436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1437]),
        .S(self_sf7[1437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1438]),
        .S(self_sf7[1438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1439]),
        .S(self_sf7[1439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[143]),
        .S(self_sf7[143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1440]),
        .S(self_sf7[1440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1441]),
        .S(self_sf7[1441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1442]),
        .S(self_sf7[1442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1443]),
        .S(self_sf7[1443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1444]),
        .S(self_sf7[1444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1445]),
        .S(self_sf7[1445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1446]),
        .S(self_sf7[1446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1447]),
        .S(self_sf7[1447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1448]),
        .S(self_sf7[1448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1449]),
        .S(self_sf7[1449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[144]),
        .S(self_sf7[144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1450]),
        .S(self_sf7[1450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1451]),
        .S(self_sf7[1451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1452]),
        .S(self_sf7[1452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1453]),
        .S(self_sf7[1453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1454]),
        .S(self_sf7[1454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1455]),
        .S(self_sf7[1455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1456]),
        .S(self_sf7[1456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1457]),
        .S(self_sf7[1457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1458]),
        .S(self_sf7[1458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1459]),
        .S(self_sf7[1459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[145]),
        .S(self_sf7[145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1460]),
        .S(self_sf7[1460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1461]),
        .S(self_sf7[1461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1462]),
        .S(self_sf7[1462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1463]),
        .S(self_sf7[1463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1464]),
        .S(self_sf7[1464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1465]),
        .S(self_sf7[1465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1466]),
        .S(self_sf7[1466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1467]),
        .S(self_sf7[1467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1468]),
        .S(self_sf7[1468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1469]),
        .S(self_sf7[1469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[146]),
        .S(self_sf7[146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1470]),
        .S(self_sf7[1470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1471]),
        .S(self_sf7[1471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1472]),
        .S(self_sf7[1472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1473]),
        .S(self_sf7[1473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1474]),
        .S(self_sf7[1474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1475]),
        .S(self_sf7[1475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1476]),
        .S(self_sf7[1476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1477]),
        .S(self_sf7[1477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1478]),
        .S(self_sf7[1478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1479]),
        .S(self_sf7[1479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[147]),
        .S(self_sf7[147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1480]),
        .S(self_sf7[1480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1481]),
        .S(self_sf7[1481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1482]),
        .S(self_sf7[1482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1483]),
        .S(self_sf7[1483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1484]),
        .S(self_sf7[1484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1485]),
        .S(self_sf7[1485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1486]),
        .S(self_sf7[1486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1487]),
        .S(self_sf7[1487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1488]),
        .S(self_sf7[1488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1489]),
        .S(self_sf7[1489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[148]),
        .S(self_sf7[148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1490]),
        .S(self_sf7[1490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1491]),
        .S(self_sf7[1491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1492]),
        .S(self_sf7[1492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1493]),
        .S(self_sf7[1493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1494]),
        .S(self_sf7[1494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1495]),
        .S(self_sf7[1495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1496]),
        .S(self_sf7[1496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1497]),
        .S(self_sf7[1497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1498]),
        .S(self_sf7[1498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1499]),
        .S(self_sf7[1499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[149]),
        .S(self_sf7[149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[14].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[14]),
        .S(self_sf7[14]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1500]),
        .S(self_sf7[1500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1501]),
        .S(self_sf7[1501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1502]),
        .S(self_sf7[1502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1503]),
        .S(self_sf7[1503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1504]),
        .S(self_sf7[1504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1505]),
        .S(self_sf7[1505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1506]),
        .S(self_sf7[1506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1507]),
        .S(self_sf7[1507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1508]),
        .S(self_sf7[1508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1509]),
        .S(self_sf7[1509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[150]),
        .S(self_sf7[150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1510]),
        .S(self_sf7[1510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1511]),
        .S(self_sf7[1511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1512]),
        .S(self_sf7[1512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1513]),
        .S(self_sf7[1513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1514]),
        .S(self_sf7[1514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1515]),
        .S(self_sf7[1515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1516]),
        .S(self_sf7[1516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1517]),
        .S(self_sf7[1517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1518]),
        .S(self_sf7[1518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1519]),
        .S(self_sf7[1519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[151]),
        .S(self_sf7[151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1520]),
        .S(self_sf7[1520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1521]),
        .S(self_sf7[1521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1522]),
        .S(self_sf7[1522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1523]),
        .S(self_sf7[1523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1524]),
        .S(self_sf7[1524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1525]),
        .S(self_sf7[1525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1526]),
        .S(self_sf7[1526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1527]),
        .S(self_sf7[1527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1528]),
        .S(self_sf7[1528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1529]),
        .S(self_sf7[1529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[152]),
        .S(self_sf7[152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1530]),
        .S(self_sf7[1530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1531]),
        .S(self_sf7[1531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1532]),
        .S(self_sf7[1532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1533]),
        .S(self_sf7[1533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1534]),
        .S(self_sf7[1534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1535]),
        .S(self_sf7[1535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1536]),
        .S(self_sf7[1536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1537]),
        .S(self_sf7[1537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1538]),
        .S(self_sf7[1538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1539]),
        .S(self_sf7[1539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[153]),
        .S(self_sf7[153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1540]),
        .S(self_sf7[1540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1541]),
        .S(self_sf7[1541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1542]),
        .S(self_sf7[1542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1543]),
        .S(self_sf7[1543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1544]),
        .S(self_sf7[1544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1545]),
        .S(self_sf7[1545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1546]),
        .S(self_sf7[1546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1547]),
        .S(self_sf7[1547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1548]),
        .S(self_sf7[1548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1549]),
        .S(self_sf7[1549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[154]),
        .S(self_sf7[154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1550]),
        .S(self_sf7[1550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1551]),
        .S(self_sf7[1551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1552]),
        .S(self_sf7[1552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1553]),
        .S(self_sf7[1553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1554]),
        .S(self_sf7[1554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1555]),
        .S(self_sf7[1555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1556]),
        .S(self_sf7[1556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1557]),
        .S(self_sf7[1557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1558]),
        .S(self_sf7[1558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1559]),
        .S(self_sf7[1559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[155]),
        .S(self_sf7[155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1560]),
        .S(self_sf7[1560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1561]),
        .S(self_sf7[1561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1562]),
        .S(self_sf7[1562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1563]),
        .S(self_sf7[1563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1564]),
        .S(self_sf7[1564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1565]),
        .S(self_sf7[1565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1566]),
        .S(self_sf7[1566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1567]),
        .S(self_sf7[1567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1568]),
        .S(self_sf7[1568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1569]),
        .S(self_sf7[1569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[156]),
        .S(self_sf7[156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1570]),
        .S(self_sf7[1570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1571]),
        .S(self_sf7[1571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1572]),
        .S(self_sf7[1572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1573]),
        .S(self_sf7[1573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1574]),
        .S(self_sf7[1574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1575]),
        .S(self_sf7[1575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1576]),
        .S(self_sf7[1576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1577]),
        .S(self_sf7[1577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1578]),
        .S(self_sf7[1578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1579]),
        .S(self_sf7[1579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[157]),
        .S(self_sf7[157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1580]),
        .S(self_sf7[1580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1581]),
        .S(self_sf7[1581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1582]),
        .S(self_sf7[1582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1583]),
        .S(self_sf7[1583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1584]),
        .S(self_sf7[1584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1585]),
        .S(self_sf7[1585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1586]),
        .S(self_sf7[1586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1587]),
        .S(self_sf7[1587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1588]),
        .S(self_sf7[1588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1589]),
        .S(self_sf7[1589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[158]),
        .S(self_sf7[158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1590]),
        .S(self_sf7[1590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1591]),
        .S(self_sf7[1591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1592]),
        .S(self_sf7[1592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1593]),
        .S(self_sf7[1593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1594]),
        .S(self_sf7[1594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1595]),
        .S(self_sf7[1595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1596]),
        .S(self_sf7[1596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1597]),
        .S(self_sf7[1597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1598]),
        .S(self_sf7[1598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1599]),
        .S(self_sf7[1599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[159]),
        .S(self_sf7[159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[15].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[15]),
        .S(self_sf7[15]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1600]),
        .S(self_sf7[1600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1601]),
        .S(self_sf7[1601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1602]),
        .S(self_sf7[1602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1603]),
        .S(self_sf7[1603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1604]),
        .S(self_sf7[1604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1605]),
        .S(self_sf7[1605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1606]),
        .S(self_sf7[1606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1607]),
        .S(self_sf7[1607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1608]),
        .S(self_sf7[1608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1609]),
        .S(self_sf7[1609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[160]),
        .S(self_sf7[160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1610]),
        .S(self_sf7[1610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1611]),
        .S(self_sf7[1611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1612]),
        .S(self_sf7[1612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1613]),
        .S(self_sf7[1613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1614]),
        .S(self_sf7[1614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1615]),
        .S(self_sf7[1615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1616]),
        .S(self_sf7[1616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1617]),
        .S(self_sf7[1617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1618]),
        .S(self_sf7[1618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1619]),
        .S(self_sf7[1619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[161]),
        .S(self_sf7[161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1620]),
        .S(self_sf7[1620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1621]),
        .S(self_sf7[1621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1622]),
        .S(self_sf7[1622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1623]),
        .S(self_sf7[1623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1624]),
        .S(self_sf7[1624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1625]),
        .S(self_sf7[1625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1626]),
        .S(self_sf7[1626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1627]),
        .S(self_sf7[1627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1628]),
        .S(self_sf7[1628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1629]),
        .S(self_sf7[1629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[162]),
        .S(self_sf7[162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1630]),
        .S(self_sf7[1630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1631]),
        .S(self_sf7[1631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1632]),
        .S(self_sf7[1632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1633]),
        .S(self_sf7[1633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1634]),
        .S(self_sf7[1634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1635]),
        .S(self_sf7[1635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1636]),
        .S(self_sf7[1636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1637]),
        .S(self_sf7[1637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1638]),
        .S(self_sf7[1638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1639]),
        .S(self_sf7[1639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[163]),
        .S(self_sf7[163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1640]),
        .S(self_sf7[1640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1641]),
        .S(self_sf7[1641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1642]),
        .S(self_sf7[1642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1643]),
        .S(self_sf7[1643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1644]),
        .S(self_sf7[1644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1645]),
        .S(self_sf7[1645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1646]),
        .S(self_sf7[1646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1647]),
        .S(self_sf7[1647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1648]),
        .S(self_sf7[1648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1649]),
        .S(self_sf7[1649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[164]),
        .S(self_sf7[164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1650]),
        .S(self_sf7[1650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1651]),
        .S(self_sf7[1651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1652]),
        .S(self_sf7[1652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1653]),
        .S(self_sf7[1653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1654]),
        .S(self_sf7[1654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1655]),
        .S(self_sf7[1655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1656]),
        .S(self_sf7[1656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1657]),
        .S(self_sf7[1657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1658]),
        .S(self_sf7[1658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1659]),
        .S(self_sf7[1659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[165]),
        .S(self_sf7[165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1660]),
        .S(self_sf7[1660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1661]),
        .S(self_sf7[1661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1662]),
        .S(self_sf7[1662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1663]),
        .S(self_sf7[1663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1664]),
        .S(self_sf7[1664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1665]),
        .S(self_sf7[1665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1666]),
        .S(self_sf7[1666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1667]),
        .S(self_sf7[1667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1668]),
        .S(self_sf7[1668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1669]),
        .S(self_sf7[1669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[166]),
        .S(self_sf7[166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1670]),
        .S(self_sf7[1670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1671]),
        .S(self_sf7[1671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1672]),
        .S(self_sf7[1672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1673]),
        .S(self_sf7[1673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1674]),
        .S(self_sf7[1674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1675]),
        .S(self_sf7[1675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1676]),
        .S(self_sf7[1676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1677]),
        .S(self_sf7[1677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1678]),
        .S(self_sf7[1678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1679]),
        .S(self_sf7[1679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[167]),
        .S(self_sf7[167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1680]),
        .S(self_sf7[1680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1681]),
        .S(self_sf7[1681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1682]),
        .S(self_sf7[1682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1683]),
        .S(self_sf7[1683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1684]),
        .S(self_sf7[1684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1685]),
        .S(self_sf7[1685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1686]),
        .S(self_sf7[1686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1687]),
        .S(self_sf7[1687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1688]),
        .S(self_sf7[1688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1689]),
        .S(self_sf7[1689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[168]),
        .S(self_sf7[168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1690]),
        .S(self_sf7[1690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1691]),
        .S(self_sf7[1691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1692]),
        .S(self_sf7[1692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1693]),
        .S(self_sf7[1693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1694]),
        .S(self_sf7[1694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1695]),
        .S(self_sf7[1695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1696]),
        .S(self_sf7[1696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1697]),
        .S(self_sf7[1697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1698]),
        .S(self_sf7[1698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1699]),
        .S(self_sf7[1699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[169]),
        .S(self_sf7[169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[16].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[16]),
        .S(self_sf7[16]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1700]),
        .S(self_sf7[1700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1701]),
        .S(self_sf7[1701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1702]),
        .S(self_sf7[1702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1703]),
        .S(self_sf7[1703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1704]),
        .S(self_sf7[1704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1705]),
        .S(self_sf7[1705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1706]),
        .S(self_sf7[1706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1707]),
        .S(self_sf7[1707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1708]),
        .S(self_sf7[1708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1709]),
        .S(self_sf7[1709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[170]),
        .S(self_sf7[170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1710]),
        .S(self_sf7[1710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1711]),
        .S(self_sf7[1711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1712]),
        .S(self_sf7[1712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1713]),
        .S(self_sf7[1713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1714]),
        .S(self_sf7[1714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1715]),
        .S(self_sf7[1715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1716]),
        .S(self_sf7[1716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1717]),
        .S(self_sf7[1717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1718]),
        .S(self_sf7[1718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1719]),
        .S(self_sf7[1719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[171]),
        .S(self_sf7[171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1720]),
        .S(self_sf7[1720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1721]),
        .S(self_sf7[1721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1722]),
        .S(self_sf7[1722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1723]),
        .S(self_sf7[1723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1724]),
        .S(self_sf7[1724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1725]),
        .S(self_sf7[1725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1726]),
        .S(self_sf7[1726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1727]),
        .S(self_sf7[1727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1728]),
        .S(self_sf7[1728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1729]),
        .S(self_sf7[1729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[172]),
        .S(self_sf7[172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1730]),
        .S(self_sf7[1730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1731]),
        .S(self_sf7[1731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1732]),
        .S(self_sf7[1732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1733]),
        .S(self_sf7[1733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1734]),
        .S(self_sf7[1734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1735]),
        .S(self_sf7[1735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1736]),
        .S(self_sf7[1736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1737]),
        .S(self_sf7[1737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1738]),
        .S(self_sf7[1738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1739]),
        .S(self_sf7[1739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[173]),
        .S(self_sf7[173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1740]),
        .S(self_sf7[1740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1741]),
        .S(self_sf7[1741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1742]),
        .S(self_sf7[1742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1743]),
        .S(self_sf7[1743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1744]),
        .S(self_sf7[1744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1745]),
        .S(self_sf7[1745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1746]),
        .S(self_sf7[1746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1747]),
        .S(self_sf7[1747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1748]),
        .S(self_sf7[1748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1749]),
        .S(self_sf7[1749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[174]),
        .S(self_sf7[174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1750]),
        .S(self_sf7[1750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1751]),
        .S(self_sf7[1751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1752]),
        .S(self_sf7[1752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1753]),
        .S(self_sf7[1753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1754]),
        .S(self_sf7[1754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1755]),
        .S(self_sf7[1755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1756]),
        .S(self_sf7[1756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1757]),
        .S(self_sf7[1757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1758]),
        .S(self_sf7[1758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1759]),
        .S(self_sf7[1759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[175]),
        .S(self_sf7[175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1760]),
        .S(self_sf7[1760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1761]),
        .S(self_sf7[1761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1762]),
        .S(self_sf7[1762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1763]),
        .S(self_sf7[1763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1764]),
        .S(self_sf7[1764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1765]),
        .S(self_sf7[1765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1766]),
        .S(self_sf7[1766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1767]),
        .S(self_sf7[1767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1768]),
        .S(self_sf7[1768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1769]),
        .S(self_sf7[1769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[176]),
        .S(self_sf7[176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1770]),
        .S(self_sf7[1770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1771]),
        .S(self_sf7[1771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1772]),
        .S(self_sf7[1772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1773]),
        .S(self_sf7[1773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1774]),
        .S(self_sf7[1774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1775]),
        .S(self_sf7[1775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1776]),
        .S(self_sf7[1776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1777]),
        .S(self_sf7[1777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1778]),
        .S(self_sf7[1778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1779]),
        .S(self_sf7[1779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[177]),
        .S(self_sf7[177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1780]),
        .S(self_sf7[1780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1781]),
        .S(self_sf7[1781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1782]),
        .S(self_sf7[1782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1783]),
        .S(self_sf7[1783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1784]),
        .S(self_sf7[1784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1785]),
        .S(self_sf7[1785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1786]),
        .S(self_sf7[1786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1787]),
        .S(self_sf7[1787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1788]),
        .S(self_sf7[1788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1789]),
        .S(self_sf7[1789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[178]),
        .S(self_sf7[178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1790]),
        .S(self_sf7[1790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1791]),
        .S(self_sf7[1791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1792]),
        .S(self_sf7[1792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1793]),
        .S(self_sf7[1793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1794]),
        .S(self_sf7[1794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1795]),
        .S(self_sf7[1795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1796]),
        .S(self_sf7[1796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1797]),
        .S(self_sf7[1797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1798]),
        .S(self_sf7[1798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1799]),
        .S(self_sf7[1799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[179]),
        .S(self_sf7[179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[17].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[17]),
        .S(self_sf7[17]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[180]),
        .S(self_sf7[180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[181]),
        .S(self_sf7[181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[182]),
        .S(self_sf7[182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[183]),
        .S(self_sf7[183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[184]),
        .S(self_sf7[184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[185]),
        .S(self_sf7[185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[186]),
        .S(self_sf7[186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[187]),
        .S(self_sf7[187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[188]),
        .S(self_sf7[188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[189]),
        .S(self_sf7[189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[18].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[18]),
        .S(self_sf7[18]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[190]),
        .S(self_sf7[190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[191]),
        .S(self_sf7[191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[192]),
        .S(self_sf7[192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[193]),
        .S(self_sf7[193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[194]),
        .S(self_sf7[194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[195]),
        .S(self_sf7[195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[196]),
        .S(self_sf7[196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[197]),
        .S(self_sf7[197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[198]),
        .S(self_sf7[198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[199]),
        .S(self_sf7[199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[19].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[19]),
        .S(self_sf7[19]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1]),
        .S(info_sf7[1]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[200]),
        .S(self_sf7[200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[201]),
        .S(self_sf7[201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[202]),
        .S(self_sf7[202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[203]),
        .S(self_sf7[203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[204]),
        .S(self_sf7[204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[205]),
        .S(self_sf7[205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[206]),
        .S(self_sf7[206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[207]),
        .S(self_sf7[207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[208]),
        .S(self_sf7[208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[209]),
        .S(self_sf7[209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[20].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[20]),
        .S(self_sf7[20]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[210]),
        .S(self_sf7[210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[211]),
        .S(self_sf7[211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[212]),
        .S(self_sf7[212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[213]),
        .S(self_sf7[213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[214]),
        .S(self_sf7[214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[215]),
        .S(self_sf7[215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[216]),
        .S(self_sf7[216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[217]),
        .S(self_sf7[217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[218]),
        .S(self_sf7[218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[219]),
        .S(self_sf7[219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[21].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[21]),
        .S(self_sf7[21]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[220]),
        .S(self_sf7[220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[221]),
        .S(self_sf7[221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[222]),
        .S(self_sf7[222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[223]),
        .S(self_sf7[223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[224]),
        .S(self_sf7[224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[225]),
        .S(self_sf7[225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[226]),
        .S(self_sf7[226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[227]),
        .S(self_sf7[227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[228]),
        .S(self_sf7[228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[229]),
        .S(self_sf7[229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[22].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[22]),
        .S(self_sf7[22]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[230]),
        .S(self_sf7[230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[231]),
        .S(self_sf7[231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[232]),
        .S(self_sf7[232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[233]),
        .S(self_sf7[233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[234]),
        .S(self_sf7[234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[235]),
        .S(self_sf7[235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[236]),
        .S(self_sf7[236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[237]),
        .S(self_sf7[237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[238]),
        .S(self_sf7[238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[239]),
        .S(self_sf7[239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[23].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[23]),
        .S(self_sf7[23]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[240]),
        .S(self_sf7[240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[241]),
        .S(self_sf7[241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[242]),
        .S(self_sf7[242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[243]),
        .S(self_sf7[243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[244]),
        .S(self_sf7[244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[245]),
        .S(self_sf7[245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[246]),
        .S(self_sf7[246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[247]),
        .S(self_sf7[247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[248]),
        .S(self_sf7[248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[249]),
        .S(self_sf7[249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[24].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[24]),
        .S(self_sf7[24]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[250]),
        .S(self_sf7[250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[251]),
        .S(self_sf7[251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[252]),
        .S(self_sf7[252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[253]),
        .S(self_sf7[253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[254]),
        .S(self_sf7[254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[255]),
        .S(self_sf7[255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[256]),
        .S(self_sf7[256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[257]),
        .S(self_sf7[257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[258]),
        .S(self_sf7[258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[259]),
        .S(self_sf7[259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[25].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[25]),
        .S(self_sf7[25]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[260]),
        .S(self_sf7[260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[261]),
        .S(self_sf7[261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[262]),
        .S(self_sf7[262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[263]),
        .S(self_sf7[263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[264]),
        .S(self_sf7[264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[265]),
        .S(self_sf7[265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[266]),
        .S(self_sf7[266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[267]),
        .S(self_sf7[267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[268]),
        .S(self_sf7[268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[269]),
        .S(self_sf7[269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[26].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[26]),
        .S(self_sf7[26]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[270]),
        .S(self_sf7[270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[271]),
        .S(self_sf7[271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[272]),
        .S(self_sf7[272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[273]),
        .S(self_sf7[273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[274]),
        .S(self_sf7[274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[275]),
        .S(self_sf7[275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[276]),
        .S(self_sf7[276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[277]),
        .S(self_sf7[277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[278]),
        .S(self_sf7[278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[279]),
        .S(self_sf7[279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[27].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[27]),
        .S(self_sf7[27]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[280]),
        .S(self_sf7[280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[281]),
        .S(self_sf7[281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[282]),
        .S(self_sf7[282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[283]),
        .S(self_sf7[283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[284]),
        .S(self_sf7[284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[285]),
        .S(self_sf7[285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[286]),
        .S(self_sf7[286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[287]),
        .S(self_sf7[287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[288]),
        .S(self_sf7[288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[289]),
        .S(self_sf7[289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[28].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[28]),
        .S(self_sf7[28]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[290]),
        .S(self_sf7[290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[291]),
        .S(self_sf7[291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[292]),
        .S(self_sf7[292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[293]),
        .S(self_sf7[293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[294]),
        .S(self_sf7[294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[295]),
        .S(self_sf7[295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[296]),
        .S(self_sf7[296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[297]),
        .S(self_sf7[297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[298]),
        .S(self_sf7[298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[299]),
        .S(self_sf7[299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[29].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[29]),
        .S(self_sf7[29]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[2].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[2]),
        .S(info_sf7[2]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[300]),
        .S(self_sf7[300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[301]),
        .S(self_sf7[301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[302]),
        .S(self_sf7[302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[303]),
        .S(self_sf7[303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[304]),
        .S(self_sf7[304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[305]),
        .S(self_sf7[305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[306]),
        .S(self_sf7[306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[307]),
        .S(self_sf7[307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[308]),
        .S(self_sf7[308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[309]),
        .S(self_sf7[309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[30].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[30]),
        .S(self_sf7[30]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[310]),
        .S(self_sf7[310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[311]),
        .S(self_sf7[311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[312]),
        .S(self_sf7[312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[313]),
        .S(self_sf7[313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[314]),
        .S(self_sf7[314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[315]),
        .S(self_sf7[315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[316]),
        .S(self_sf7[316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[317]),
        .S(self_sf7[317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[318]),
        .S(self_sf7[318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[319]),
        .S(self_sf7[319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[31].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[31]),
        .S(self_sf7[31]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[320]),
        .S(self_sf7[320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[321]),
        .S(self_sf7[321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[322]),
        .S(self_sf7[322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[323]),
        .S(self_sf7[323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[324]),
        .S(self_sf7[324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[325]),
        .S(self_sf7[325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[326]),
        .S(self_sf7[326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[327]),
        .S(self_sf7[327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[328]),
        .S(self_sf7[328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[329]),
        .S(self_sf7[329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[32].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[32]),
        .S(self_sf7[32]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[330]),
        .S(self_sf7[330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[331]),
        .S(self_sf7[331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[332]),
        .S(self_sf7[332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[333]),
        .S(self_sf7[333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[334]),
        .S(self_sf7[334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[335]),
        .S(self_sf7[335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[336]),
        .S(self_sf7[336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[337]),
        .S(self_sf7[337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[338]),
        .S(self_sf7[338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[339]),
        .S(self_sf7[339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[33].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[33]),
        .S(self_sf7[33]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[340]),
        .S(self_sf7[340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[341]),
        .S(self_sf7[341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[342]),
        .S(self_sf7[342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[343]),
        .S(self_sf7[343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[344]),
        .S(self_sf7[344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[345]),
        .S(self_sf7[345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[346]),
        .S(self_sf7[346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[347]),
        .S(self_sf7[347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[348]),
        .S(self_sf7[348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[349]),
        .S(self_sf7[349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[34].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[34]),
        .S(self_sf7[34]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[350]),
        .S(self_sf7[350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[351]),
        .S(self_sf7[351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[352]),
        .S(self_sf7[352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[353]),
        .S(self_sf7[353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[354]),
        .S(self_sf7[354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[355]),
        .S(self_sf7[355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[356]),
        .S(self_sf7[356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[357]),
        .S(self_sf7[357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[358]),
        .S(self_sf7[358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[359]),
        .S(self_sf7[359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[35].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[35]),
        .S(self_sf7[35]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[360]),
        .S(self_sf7[360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[361]),
        .S(self_sf7[361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[362]),
        .S(self_sf7[362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[363]),
        .S(self_sf7[363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[364]),
        .S(self_sf7[364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[365]),
        .S(self_sf7[365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[366]),
        .S(self_sf7[366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[367]),
        .S(self_sf7[367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[368]),
        .S(self_sf7[368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[369]),
        .S(self_sf7[369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[36].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[36]),
        .S(self_sf7[36]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[370]),
        .S(self_sf7[370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[371]),
        .S(self_sf7[371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[372]),
        .S(self_sf7[372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[373]),
        .S(self_sf7[373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[374]),
        .S(self_sf7[374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[375]),
        .S(self_sf7[375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[376]),
        .S(self_sf7[376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[377]),
        .S(self_sf7[377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[378]),
        .S(self_sf7[378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[379]),
        .S(self_sf7[379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[37].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[37]),
        .S(self_sf7[37]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[380]),
        .S(self_sf7[380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[381]),
        .S(self_sf7[381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[382]),
        .S(self_sf7[382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[383]),
        .S(self_sf7[383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[384]),
        .S(self_sf7[384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[385]),
        .S(self_sf7[385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[386]),
        .S(self_sf7[386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[387]),
        .S(self_sf7[387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[388]),
        .S(self_sf7[388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[389]),
        .S(self_sf7[389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[38].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[38]),
        .S(self_sf7[38]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[390]),
        .S(self_sf7[390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[391]),
        .S(self_sf7[391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[392]),
        .S(self_sf7[392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[393]),
        .S(self_sf7[393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[394]),
        .S(self_sf7[394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[395]),
        .S(self_sf7[395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[396]),
        .S(self_sf7[396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[397]),
        .S(self_sf7[397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[398]),
        .S(self_sf7[398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[399]),
        .S(self_sf7[399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[39].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[39]),
        .S(self_sf7[39]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[3].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[3]),
        .S(info_sf7[3]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[400]),
        .S(self_sf7[400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[401]),
        .S(self_sf7[401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[402]),
        .S(self_sf7[402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[403]),
        .S(self_sf7[403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[404]),
        .S(self_sf7[404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[405]),
        .S(self_sf7[405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[406]),
        .S(self_sf7[406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[407]),
        .S(self_sf7[407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[408]),
        .S(self_sf7[408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[409]),
        .S(self_sf7[409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[40].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[40]),
        .S(self_sf7[40]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[410]),
        .S(self_sf7[410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[411]),
        .S(self_sf7[411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[412]),
        .S(self_sf7[412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[413]),
        .S(self_sf7[413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[414]),
        .S(self_sf7[414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[415]),
        .S(self_sf7[415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[416]),
        .S(self_sf7[416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[417]),
        .S(self_sf7[417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[418]),
        .S(self_sf7[418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[419]),
        .S(self_sf7[419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[41].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[41]),
        .S(self_sf7[41]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[420]),
        .S(self_sf7[420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[421]),
        .S(self_sf7[421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[422]),
        .S(self_sf7[422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[423]),
        .S(self_sf7[423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[424]),
        .S(self_sf7[424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[425]),
        .S(self_sf7[425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[426]),
        .S(self_sf7[426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[427]),
        .S(self_sf7[427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[428]),
        .S(self_sf7[428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[429]),
        .S(self_sf7[429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[42].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[42]),
        .S(self_sf7[42]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[430]),
        .S(self_sf7[430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[431]),
        .S(self_sf7[431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[432]),
        .S(self_sf7[432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[433]),
        .S(self_sf7[433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[434]),
        .S(self_sf7[434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[435]),
        .S(self_sf7[435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[436]),
        .S(self_sf7[436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[437]),
        .S(self_sf7[437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[438]),
        .S(self_sf7[438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[439]),
        .S(self_sf7[439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[43].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[43]),
        .S(self_sf7[43]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[440]),
        .S(self_sf7[440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[441]),
        .S(self_sf7[441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[442]),
        .S(self_sf7[442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[443]),
        .S(self_sf7[443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[444]),
        .S(self_sf7[444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[445]),
        .S(self_sf7[445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[446]),
        .S(self_sf7[446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[447]),
        .S(self_sf7[447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[448]),
        .S(self_sf7[448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[449]),
        .S(self_sf7[449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[44].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[44]),
        .S(self_sf7[44]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[450]),
        .S(self_sf7[450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[451]),
        .S(self_sf7[451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[452]),
        .S(self_sf7[452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[453]),
        .S(self_sf7[453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[454]),
        .S(self_sf7[454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[455]),
        .S(self_sf7[455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[456]),
        .S(self_sf7[456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[457]),
        .S(self_sf7[457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[458]),
        .S(self_sf7[458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[459]),
        .S(self_sf7[459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[45].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[45]),
        .S(self_sf7[45]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[460]),
        .S(self_sf7[460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[461]),
        .S(self_sf7[461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[462]),
        .S(self_sf7[462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[463]),
        .S(self_sf7[463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[464]),
        .S(self_sf7[464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[465]),
        .S(self_sf7[465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[466]),
        .S(self_sf7[466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[467]),
        .S(self_sf7[467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[468]),
        .S(self_sf7[468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[469]),
        .S(self_sf7[469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[46].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[46]),
        .S(self_sf7[46]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[470]),
        .S(self_sf7[470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[471]),
        .S(self_sf7[471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[472]),
        .S(self_sf7[472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[473]),
        .S(self_sf7[473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[474]),
        .S(self_sf7[474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[475]),
        .S(self_sf7[475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[476]),
        .S(self_sf7[476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[477]),
        .S(self_sf7[477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[478]),
        .S(self_sf7[478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[479]),
        .S(self_sf7[479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[47].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[47]),
        .S(self_sf7[47]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[480]),
        .S(self_sf7[480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[481]),
        .S(self_sf7[481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[482]),
        .S(self_sf7[482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[483]),
        .S(self_sf7[483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[484]),
        .S(self_sf7[484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[485]),
        .S(self_sf7[485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[486]),
        .S(self_sf7[486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[487]),
        .S(self_sf7[487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[488]),
        .S(self_sf7[488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[489]),
        .S(self_sf7[489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[48].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[48]),
        .S(self_sf7[48]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[490]),
        .S(self_sf7[490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[491]),
        .S(self_sf7[491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[492]),
        .S(self_sf7[492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[493]),
        .S(self_sf7[493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[494]),
        .S(self_sf7[494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[495]),
        .S(self_sf7[495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[496]),
        .S(self_sf7[496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[497]),
        .S(self_sf7[497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[498]),
        .S(self_sf7[498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[499]),
        .S(self_sf7[499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[49].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[49]),
        .S(self_sf7[49]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[4].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[4]),
        .S(info_sf7[4]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[500]),
        .S(self_sf7[500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[501]),
        .S(self_sf7[501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[502]),
        .S(self_sf7[502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[503]),
        .S(self_sf7[503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[504]),
        .S(self_sf7[504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[505]),
        .S(self_sf7[505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[506]),
        .S(self_sf7[506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[507]),
        .S(self_sf7[507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[508]),
        .S(self_sf7[508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[509]),
        .S(self_sf7[509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[50].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[50]),
        .S(self_sf7[50]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[510]),
        .S(self_sf7[510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[511]),
        .S(self_sf7[511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[512]),
        .S(self_sf7[512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[513]),
        .S(self_sf7[513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[514]),
        .S(self_sf7[514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[515]),
        .S(self_sf7[515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[516]),
        .S(self_sf7[516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[517]),
        .S(self_sf7[517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[518]),
        .S(self_sf7[518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[519]),
        .S(self_sf7[519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[51].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[51]),
        .S(self_sf7[51]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[520]),
        .S(self_sf7[520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[521]),
        .S(self_sf7[521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[522]),
        .S(self_sf7[522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[523]),
        .S(self_sf7[523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[524]),
        .S(self_sf7[524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[525]),
        .S(self_sf7[525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[526]),
        .S(self_sf7[526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[527]),
        .S(self_sf7[527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[528]),
        .S(self_sf7[528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[529]),
        .S(self_sf7[529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[52].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[52]),
        .S(self_sf7[52]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[530]),
        .S(self_sf7[530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[531]),
        .S(self_sf7[531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[532]),
        .S(self_sf7[532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[533]),
        .S(self_sf7[533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[534]),
        .S(self_sf7[534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[535]),
        .S(self_sf7[535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[536]),
        .S(self_sf7[536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[537]),
        .S(self_sf7[537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[538]),
        .S(self_sf7[538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[539]),
        .S(self_sf7[539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[53].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[53]),
        .S(self_sf7[53]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[540]),
        .S(self_sf7[540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[541]),
        .S(self_sf7[541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[542]),
        .S(self_sf7[542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[543]),
        .S(self_sf7[543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[544]),
        .S(self_sf7[544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[545]),
        .S(self_sf7[545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[546]),
        .S(self_sf7[546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[547]),
        .S(self_sf7[547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[548]),
        .S(self_sf7[548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[549]),
        .S(self_sf7[549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[54].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[54]),
        .S(self_sf7[54]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[550]),
        .S(self_sf7[550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[551]),
        .S(self_sf7[551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[552]),
        .S(self_sf7[552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[553]),
        .S(self_sf7[553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[554]),
        .S(self_sf7[554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[555]),
        .S(self_sf7[555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[556]),
        .S(self_sf7[556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[557]),
        .S(self_sf7[557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[558]),
        .S(self_sf7[558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[559]),
        .S(self_sf7[559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[55].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[55]),
        .S(self_sf7[55]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[560]),
        .S(self_sf7[560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[561]),
        .S(self_sf7[561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[562]),
        .S(self_sf7[562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[563]),
        .S(self_sf7[563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[564]),
        .S(self_sf7[564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[565]),
        .S(self_sf7[565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[566]),
        .S(self_sf7[566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[567]),
        .S(self_sf7[567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[568]),
        .S(self_sf7[568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[569]),
        .S(self_sf7[569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[56].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[56]),
        .S(self_sf7[56]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[570]),
        .S(self_sf7[570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[571]),
        .S(self_sf7[571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[572]),
        .S(self_sf7[572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[573]),
        .S(self_sf7[573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[574]),
        .S(self_sf7[574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[575]),
        .S(self_sf7[575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[576]),
        .S(self_sf7[576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[577]),
        .S(self_sf7[577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[578]),
        .S(self_sf7[578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[579]),
        .S(self_sf7[579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[57].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[57]),
        .S(self_sf7[57]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[580]),
        .S(self_sf7[580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[581]),
        .S(self_sf7[581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[582]),
        .S(self_sf7[582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[583]),
        .S(self_sf7[583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[584]),
        .S(self_sf7[584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[585]),
        .S(self_sf7[585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[586]),
        .S(self_sf7[586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[587]),
        .S(self_sf7[587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[588]),
        .S(self_sf7[588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[589]),
        .S(self_sf7[589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[58].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[58]),
        .S(self_sf7[58]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[590]),
        .S(self_sf7[590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[591]),
        .S(self_sf7[591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[592]),
        .S(self_sf7[592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[593]),
        .S(self_sf7[593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[594]),
        .S(self_sf7[594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[595]),
        .S(self_sf7[595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[596]),
        .S(self_sf7[596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[597]),
        .S(self_sf7[597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[598]),
        .S(self_sf7[598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[599]),
        .S(self_sf7[599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[59].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[59]),
        .S(self_sf7[59]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[5].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[5]),
        .S(info_sf7[5]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[600]),
        .S(self_sf7[600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[601]),
        .S(self_sf7[601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[602]),
        .S(self_sf7[602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[603]),
        .S(self_sf7[603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[604]),
        .S(self_sf7[604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[605]),
        .S(self_sf7[605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[606]),
        .S(self_sf7[606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[607]),
        .S(self_sf7[607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[608]),
        .S(self_sf7[608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[609]),
        .S(self_sf7[609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[60].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[60]),
        .S(self_sf7[60]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[610]),
        .S(self_sf7[610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[611]),
        .S(self_sf7[611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[612]),
        .S(self_sf7[612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[613]),
        .S(self_sf7[613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[614]),
        .S(self_sf7[614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[615]),
        .S(self_sf7[615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[616]),
        .S(self_sf7[616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[617]),
        .S(self_sf7[617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[618]),
        .S(self_sf7[618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[619]),
        .S(self_sf7[619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[61].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[61]),
        .S(self_sf7[61]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[620]),
        .S(self_sf7[620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[621]),
        .S(self_sf7[621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[622]),
        .S(self_sf7[622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[623]),
        .S(self_sf7[623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[624]),
        .S(self_sf7[624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[625]),
        .S(self_sf7[625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[626]),
        .S(self_sf7[626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[627]),
        .S(self_sf7[627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[628]),
        .S(self_sf7[628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[629]),
        .S(self_sf7[629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[62].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[62]),
        .S(self_sf7[62]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[630]),
        .S(self_sf7[630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[631]),
        .S(self_sf7[631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[632]),
        .S(self_sf7[632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[633]),
        .S(self_sf7[633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[634]),
        .S(self_sf7[634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[635]),
        .S(self_sf7[635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[636]),
        .S(self_sf7[636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[637]),
        .S(self_sf7[637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[638]),
        .S(self_sf7[638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[639]),
        .S(self_sf7[639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[63].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[63]),
        .S(self_sf7[63]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[640]),
        .S(self_sf7[640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[641]),
        .S(self_sf7[641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[642]),
        .S(self_sf7[642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[643]),
        .S(self_sf7[643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[644]),
        .S(self_sf7[644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[645]),
        .S(self_sf7[645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[646]),
        .S(self_sf7[646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[647]),
        .S(self_sf7[647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[648]),
        .S(self_sf7[648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[649]),
        .S(self_sf7[649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[64].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[64]),
        .S(self_sf7[64]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[650]),
        .S(self_sf7[650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[651]),
        .S(self_sf7[651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[652]),
        .S(self_sf7[652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[653]),
        .S(self_sf7[653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[654]),
        .S(self_sf7[654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[655]),
        .S(self_sf7[655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[656]),
        .S(self_sf7[656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[657]),
        .S(self_sf7[657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[658]),
        .S(self_sf7[658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[659]),
        .S(self_sf7[659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[65].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[65]),
        .S(self_sf7[65]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[660]),
        .S(self_sf7[660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[661]),
        .S(self_sf7[661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[662]),
        .S(self_sf7[662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[663]),
        .S(self_sf7[663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[664]),
        .S(self_sf7[664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[665]),
        .S(self_sf7[665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[666]),
        .S(self_sf7[666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[667]),
        .S(self_sf7[667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[668]),
        .S(self_sf7[668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[669]),
        .S(self_sf7[669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[66].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[66]),
        .S(self_sf7[66]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[670]),
        .S(self_sf7[670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[671]),
        .S(self_sf7[671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[672]),
        .S(self_sf7[672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[673]),
        .S(self_sf7[673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[674]),
        .S(self_sf7[674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[675]),
        .S(self_sf7[675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[676]),
        .S(self_sf7[676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[677]),
        .S(self_sf7[677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[678]),
        .S(self_sf7[678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[679]),
        .S(self_sf7[679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[67].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[67]),
        .S(self_sf7[67]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[680]),
        .S(self_sf7[680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[681]),
        .S(self_sf7[681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[682]),
        .S(self_sf7[682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[683]),
        .S(self_sf7[683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[684]),
        .S(self_sf7[684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[685]),
        .S(self_sf7[685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[686]),
        .S(self_sf7[686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[687]),
        .S(self_sf7[687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[688]),
        .S(self_sf7[688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[689]),
        .S(self_sf7[689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[68].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[68]),
        .S(self_sf7[68]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[690]),
        .S(self_sf7[690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[691]),
        .S(self_sf7[691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[692]),
        .S(self_sf7[692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[693]),
        .S(self_sf7[693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[694]),
        .S(self_sf7[694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[695]),
        .S(self_sf7[695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[696]),
        .S(self_sf7[696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[697]),
        .S(self_sf7[697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[698]),
        .S(self_sf7[698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[699]),
        .S(self_sf7[699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[69].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[69]),
        .S(self_sf7[69]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[6].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[6]),
        .S(info_sf7[6]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[700]),
        .S(self_sf7[700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[701]),
        .S(self_sf7[701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[702]),
        .S(self_sf7[702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[703]),
        .S(self_sf7[703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[704]),
        .S(self_sf7[704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[705]),
        .S(self_sf7[705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[706]),
        .S(self_sf7[706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[707]),
        .S(self_sf7[707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[708]),
        .S(self_sf7[708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[709]),
        .S(self_sf7[709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[70].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[70]),
        .S(self_sf7[70]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[710]),
        .S(self_sf7[710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[711]),
        .S(self_sf7[711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[712]),
        .S(self_sf7[712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[713]),
        .S(self_sf7[713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[714]),
        .S(self_sf7[714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[715]),
        .S(self_sf7[715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[716]),
        .S(self_sf7[716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[717]),
        .S(self_sf7[717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[718]),
        .S(self_sf7[718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[719]),
        .S(self_sf7[719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[71].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[71]),
        .S(self_sf7[71]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[720]),
        .S(self_sf7[720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[721]),
        .S(self_sf7[721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[722]),
        .S(self_sf7[722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[723]),
        .S(self_sf7[723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[724]),
        .S(self_sf7[724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[725]),
        .S(self_sf7[725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[726]),
        .S(self_sf7[726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[727]),
        .S(self_sf7[727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[728]),
        .S(self_sf7[728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[729]),
        .S(self_sf7[729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[72].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[72]),
        .S(self_sf7[72]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[730]),
        .S(self_sf7[730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[731]),
        .S(self_sf7[731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[732]),
        .S(self_sf7[732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[733]),
        .S(self_sf7[733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[734]),
        .S(self_sf7[734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[735]),
        .S(self_sf7[735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[736]),
        .S(self_sf7[736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[737]),
        .S(self_sf7[737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[738]),
        .S(self_sf7[738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[739]),
        .S(self_sf7[739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[73].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[73]),
        .S(self_sf7[73]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[740]),
        .S(self_sf7[740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[741]),
        .S(self_sf7[741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[742]),
        .S(self_sf7[742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[743]),
        .S(self_sf7[743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[744]),
        .S(self_sf7[744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[745]),
        .S(self_sf7[745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[746]),
        .S(self_sf7[746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[747]),
        .S(self_sf7[747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[748]),
        .S(self_sf7[748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[749]),
        .S(self_sf7[749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[74].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[74]),
        .S(self_sf7[74]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[750]),
        .S(self_sf7[750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[751]),
        .S(self_sf7[751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[752]),
        .S(self_sf7[752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[753]),
        .S(self_sf7[753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[754]),
        .S(self_sf7[754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[755]),
        .S(self_sf7[755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[756]),
        .S(self_sf7[756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[757]),
        .S(self_sf7[757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[758]),
        .S(self_sf7[758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[759]),
        .S(self_sf7[759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[75].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[75]),
        .S(self_sf7[75]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[760]),
        .S(self_sf7[760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[761]),
        .S(self_sf7[761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[762]),
        .S(self_sf7[762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[763]),
        .S(self_sf7[763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[764]),
        .S(self_sf7[764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[765]),
        .S(self_sf7[765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[766]),
        .S(self_sf7[766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[767]),
        .S(self_sf7[767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[768]),
        .S(self_sf7[768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[769]),
        .S(self_sf7[769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[76].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[76]),
        .S(self_sf7[76]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[770]),
        .S(self_sf7[770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[771]),
        .S(self_sf7[771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[772]),
        .S(self_sf7[772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[773]),
        .S(self_sf7[773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[774]),
        .S(self_sf7[774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[775]),
        .S(self_sf7[775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[776]),
        .S(self_sf7[776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[777]),
        .S(self_sf7[777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[778]),
        .S(self_sf7[778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[779]),
        .S(self_sf7[779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[77].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[77]),
        .S(self_sf7[77]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[780]),
        .S(self_sf7[780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[781]),
        .S(self_sf7[781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[782]),
        .S(self_sf7[782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[783]),
        .S(self_sf7[783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[784]),
        .S(self_sf7[784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[785]),
        .S(self_sf7[785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[786]),
        .S(self_sf7[786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[787]),
        .S(self_sf7[787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[788]),
        .S(self_sf7[788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[789]),
        .S(self_sf7[789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[78].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[78]),
        .S(self_sf7[78]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[790]),
        .S(self_sf7[790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[791]),
        .S(self_sf7[791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[792]),
        .S(self_sf7[792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[793]),
        .S(self_sf7[793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[794]),
        .S(self_sf7[794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[795]),
        .S(self_sf7[795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[796]),
        .S(self_sf7[796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[797]),
        .S(self_sf7[797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[798]),
        .S(self_sf7[798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[799]),
        .S(self_sf7[799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[79].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[79]),
        .S(self_sf7[79]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[7].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[7]),
        .S(info_sf7[7]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[800].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[800]),
        .S(self_sf7[800]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[801].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[801]),
        .S(self_sf7[801]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[802].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[802]),
        .S(self_sf7[802]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[803].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[803]),
        .S(self_sf7[803]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[804].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[804]),
        .S(self_sf7[804]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[805].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[805]),
        .S(self_sf7[805]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[806].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[806]),
        .S(self_sf7[806]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[807].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[807]),
        .S(self_sf7[807]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[808].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[808]),
        .S(self_sf7[808]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[809].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[809]),
        .S(self_sf7[809]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[80].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[80]),
        .S(self_sf7[80]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[810].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[810]),
        .S(self_sf7[810]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[811].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[811]),
        .S(self_sf7[811]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[812].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[812]),
        .S(self_sf7[812]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[813].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[813]),
        .S(self_sf7[813]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[814].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[814]),
        .S(self_sf7[814]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[815].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[815]),
        .S(self_sf7[815]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[816].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[816]),
        .S(self_sf7[816]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[817].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[817]),
        .S(self_sf7[817]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[818].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[818]),
        .S(self_sf7[818]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[819].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[819]),
        .S(self_sf7[819]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[81].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[81]),
        .S(self_sf7[81]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[820].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[820]),
        .S(self_sf7[820]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[821].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[821]),
        .S(self_sf7[821]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[822].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[822]),
        .S(self_sf7[822]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[823].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[823]),
        .S(self_sf7[823]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[824].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[824]),
        .S(self_sf7[824]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[825].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[825]),
        .S(self_sf7[825]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[826].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[826]),
        .S(self_sf7[826]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[827].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[827]),
        .S(self_sf7[827]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[828].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[828]),
        .S(self_sf7[828]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[829].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[829]),
        .S(self_sf7[829]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[82].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[82]),
        .S(self_sf7[82]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[830].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[830]),
        .S(self_sf7[830]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[831].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[831]),
        .S(self_sf7[831]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[832].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[832]),
        .S(self_sf7[832]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[833].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[833]),
        .S(self_sf7[833]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[834].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[834]),
        .S(self_sf7[834]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[835].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[835]),
        .S(self_sf7[835]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[836].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[836]),
        .S(self_sf7[836]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[837].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[837]),
        .S(self_sf7[837]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[838].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[838]),
        .S(self_sf7[838]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[839].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[839]),
        .S(self_sf7[839]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[83].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[83]),
        .S(self_sf7[83]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[840].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[840]),
        .S(self_sf7[840]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[841].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[841]),
        .S(self_sf7[841]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[842].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[842]),
        .S(self_sf7[842]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[843].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[843]),
        .S(self_sf7[843]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[844].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[844]),
        .S(self_sf7[844]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[845].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[845]),
        .S(self_sf7[845]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[846].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[846]),
        .S(self_sf7[846]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[847].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[847]),
        .S(self_sf7[847]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[848].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[848]),
        .S(self_sf7[848]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[849].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[849]),
        .S(self_sf7[849]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[84].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[84]),
        .S(self_sf7[84]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[850].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[850]),
        .S(self_sf7[850]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[851].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[851]),
        .S(self_sf7[851]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[852].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[852]),
        .S(self_sf7[852]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[853].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[853]),
        .S(self_sf7[853]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[854].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[854]),
        .S(self_sf7[854]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[855].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[855]),
        .S(self_sf7[855]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[856].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[856]),
        .S(self_sf7[856]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[857].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[857]),
        .S(self_sf7[857]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[858].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[858]),
        .S(self_sf7[858]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[859].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[859]),
        .S(self_sf7[859]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[85].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[85]),
        .S(self_sf7[85]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[860].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[860]),
        .S(self_sf7[860]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[861].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[861]),
        .S(self_sf7[861]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[862].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[862]),
        .S(self_sf7[862]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[863].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[863]),
        .S(self_sf7[863]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[864].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[864]),
        .S(self_sf7[864]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[865].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[865]),
        .S(self_sf7[865]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[866].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[866]),
        .S(self_sf7[866]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[867].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[867]),
        .S(self_sf7[867]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[868].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[868]),
        .S(self_sf7[868]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[869].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[869]),
        .S(self_sf7[869]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[86].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[86]),
        .S(self_sf7[86]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[870].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[870]),
        .S(self_sf7[870]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[871].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[871]),
        .S(self_sf7[871]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[872].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[872]),
        .S(self_sf7[872]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[873].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[873]),
        .S(self_sf7[873]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[874].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[874]),
        .S(self_sf7[874]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[875].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[875]),
        .S(self_sf7[875]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[876].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[876]),
        .S(self_sf7[876]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[877].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[877]),
        .S(self_sf7[877]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[878].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[878]),
        .S(self_sf7[878]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[879].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[879]),
        .S(self_sf7[879]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[87].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[87]),
        .S(self_sf7[87]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[880].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[880]),
        .S(self_sf7[880]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[881].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[881]),
        .S(self_sf7[881]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[882].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[882]),
        .S(self_sf7[882]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[883].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[883]),
        .S(self_sf7[883]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[884].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[884]),
        .S(self_sf7[884]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[885].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[885]),
        .S(self_sf7[885]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[886].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[886]),
        .S(self_sf7[886]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[887].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[887]),
        .S(self_sf7[887]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[888].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[888]),
        .S(self_sf7[888]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[889].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[889]),
        .S(self_sf7[889]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[88].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[88]),
        .S(self_sf7[88]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[890].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[890]),
        .S(self_sf7[890]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[891].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[891]),
        .S(self_sf7[891]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[892].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[892]),
        .S(self_sf7[892]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[893].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[893]),
        .S(self_sf7[893]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[894].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[894]),
        .S(self_sf7[894]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[895].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[895]),
        .S(self_sf7[895]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[896].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[896]),
        .S(self_sf7[896]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[897].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[897]),
        .S(self_sf7[897]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[898].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[898]),
        .S(self_sf7[898]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[899].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[899]),
        .S(self_sf7[899]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[89].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[89]),
        .S(self_sf7[89]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[8].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[8]),
        .S(self_sf7[8]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[900].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[900]),
        .S(self_sf7[900]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[901].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[901]),
        .S(self_sf7[901]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[902].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[902]),
        .S(self_sf7[902]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[903].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[903]),
        .S(self_sf7[903]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[904].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[904]),
        .S(self_sf7[904]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[905].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[905]),
        .S(self_sf7[905]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[906].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[906]),
        .S(self_sf7[906]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[907].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[907]),
        .S(self_sf7[907]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[908].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[908]),
        .S(self_sf7[908]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[909].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[909]),
        .S(self_sf7[909]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[90].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[90]),
        .S(self_sf7[90]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[910].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[910]),
        .S(self_sf7[910]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[911].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[911]),
        .S(self_sf7[911]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[912].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[912]),
        .S(self_sf7[912]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[913].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[913]),
        .S(self_sf7[913]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[914].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[914]),
        .S(self_sf7[914]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[915].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[915]),
        .S(self_sf7[915]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[916].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[916]),
        .S(self_sf7[916]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[917].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[917]),
        .S(self_sf7[917]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[918].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[918]),
        .S(self_sf7[918]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[919].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[919]),
        .S(self_sf7[919]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[91].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[91]),
        .S(self_sf7[91]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[920].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[920]),
        .S(self_sf7[920]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[921].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[921]),
        .S(self_sf7[921]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[922].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[922]),
        .S(self_sf7[922]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[923].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[923]),
        .S(self_sf7[923]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[924].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[924]),
        .S(self_sf7[924]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[925].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[925]),
        .S(self_sf7[925]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[926].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[926]),
        .S(self_sf7[926]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[927].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[927]),
        .S(self_sf7[927]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[928].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[928]),
        .S(self_sf7[928]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[929].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[929]),
        .S(self_sf7[929]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[92].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[92]),
        .S(self_sf7[92]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[930].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[930]),
        .S(self_sf7[930]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[931].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[931]),
        .S(self_sf7[931]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[932].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[932]),
        .S(self_sf7[932]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[933].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[933]),
        .S(self_sf7[933]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[934].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[934]),
        .S(self_sf7[934]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[935].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[935]),
        .S(self_sf7[935]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[936].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[936]),
        .S(self_sf7[936]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[937].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[937]),
        .S(self_sf7[937]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[938].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[938]),
        .S(self_sf7[938]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[939].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[939]),
        .S(self_sf7[939]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[93].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[93]),
        .S(self_sf7[93]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[940].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[940]),
        .S(self_sf7[940]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[941].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[941]),
        .S(self_sf7[941]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[942].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[942]),
        .S(self_sf7[942]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[943].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[943]),
        .S(self_sf7[943]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[944].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[944]),
        .S(self_sf7[944]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[945].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[945]),
        .S(self_sf7[945]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[946].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[946]),
        .S(self_sf7[946]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[947].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[947]),
        .S(self_sf7[947]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[948].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[948]),
        .S(self_sf7[948]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[949].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[949]),
        .S(self_sf7[949]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[94].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[94]),
        .S(self_sf7[94]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[950].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[950]),
        .S(self_sf7[950]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[951].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[951]),
        .S(self_sf7[951]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[952].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[952]),
        .S(self_sf7[952]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[953].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[953]),
        .S(self_sf7[953]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[954].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[954]),
        .S(self_sf7[954]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[955].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[955]),
        .S(self_sf7[955]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[956].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[956]),
        .S(self_sf7[956]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[957].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[957]),
        .S(self_sf7[957]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[958].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[958]),
        .S(self_sf7[958]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[959].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[959]),
        .S(self_sf7[959]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[95].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[95]),
        .S(self_sf7[95]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[960].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[960]),
        .S(self_sf7[960]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[961].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[961]),
        .S(self_sf7[961]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[962].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[962]),
        .S(self_sf7[962]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[963].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[963]),
        .S(self_sf7[963]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[964].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[964]),
        .S(self_sf7[964]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[965].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[965]),
        .S(self_sf7[965]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[966].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[966]),
        .S(self_sf7[966]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[967].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[967]),
        .S(self_sf7[967]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[968].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[968]),
        .S(self_sf7[968]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[969].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[969]),
        .S(self_sf7[969]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[96].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[96]),
        .S(self_sf7[96]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[970].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[970]),
        .S(self_sf7[970]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[971].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[971]),
        .S(self_sf7[971]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[972].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[972]),
        .S(self_sf7[972]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[973].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[973]),
        .S(self_sf7[973]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[974].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[974]),
        .S(self_sf7[974]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[975].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[975]),
        .S(self_sf7[975]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[976].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[976]),
        .S(self_sf7[976]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[977].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[977]),
        .S(self_sf7[977]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[978].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[978]),
        .S(self_sf7[978]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[979].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[979]),
        .S(self_sf7[979]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[97].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[97]),
        .S(self_sf7[97]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[980].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[980]),
        .S(self_sf7[980]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[981].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[981]),
        .S(self_sf7[981]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[982].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[982]),
        .S(self_sf7[982]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[983].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[983]),
        .S(self_sf7[983]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[984].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[984]),
        .S(self_sf7[984]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[985].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[985]),
        .S(self_sf7[985]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[986].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[986]),
        .S(self_sf7[986]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[987].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[987]),
        .S(self_sf7[987]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[988].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[988]),
        .S(self_sf7[988]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[989].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[989]),
        .S(self_sf7[989]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[98].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[98]),
        .S(self_sf7[98]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[990].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[990]),
        .S(self_sf7[990]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[991].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[991]),
        .S(self_sf7[991]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[992].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[992]),
        .S(self_sf7[992]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[993].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[993]),
        .S(self_sf7[993]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[994].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[994]),
        .S(self_sf7[994]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[995].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[995]),
        .S(self_sf7[995]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[996].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[996]),
        .S(self_sf7[996]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[997].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[997]),
        .S(self_sf7[997]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[998].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[998]),
        .S(self_sf7[998]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[999].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[999]),
        .S(self_sf7[999]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[99].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[99]),
        .S(self_sf7[99]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[9].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[9]),
        .S(self_sf7[9]));
  (* BOX_TYPE = "black_box" *) 
  MUXF8 \activity_ROsf8[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf8[0]),
        .S(self_sf8[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF9 \activity_ROsf9[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf9[0]),
        .S(self_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_0
       (.I0(1'b0),
        .O(self_sf7[1802]));
  LUT1 #(
    .INIT(2'h2)) 
    i_1
       (.I0(1'b0),
        .O(self_sf7[1801]));
  LUT1 #(
    .INIT(2'h2)) 
    i_10
       (.I0(1'b0),
        .O(info_sf8[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_11
       (.I0(1'b0),
        .O(info_sf8[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_12
       (.I0(1'b0),
        .O(info_sf8[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_13
       (.I0(1'b0),
        .O(info_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_14
       (.I0(1'b0),
        .O(info_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_15
       (.I0(1'b0),
        .O(info_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_16
       (.I0(1'b0),
        .O(info_sf8[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_17
       (.I0(1'b0),
        .O(info_sf9[7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_18
       (.I0(1'b0),
        .O(info_sf9[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_19
       (.I0(1'b0),
        .O(info_sf9[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_2
       (.I0(1'b0),
        .O(self_sf7[1800]));
  LUT1 #(
    .INIT(2'h2)) 
    i_20
       (.I0(1'b0),
        .O(info_sf9[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_21
       (.I0(1'b0),
        .O(info_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_22
       (.I0(1'b0),
        .O(info_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_23
       (.I0(1'b0),
        .O(info_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_24
       (.I0(1'b0),
        .O(info_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_3
       (.I0(1'b0),
        .O(self_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_4
       (.I0(1'b0),
        .O(self_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_5
       (.I0(1'b0),
        .O(self_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_6
       (.I0(1'b0),
        .O(self_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_7
       (.I0(1'b0),
        .O(self_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_8
       (.I0(1'b0),
        .O(self_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_9
       (.I0(1'b0),
        .O(info_sf8[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst
       (.I0(self_sf7[7]),
        .O(info_sf7[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__0
       (.I0(self_sf7[6]),
        .O(info_sf7[6]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__1
       (.I0(self_sf7[5]),
        .O(info_sf7[5]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__2
       (.I0(self_sf7[4]),
        .O(info_sf7[4]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__3
       (.I0(self_sf7[3]),
        .O(info_sf7[3]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__4
       (.I0(self_sf7[2]),
        .O(info_sf7[2]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__5
       (.I0(self_sf7[1]),
        .O(info_sf7[1]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__6
       (.I0(self_sf7[0]),
        .O(info_sf7[0]));
endmodule

(* ORIG_REF_NAME = "muxer" *) (* box_type = "black_box" *) (* dont_touch = "true" *) 
module switch_elements_muxer__7
   (enable_i,
    info_o);
  input enable_i;
  output info_o;

  wire enable_i;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf7;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf8;
  (* RTL_KEEP = "true" *) (* S *) wire [7:0]info_sf9;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [1802:0]self_sf7;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf8;
  (* ALLOW_COMBINATORIAL_LOOPS *) (* RTL_KEEP = "true" *) (* S *) 
  (* equivalent_register_removal = "no" *) wire [3:0]self_sf9;

  assign info_o = info_sf7[1];
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[0]),
        .S(info_sf7[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1000].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1000]),
        .S(self_sf7[1000]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1001].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1001]),
        .S(self_sf7[1001]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1002].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1002]),
        .S(self_sf7[1002]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1003].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1003]),
        .S(self_sf7[1003]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1004].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1004]),
        .S(self_sf7[1004]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1005].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1005]),
        .S(self_sf7[1005]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1006].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1006]),
        .S(self_sf7[1006]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1007].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1007]),
        .S(self_sf7[1007]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1008].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1008]),
        .S(self_sf7[1008]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1009].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1009]),
        .S(self_sf7[1009]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[100]),
        .S(self_sf7[100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1010].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1010]),
        .S(self_sf7[1010]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1011].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1011]),
        .S(self_sf7[1011]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1012].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1012]),
        .S(self_sf7[1012]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1013].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1013]),
        .S(self_sf7[1013]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1014].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1014]),
        .S(self_sf7[1014]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1015].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1015]),
        .S(self_sf7[1015]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1016].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1016]),
        .S(self_sf7[1016]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1017].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1017]),
        .S(self_sf7[1017]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1018].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1018]),
        .S(self_sf7[1018]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1019].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1019]),
        .S(self_sf7[1019]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[101]),
        .S(self_sf7[101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1020].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1020]),
        .S(self_sf7[1020]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1021].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1021]),
        .S(self_sf7[1021]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1022].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1022]),
        .S(self_sf7[1022]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1023].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1023]),
        .S(self_sf7[1023]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1024].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1024]),
        .S(self_sf7[1024]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1025].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1025]),
        .S(self_sf7[1025]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1026].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1026]),
        .S(self_sf7[1026]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1027].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1027]),
        .S(self_sf7[1027]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1028].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1028]),
        .S(self_sf7[1028]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1029].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1029]),
        .S(self_sf7[1029]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[102]),
        .S(self_sf7[102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1030].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1030]),
        .S(self_sf7[1030]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1031].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1031]),
        .S(self_sf7[1031]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1032].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1032]),
        .S(self_sf7[1032]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1033].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1033]),
        .S(self_sf7[1033]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1034].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1034]),
        .S(self_sf7[1034]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1035].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1035]),
        .S(self_sf7[1035]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1036].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1036]),
        .S(self_sf7[1036]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1037].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1037]),
        .S(self_sf7[1037]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1038].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1038]),
        .S(self_sf7[1038]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1039].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1039]),
        .S(self_sf7[1039]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[103]),
        .S(self_sf7[103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1040].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1040]),
        .S(self_sf7[1040]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1041].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1041]),
        .S(self_sf7[1041]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1042].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1042]),
        .S(self_sf7[1042]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1043].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1043]),
        .S(self_sf7[1043]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1044].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1044]),
        .S(self_sf7[1044]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1045].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1045]),
        .S(self_sf7[1045]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1046].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1046]),
        .S(self_sf7[1046]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1047].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1047]),
        .S(self_sf7[1047]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1048].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1048]),
        .S(self_sf7[1048]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1049].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1049]),
        .S(self_sf7[1049]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[104]),
        .S(self_sf7[104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1050].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1050]),
        .S(self_sf7[1050]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1051].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1051]),
        .S(self_sf7[1051]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1052].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1052]),
        .S(self_sf7[1052]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1053].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1053]),
        .S(self_sf7[1053]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1054].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1054]),
        .S(self_sf7[1054]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1055].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1055]),
        .S(self_sf7[1055]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1056].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1056]),
        .S(self_sf7[1056]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1057].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1057]),
        .S(self_sf7[1057]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1058].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1058]),
        .S(self_sf7[1058]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1059].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1059]),
        .S(self_sf7[1059]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[105]),
        .S(self_sf7[105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1060].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1060]),
        .S(self_sf7[1060]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1061].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1061]),
        .S(self_sf7[1061]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1062].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1062]),
        .S(self_sf7[1062]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1063].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1063]),
        .S(self_sf7[1063]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1064].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1064]),
        .S(self_sf7[1064]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1065].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1065]),
        .S(self_sf7[1065]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1066].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1066]),
        .S(self_sf7[1066]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1067].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1067]),
        .S(self_sf7[1067]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1068].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1068]),
        .S(self_sf7[1068]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1069].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1069]),
        .S(self_sf7[1069]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[106]),
        .S(self_sf7[106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1070].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1070]),
        .S(self_sf7[1070]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1071].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1071]),
        .S(self_sf7[1071]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1072].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1072]),
        .S(self_sf7[1072]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1073].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1073]),
        .S(self_sf7[1073]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1074].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1074]),
        .S(self_sf7[1074]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1075].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1075]),
        .S(self_sf7[1075]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1076].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1076]),
        .S(self_sf7[1076]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1077].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1077]),
        .S(self_sf7[1077]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1078].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1078]),
        .S(self_sf7[1078]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1079].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1079]),
        .S(self_sf7[1079]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[107]),
        .S(self_sf7[107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1080].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1080]),
        .S(self_sf7[1080]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1081].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1081]),
        .S(self_sf7[1081]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1082].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1082]),
        .S(self_sf7[1082]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1083].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1083]),
        .S(self_sf7[1083]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1084].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1084]),
        .S(self_sf7[1084]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1085].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1085]),
        .S(self_sf7[1085]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1086].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1086]),
        .S(self_sf7[1086]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1087].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1087]),
        .S(self_sf7[1087]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1088].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1088]),
        .S(self_sf7[1088]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1089].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1089]),
        .S(self_sf7[1089]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[108]),
        .S(self_sf7[108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1090].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1090]),
        .S(self_sf7[1090]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1091].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1091]),
        .S(self_sf7[1091]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1092].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1092]),
        .S(self_sf7[1092]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1093].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1093]),
        .S(self_sf7[1093]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1094].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1094]),
        .S(self_sf7[1094]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1095].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1095]),
        .S(self_sf7[1095]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1096].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1096]),
        .S(self_sf7[1096]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1097].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1097]),
        .S(self_sf7[1097]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1098].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1098]),
        .S(self_sf7[1098]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1099].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1099]),
        .S(self_sf7[1099]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[109]),
        .S(self_sf7[109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[10].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[10]),
        .S(self_sf7[10]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1100].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1100]),
        .S(self_sf7[1100]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1101].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1101]),
        .S(self_sf7[1101]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1102].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1102]),
        .S(self_sf7[1102]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1103].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1103]),
        .S(self_sf7[1103]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1104].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1104]),
        .S(self_sf7[1104]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1105].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1105]),
        .S(self_sf7[1105]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1106].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1106]),
        .S(self_sf7[1106]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1107].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1107]),
        .S(self_sf7[1107]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1108].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1108]),
        .S(self_sf7[1108]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1109].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1109]),
        .S(self_sf7[1109]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[110]),
        .S(self_sf7[110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1110].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1110]),
        .S(self_sf7[1110]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1111]),
        .S(self_sf7[1111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1112]),
        .S(self_sf7[1112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1113]),
        .S(self_sf7[1113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1114]),
        .S(self_sf7[1114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1115]),
        .S(self_sf7[1115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1116]),
        .S(self_sf7[1116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1117]),
        .S(self_sf7[1117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1118]),
        .S(self_sf7[1118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1119]),
        .S(self_sf7[1119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[111].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[111]),
        .S(self_sf7[111]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1120]),
        .S(self_sf7[1120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1121]),
        .S(self_sf7[1121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1122]),
        .S(self_sf7[1122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1123]),
        .S(self_sf7[1123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1124]),
        .S(self_sf7[1124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1125]),
        .S(self_sf7[1125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1126]),
        .S(self_sf7[1126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1127]),
        .S(self_sf7[1127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1128]),
        .S(self_sf7[1128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1129]),
        .S(self_sf7[1129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[112].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[112]),
        .S(self_sf7[112]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1130]),
        .S(self_sf7[1130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1131]),
        .S(self_sf7[1131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1132]),
        .S(self_sf7[1132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1133]),
        .S(self_sf7[1133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1134]),
        .S(self_sf7[1134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1135]),
        .S(self_sf7[1135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1136]),
        .S(self_sf7[1136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1137]),
        .S(self_sf7[1137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1138]),
        .S(self_sf7[1138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1139]),
        .S(self_sf7[1139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[113].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[113]),
        .S(self_sf7[113]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1140]),
        .S(self_sf7[1140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1141]),
        .S(self_sf7[1141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1142]),
        .S(self_sf7[1142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1143]),
        .S(self_sf7[1143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1144]),
        .S(self_sf7[1144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1145]),
        .S(self_sf7[1145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1146]),
        .S(self_sf7[1146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1147]),
        .S(self_sf7[1147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1148]),
        .S(self_sf7[1148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1149]),
        .S(self_sf7[1149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[114].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[114]),
        .S(self_sf7[114]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1150]),
        .S(self_sf7[1150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1151]),
        .S(self_sf7[1151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1152]),
        .S(self_sf7[1152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1153]),
        .S(self_sf7[1153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1154]),
        .S(self_sf7[1154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1155]),
        .S(self_sf7[1155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1156]),
        .S(self_sf7[1156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1157]),
        .S(self_sf7[1157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1158]),
        .S(self_sf7[1158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1159]),
        .S(self_sf7[1159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[115].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[115]),
        .S(self_sf7[115]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1160]),
        .S(self_sf7[1160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1161]),
        .S(self_sf7[1161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1162]),
        .S(self_sf7[1162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1163]),
        .S(self_sf7[1163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1164]),
        .S(self_sf7[1164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1165]),
        .S(self_sf7[1165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1166]),
        .S(self_sf7[1166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1167]),
        .S(self_sf7[1167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1168]),
        .S(self_sf7[1168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1169]),
        .S(self_sf7[1169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[116].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[116]),
        .S(self_sf7[116]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1170]),
        .S(self_sf7[1170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1171]),
        .S(self_sf7[1171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1172]),
        .S(self_sf7[1172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1173]),
        .S(self_sf7[1173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1174]),
        .S(self_sf7[1174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1175]),
        .S(self_sf7[1175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1176]),
        .S(self_sf7[1176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1177]),
        .S(self_sf7[1177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1178]),
        .S(self_sf7[1178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1179]),
        .S(self_sf7[1179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[117].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[117]),
        .S(self_sf7[117]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1180]),
        .S(self_sf7[1180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1181]),
        .S(self_sf7[1181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1182]),
        .S(self_sf7[1182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1183]),
        .S(self_sf7[1183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1184]),
        .S(self_sf7[1184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1185]),
        .S(self_sf7[1185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1186]),
        .S(self_sf7[1186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1187]),
        .S(self_sf7[1187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1188]),
        .S(self_sf7[1188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1189]),
        .S(self_sf7[1189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[118].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[118]),
        .S(self_sf7[118]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1190]),
        .S(self_sf7[1190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1191]),
        .S(self_sf7[1191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1192]),
        .S(self_sf7[1192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1193]),
        .S(self_sf7[1193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1194]),
        .S(self_sf7[1194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1195]),
        .S(self_sf7[1195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1196]),
        .S(self_sf7[1196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1197]),
        .S(self_sf7[1197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1198]),
        .S(self_sf7[1198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1199]),
        .S(self_sf7[1199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[119].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[119]),
        .S(self_sf7[119]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[11].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[11]),
        .S(self_sf7[11]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1200]),
        .S(self_sf7[1200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1201]),
        .S(self_sf7[1201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1202]),
        .S(self_sf7[1202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1203]),
        .S(self_sf7[1203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1204]),
        .S(self_sf7[1204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1205]),
        .S(self_sf7[1205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1206]),
        .S(self_sf7[1206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1207]),
        .S(self_sf7[1207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1208]),
        .S(self_sf7[1208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1209]),
        .S(self_sf7[1209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[120].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[120]),
        .S(self_sf7[120]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1210]),
        .S(self_sf7[1210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1211]),
        .S(self_sf7[1211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1212]),
        .S(self_sf7[1212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1213]),
        .S(self_sf7[1213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1214]),
        .S(self_sf7[1214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1215]),
        .S(self_sf7[1215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1216]),
        .S(self_sf7[1216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1217]),
        .S(self_sf7[1217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1218]),
        .S(self_sf7[1218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1219]),
        .S(self_sf7[1219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[121].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[121]),
        .S(self_sf7[121]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1220]),
        .S(self_sf7[1220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1221]),
        .S(self_sf7[1221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1222]),
        .S(self_sf7[1222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1223]),
        .S(self_sf7[1223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1224]),
        .S(self_sf7[1224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1225]),
        .S(self_sf7[1225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1226]),
        .S(self_sf7[1226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1227]),
        .S(self_sf7[1227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1228]),
        .S(self_sf7[1228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1229]),
        .S(self_sf7[1229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[122].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[122]),
        .S(self_sf7[122]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1230]),
        .S(self_sf7[1230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1231]),
        .S(self_sf7[1231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1232]),
        .S(self_sf7[1232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1233]),
        .S(self_sf7[1233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1234]),
        .S(self_sf7[1234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1235]),
        .S(self_sf7[1235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1236]),
        .S(self_sf7[1236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1237]),
        .S(self_sf7[1237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1238]),
        .S(self_sf7[1238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1239]),
        .S(self_sf7[1239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[123].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[123]),
        .S(self_sf7[123]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1240]),
        .S(self_sf7[1240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1241]),
        .S(self_sf7[1241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1242]),
        .S(self_sf7[1242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1243]),
        .S(self_sf7[1243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1244]),
        .S(self_sf7[1244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1245]),
        .S(self_sf7[1245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1246]),
        .S(self_sf7[1246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1247]),
        .S(self_sf7[1247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1248]),
        .S(self_sf7[1248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1249]),
        .S(self_sf7[1249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[124].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[124]),
        .S(self_sf7[124]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1250]),
        .S(self_sf7[1250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1251]),
        .S(self_sf7[1251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1252]),
        .S(self_sf7[1252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1253]),
        .S(self_sf7[1253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1254]),
        .S(self_sf7[1254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1255]),
        .S(self_sf7[1255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1256]),
        .S(self_sf7[1256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1257]),
        .S(self_sf7[1257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1258]),
        .S(self_sf7[1258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1259]),
        .S(self_sf7[1259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[125].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[125]),
        .S(self_sf7[125]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1260]),
        .S(self_sf7[1260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1261]),
        .S(self_sf7[1261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1262]),
        .S(self_sf7[1262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1263]),
        .S(self_sf7[1263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1264]),
        .S(self_sf7[1264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1265]),
        .S(self_sf7[1265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1266]),
        .S(self_sf7[1266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1267]),
        .S(self_sf7[1267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1268]),
        .S(self_sf7[1268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1269]),
        .S(self_sf7[1269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[126].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[126]),
        .S(self_sf7[126]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1270]),
        .S(self_sf7[1270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1271]),
        .S(self_sf7[1271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1272]),
        .S(self_sf7[1272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1273]),
        .S(self_sf7[1273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1274]),
        .S(self_sf7[1274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1275]),
        .S(self_sf7[1275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1276]),
        .S(self_sf7[1276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1277]),
        .S(self_sf7[1277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1278]),
        .S(self_sf7[1278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1279]),
        .S(self_sf7[1279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[127].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[127]),
        .S(self_sf7[127]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1280]),
        .S(self_sf7[1280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1281]),
        .S(self_sf7[1281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1282]),
        .S(self_sf7[1282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1283]),
        .S(self_sf7[1283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1284]),
        .S(self_sf7[1284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1285]),
        .S(self_sf7[1285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1286]),
        .S(self_sf7[1286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1287]),
        .S(self_sf7[1287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1288]),
        .S(self_sf7[1288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1289]),
        .S(self_sf7[1289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[128].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[128]),
        .S(self_sf7[128]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1290]),
        .S(self_sf7[1290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1291]),
        .S(self_sf7[1291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1292]),
        .S(self_sf7[1292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1293]),
        .S(self_sf7[1293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1294]),
        .S(self_sf7[1294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1295]),
        .S(self_sf7[1295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1296]),
        .S(self_sf7[1296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1297]),
        .S(self_sf7[1297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1298]),
        .S(self_sf7[1298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1299]),
        .S(self_sf7[1299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[129].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[129]),
        .S(self_sf7[129]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[12].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[12]),
        .S(self_sf7[12]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1300]),
        .S(self_sf7[1300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1301]),
        .S(self_sf7[1301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1302]),
        .S(self_sf7[1302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1303]),
        .S(self_sf7[1303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1304]),
        .S(self_sf7[1304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1305]),
        .S(self_sf7[1305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1306]),
        .S(self_sf7[1306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1307]),
        .S(self_sf7[1307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1308]),
        .S(self_sf7[1308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1309]),
        .S(self_sf7[1309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[130].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[130]),
        .S(self_sf7[130]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1310]),
        .S(self_sf7[1310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1311]),
        .S(self_sf7[1311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1312]),
        .S(self_sf7[1312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1313]),
        .S(self_sf7[1313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1314]),
        .S(self_sf7[1314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1315]),
        .S(self_sf7[1315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1316]),
        .S(self_sf7[1316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1317]),
        .S(self_sf7[1317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1318]),
        .S(self_sf7[1318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1319]),
        .S(self_sf7[1319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[131].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[131]),
        .S(self_sf7[131]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1320]),
        .S(self_sf7[1320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1321]),
        .S(self_sf7[1321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1322]),
        .S(self_sf7[1322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1323]),
        .S(self_sf7[1323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1324]),
        .S(self_sf7[1324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1325]),
        .S(self_sf7[1325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1326]),
        .S(self_sf7[1326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1327]),
        .S(self_sf7[1327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1328]),
        .S(self_sf7[1328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1329]),
        .S(self_sf7[1329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[132].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[132]),
        .S(self_sf7[132]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1330]),
        .S(self_sf7[1330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1331]),
        .S(self_sf7[1331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1332]),
        .S(self_sf7[1332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1333]),
        .S(self_sf7[1333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1334]),
        .S(self_sf7[1334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1335]),
        .S(self_sf7[1335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1336]),
        .S(self_sf7[1336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1337]),
        .S(self_sf7[1337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1338]),
        .S(self_sf7[1338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1339]),
        .S(self_sf7[1339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[133].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[133]),
        .S(self_sf7[133]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1340]),
        .S(self_sf7[1340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1341]),
        .S(self_sf7[1341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1342]),
        .S(self_sf7[1342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1343]),
        .S(self_sf7[1343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1344]),
        .S(self_sf7[1344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1345]),
        .S(self_sf7[1345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1346]),
        .S(self_sf7[1346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1347]),
        .S(self_sf7[1347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1348]),
        .S(self_sf7[1348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1349]),
        .S(self_sf7[1349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[134].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[134]),
        .S(self_sf7[134]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1350]),
        .S(self_sf7[1350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1351]),
        .S(self_sf7[1351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1352]),
        .S(self_sf7[1352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1353]),
        .S(self_sf7[1353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1354]),
        .S(self_sf7[1354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1355]),
        .S(self_sf7[1355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1356]),
        .S(self_sf7[1356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1357]),
        .S(self_sf7[1357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1358]),
        .S(self_sf7[1358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1359]),
        .S(self_sf7[1359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[135].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[135]),
        .S(self_sf7[135]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1360]),
        .S(self_sf7[1360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1361]),
        .S(self_sf7[1361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1362]),
        .S(self_sf7[1362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1363]),
        .S(self_sf7[1363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1364]),
        .S(self_sf7[1364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1365]),
        .S(self_sf7[1365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1366]),
        .S(self_sf7[1366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1367]),
        .S(self_sf7[1367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1368]),
        .S(self_sf7[1368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1369]),
        .S(self_sf7[1369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[136].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[136]),
        .S(self_sf7[136]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1370]),
        .S(self_sf7[1370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1371]),
        .S(self_sf7[1371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1372]),
        .S(self_sf7[1372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1373]),
        .S(self_sf7[1373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1374]),
        .S(self_sf7[1374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1375]),
        .S(self_sf7[1375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1376]),
        .S(self_sf7[1376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1377]),
        .S(self_sf7[1377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1378]),
        .S(self_sf7[1378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1379]),
        .S(self_sf7[1379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[137].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[137]),
        .S(self_sf7[137]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1380]),
        .S(self_sf7[1380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1381]),
        .S(self_sf7[1381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1382]),
        .S(self_sf7[1382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1383]),
        .S(self_sf7[1383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1384]),
        .S(self_sf7[1384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1385]),
        .S(self_sf7[1385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1386]),
        .S(self_sf7[1386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1387]),
        .S(self_sf7[1387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1388]),
        .S(self_sf7[1388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1389]),
        .S(self_sf7[1389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[138].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[138]),
        .S(self_sf7[138]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1390]),
        .S(self_sf7[1390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1391]),
        .S(self_sf7[1391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1392]),
        .S(self_sf7[1392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1393]),
        .S(self_sf7[1393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1394]),
        .S(self_sf7[1394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1395]),
        .S(self_sf7[1395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1396]),
        .S(self_sf7[1396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1397]),
        .S(self_sf7[1397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1398]),
        .S(self_sf7[1398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1399]),
        .S(self_sf7[1399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[139].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[139]),
        .S(self_sf7[139]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[13].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[13]),
        .S(self_sf7[13]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1400]),
        .S(self_sf7[1400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1401]),
        .S(self_sf7[1401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1402]),
        .S(self_sf7[1402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1403]),
        .S(self_sf7[1403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1404]),
        .S(self_sf7[1404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1405]),
        .S(self_sf7[1405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1406]),
        .S(self_sf7[1406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1407]),
        .S(self_sf7[1407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1408]),
        .S(self_sf7[1408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1409]),
        .S(self_sf7[1409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[140].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[140]),
        .S(self_sf7[140]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1410]),
        .S(self_sf7[1410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1411]),
        .S(self_sf7[1411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1412]),
        .S(self_sf7[1412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1413]),
        .S(self_sf7[1413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1414]),
        .S(self_sf7[1414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1415]),
        .S(self_sf7[1415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1416]),
        .S(self_sf7[1416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1417]),
        .S(self_sf7[1417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1418]),
        .S(self_sf7[1418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1419]),
        .S(self_sf7[1419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[141].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[141]),
        .S(self_sf7[141]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1420]),
        .S(self_sf7[1420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1421]),
        .S(self_sf7[1421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1422]),
        .S(self_sf7[1422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1423]),
        .S(self_sf7[1423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1424]),
        .S(self_sf7[1424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1425]),
        .S(self_sf7[1425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1426]),
        .S(self_sf7[1426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1427]),
        .S(self_sf7[1427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1428]),
        .S(self_sf7[1428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1429]),
        .S(self_sf7[1429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[142].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[142]),
        .S(self_sf7[142]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1430]),
        .S(self_sf7[1430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1431]),
        .S(self_sf7[1431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1432]),
        .S(self_sf7[1432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1433]),
        .S(self_sf7[1433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1434]),
        .S(self_sf7[1434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1435]),
        .S(self_sf7[1435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1436]),
        .S(self_sf7[1436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1437]),
        .S(self_sf7[1437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1438]),
        .S(self_sf7[1438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1439]),
        .S(self_sf7[1439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[143].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[143]),
        .S(self_sf7[143]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1440]),
        .S(self_sf7[1440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1441]),
        .S(self_sf7[1441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1442]),
        .S(self_sf7[1442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1443]),
        .S(self_sf7[1443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1444]),
        .S(self_sf7[1444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1445]),
        .S(self_sf7[1445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1446]),
        .S(self_sf7[1446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1447]),
        .S(self_sf7[1447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1448]),
        .S(self_sf7[1448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1449]),
        .S(self_sf7[1449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[144].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[144]),
        .S(self_sf7[144]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1450]),
        .S(self_sf7[1450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1451]),
        .S(self_sf7[1451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1452]),
        .S(self_sf7[1452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1453]),
        .S(self_sf7[1453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1454]),
        .S(self_sf7[1454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1455]),
        .S(self_sf7[1455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1456]),
        .S(self_sf7[1456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1457]),
        .S(self_sf7[1457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1458]),
        .S(self_sf7[1458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1459]),
        .S(self_sf7[1459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[145].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[145]),
        .S(self_sf7[145]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1460]),
        .S(self_sf7[1460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1461]),
        .S(self_sf7[1461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1462]),
        .S(self_sf7[1462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1463]),
        .S(self_sf7[1463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1464]),
        .S(self_sf7[1464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1465]),
        .S(self_sf7[1465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1466]),
        .S(self_sf7[1466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1467]),
        .S(self_sf7[1467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1468]),
        .S(self_sf7[1468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1469]),
        .S(self_sf7[1469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[146].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[146]),
        .S(self_sf7[146]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1470]),
        .S(self_sf7[1470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1471]),
        .S(self_sf7[1471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1472]),
        .S(self_sf7[1472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1473]),
        .S(self_sf7[1473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1474]),
        .S(self_sf7[1474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1475]),
        .S(self_sf7[1475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1476]),
        .S(self_sf7[1476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1477]),
        .S(self_sf7[1477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1478]),
        .S(self_sf7[1478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1479]),
        .S(self_sf7[1479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[147].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[147]),
        .S(self_sf7[147]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1480]),
        .S(self_sf7[1480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1481]),
        .S(self_sf7[1481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1482]),
        .S(self_sf7[1482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1483]),
        .S(self_sf7[1483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1484]),
        .S(self_sf7[1484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1485]),
        .S(self_sf7[1485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1486]),
        .S(self_sf7[1486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1487]),
        .S(self_sf7[1487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1488]),
        .S(self_sf7[1488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1489]),
        .S(self_sf7[1489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[148].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[148]),
        .S(self_sf7[148]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1490]),
        .S(self_sf7[1490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1491]),
        .S(self_sf7[1491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1492]),
        .S(self_sf7[1492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1493]),
        .S(self_sf7[1493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1494]),
        .S(self_sf7[1494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1495]),
        .S(self_sf7[1495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1496]),
        .S(self_sf7[1496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1497]),
        .S(self_sf7[1497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1498]),
        .S(self_sf7[1498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1499]),
        .S(self_sf7[1499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[149].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[149]),
        .S(self_sf7[149]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[14].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[14]),
        .S(self_sf7[14]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1500]),
        .S(self_sf7[1500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1501]),
        .S(self_sf7[1501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1502]),
        .S(self_sf7[1502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1503]),
        .S(self_sf7[1503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1504]),
        .S(self_sf7[1504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1505]),
        .S(self_sf7[1505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1506]),
        .S(self_sf7[1506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1507]),
        .S(self_sf7[1507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1508]),
        .S(self_sf7[1508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1509]),
        .S(self_sf7[1509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[150].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[150]),
        .S(self_sf7[150]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1510]),
        .S(self_sf7[1510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1511]),
        .S(self_sf7[1511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1512]),
        .S(self_sf7[1512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1513]),
        .S(self_sf7[1513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1514]),
        .S(self_sf7[1514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1515]),
        .S(self_sf7[1515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1516]),
        .S(self_sf7[1516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1517]),
        .S(self_sf7[1517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1518]),
        .S(self_sf7[1518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1519]),
        .S(self_sf7[1519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[151].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[151]),
        .S(self_sf7[151]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1520]),
        .S(self_sf7[1520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1521]),
        .S(self_sf7[1521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1522]),
        .S(self_sf7[1522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1523]),
        .S(self_sf7[1523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1524]),
        .S(self_sf7[1524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1525]),
        .S(self_sf7[1525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1526]),
        .S(self_sf7[1526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1527]),
        .S(self_sf7[1527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1528]),
        .S(self_sf7[1528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1529]),
        .S(self_sf7[1529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[152].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[152]),
        .S(self_sf7[152]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1530]),
        .S(self_sf7[1530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1531]),
        .S(self_sf7[1531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1532]),
        .S(self_sf7[1532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1533]),
        .S(self_sf7[1533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1534]),
        .S(self_sf7[1534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1535]),
        .S(self_sf7[1535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1536]),
        .S(self_sf7[1536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1537]),
        .S(self_sf7[1537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1538]),
        .S(self_sf7[1538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1539]),
        .S(self_sf7[1539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[153].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[153]),
        .S(self_sf7[153]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1540]),
        .S(self_sf7[1540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1541]),
        .S(self_sf7[1541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1542]),
        .S(self_sf7[1542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1543]),
        .S(self_sf7[1543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1544]),
        .S(self_sf7[1544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1545]),
        .S(self_sf7[1545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1546]),
        .S(self_sf7[1546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1547]),
        .S(self_sf7[1547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1548]),
        .S(self_sf7[1548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1549]),
        .S(self_sf7[1549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[154].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[154]),
        .S(self_sf7[154]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1550]),
        .S(self_sf7[1550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1551]),
        .S(self_sf7[1551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1552]),
        .S(self_sf7[1552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1553]),
        .S(self_sf7[1553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1554]),
        .S(self_sf7[1554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1555]),
        .S(self_sf7[1555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1556]),
        .S(self_sf7[1556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1557]),
        .S(self_sf7[1557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1558]),
        .S(self_sf7[1558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1559]),
        .S(self_sf7[1559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[155].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[155]),
        .S(self_sf7[155]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1560]),
        .S(self_sf7[1560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1561]),
        .S(self_sf7[1561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1562]),
        .S(self_sf7[1562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1563]),
        .S(self_sf7[1563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1564]),
        .S(self_sf7[1564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1565]),
        .S(self_sf7[1565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1566]),
        .S(self_sf7[1566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1567]),
        .S(self_sf7[1567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1568]),
        .S(self_sf7[1568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1569]),
        .S(self_sf7[1569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[156].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[156]),
        .S(self_sf7[156]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1570]),
        .S(self_sf7[1570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1571]),
        .S(self_sf7[1571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1572]),
        .S(self_sf7[1572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1573]),
        .S(self_sf7[1573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1574]),
        .S(self_sf7[1574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1575]),
        .S(self_sf7[1575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1576]),
        .S(self_sf7[1576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1577]),
        .S(self_sf7[1577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1578]),
        .S(self_sf7[1578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1579]),
        .S(self_sf7[1579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[157].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[157]),
        .S(self_sf7[157]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1580]),
        .S(self_sf7[1580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1581]),
        .S(self_sf7[1581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1582]),
        .S(self_sf7[1582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1583]),
        .S(self_sf7[1583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1584]),
        .S(self_sf7[1584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1585]),
        .S(self_sf7[1585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1586]),
        .S(self_sf7[1586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1587]),
        .S(self_sf7[1587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1588]),
        .S(self_sf7[1588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1589]),
        .S(self_sf7[1589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[158].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[158]),
        .S(self_sf7[158]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1590]),
        .S(self_sf7[1590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1591]),
        .S(self_sf7[1591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1592]),
        .S(self_sf7[1592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1593]),
        .S(self_sf7[1593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1594]),
        .S(self_sf7[1594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1595]),
        .S(self_sf7[1595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1596]),
        .S(self_sf7[1596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1597]),
        .S(self_sf7[1597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1598]),
        .S(self_sf7[1598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1599]),
        .S(self_sf7[1599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[159].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[159]),
        .S(self_sf7[159]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[15].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[15]),
        .S(self_sf7[15]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1600]),
        .S(self_sf7[1600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1601]),
        .S(self_sf7[1601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1602]),
        .S(self_sf7[1602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1603]),
        .S(self_sf7[1603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1604]),
        .S(self_sf7[1604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1605]),
        .S(self_sf7[1605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1606]),
        .S(self_sf7[1606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1607]),
        .S(self_sf7[1607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1608]),
        .S(self_sf7[1608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1609]),
        .S(self_sf7[1609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[160].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[160]),
        .S(self_sf7[160]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1610]),
        .S(self_sf7[1610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1611]),
        .S(self_sf7[1611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1612]),
        .S(self_sf7[1612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1613]),
        .S(self_sf7[1613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1614]),
        .S(self_sf7[1614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1615]),
        .S(self_sf7[1615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1616]),
        .S(self_sf7[1616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1617]),
        .S(self_sf7[1617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1618]),
        .S(self_sf7[1618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1619]),
        .S(self_sf7[1619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[161].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[161]),
        .S(self_sf7[161]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1620]),
        .S(self_sf7[1620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1621]),
        .S(self_sf7[1621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1622]),
        .S(self_sf7[1622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1623]),
        .S(self_sf7[1623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1624]),
        .S(self_sf7[1624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1625]),
        .S(self_sf7[1625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1626]),
        .S(self_sf7[1626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1627]),
        .S(self_sf7[1627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1628]),
        .S(self_sf7[1628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1629]),
        .S(self_sf7[1629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[162].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[162]),
        .S(self_sf7[162]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1630]),
        .S(self_sf7[1630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1631]),
        .S(self_sf7[1631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1632]),
        .S(self_sf7[1632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1633]),
        .S(self_sf7[1633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1634]),
        .S(self_sf7[1634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1635]),
        .S(self_sf7[1635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1636]),
        .S(self_sf7[1636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1637]),
        .S(self_sf7[1637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1638]),
        .S(self_sf7[1638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1639]),
        .S(self_sf7[1639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[163].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[163]),
        .S(self_sf7[163]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1640]),
        .S(self_sf7[1640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1641]),
        .S(self_sf7[1641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1642]),
        .S(self_sf7[1642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1643]),
        .S(self_sf7[1643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1644]),
        .S(self_sf7[1644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1645]),
        .S(self_sf7[1645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1646]),
        .S(self_sf7[1646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1647]),
        .S(self_sf7[1647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1648]),
        .S(self_sf7[1648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1649]),
        .S(self_sf7[1649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[164].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[164]),
        .S(self_sf7[164]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1650]),
        .S(self_sf7[1650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1651]),
        .S(self_sf7[1651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1652]),
        .S(self_sf7[1652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1653]),
        .S(self_sf7[1653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1654]),
        .S(self_sf7[1654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1655]),
        .S(self_sf7[1655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1656]),
        .S(self_sf7[1656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1657]),
        .S(self_sf7[1657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1658]),
        .S(self_sf7[1658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1659]),
        .S(self_sf7[1659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[165].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[165]),
        .S(self_sf7[165]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1660]),
        .S(self_sf7[1660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1661]),
        .S(self_sf7[1661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1662]),
        .S(self_sf7[1662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1663]),
        .S(self_sf7[1663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1664]),
        .S(self_sf7[1664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1665]),
        .S(self_sf7[1665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1666]),
        .S(self_sf7[1666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1667]),
        .S(self_sf7[1667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1668]),
        .S(self_sf7[1668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1669]),
        .S(self_sf7[1669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[166].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[166]),
        .S(self_sf7[166]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1670]),
        .S(self_sf7[1670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1671]),
        .S(self_sf7[1671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1672]),
        .S(self_sf7[1672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1673]),
        .S(self_sf7[1673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1674]),
        .S(self_sf7[1674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1675]),
        .S(self_sf7[1675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1676]),
        .S(self_sf7[1676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1677]),
        .S(self_sf7[1677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1678]),
        .S(self_sf7[1678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1679]),
        .S(self_sf7[1679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[167].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[167]),
        .S(self_sf7[167]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1680]),
        .S(self_sf7[1680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1681]),
        .S(self_sf7[1681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1682]),
        .S(self_sf7[1682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1683]),
        .S(self_sf7[1683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1684]),
        .S(self_sf7[1684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1685]),
        .S(self_sf7[1685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1686]),
        .S(self_sf7[1686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1687]),
        .S(self_sf7[1687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1688]),
        .S(self_sf7[1688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1689]),
        .S(self_sf7[1689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[168].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[168]),
        .S(self_sf7[168]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1690]),
        .S(self_sf7[1690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1691]),
        .S(self_sf7[1691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1692]),
        .S(self_sf7[1692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1693]),
        .S(self_sf7[1693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1694]),
        .S(self_sf7[1694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1695]),
        .S(self_sf7[1695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1696]),
        .S(self_sf7[1696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1697]),
        .S(self_sf7[1697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1698]),
        .S(self_sf7[1698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1699]),
        .S(self_sf7[1699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[169].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[169]),
        .S(self_sf7[169]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[16].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[16]),
        .S(self_sf7[16]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1700]),
        .S(self_sf7[1700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1701]),
        .S(self_sf7[1701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1702]),
        .S(self_sf7[1702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1703]),
        .S(self_sf7[1703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1704]),
        .S(self_sf7[1704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1705]),
        .S(self_sf7[1705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1706]),
        .S(self_sf7[1706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1707]),
        .S(self_sf7[1707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1708]),
        .S(self_sf7[1708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1709]),
        .S(self_sf7[1709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[170].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[170]),
        .S(self_sf7[170]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1710]),
        .S(self_sf7[1710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1711]),
        .S(self_sf7[1711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1712]),
        .S(self_sf7[1712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1713]),
        .S(self_sf7[1713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1714]),
        .S(self_sf7[1714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1715]),
        .S(self_sf7[1715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1716]),
        .S(self_sf7[1716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1717]),
        .S(self_sf7[1717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1718]),
        .S(self_sf7[1718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1719]),
        .S(self_sf7[1719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[171].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[171]),
        .S(self_sf7[171]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1720]),
        .S(self_sf7[1720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1721]),
        .S(self_sf7[1721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1722]),
        .S(self_sf7[1722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1723]),
        .S(self_sf7[1723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1724]),
        .S(self_sf7[1724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1725]),
        .S(self_sf7[1725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1726]),
        .S(self_sf7[1726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1727]),
        .S(self_sf7[1727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1728]),
        .S(self_sf7[1728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1729]),
        .S(self_sf7[1729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[172].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[172]),
        .S(self_sf7[172]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1730]),
        .S(self_sf7[1730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1731]),
        .S(self_sf7[1731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1732]),
        .S(self_sf7[1732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1733]),
        .S(self_sf7[1733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1734]),
        .S(self_sf7[1734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1735]),
        .S(self_sf7[1735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1736]),
        .S(self_sf7[1736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1737]),
        .S(self_sf7[1737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1738]),
        .S(self_sf7[1738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1739]),
        .S(self_sf7[1739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[173].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[173]),
        .S(self_sf7[173]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1740]),
        .S(self_sf7[1740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1741]),
        .S(self_sf7[1741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1742]),
        .S(self_sf7[1742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1743]),
        .S(self_sf7[1743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1744]),
        .S(self_sf7[1744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1745]),
        .S(self_sf7[1745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1746]),
        .S(self_sf7[1746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1747]),
        .S(self_sf7[1747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1748]),
        .S(self_sf7[1748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1749]),
        .S(self_sf7[1749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[174].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[174]),
        .S(self_sf7[174]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1750]),
        .S(self_sf7[1750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1751]),
        .S(self_sf7[1751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1752]),
        .S(self_sf7[1752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1753]),
        .S(self_sf7[1753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1754]),
        .S(self_sf7[1754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1755]),
        .S(self_sf7[1755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1756]),
        .S(self_sf7[1756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1757]),
        .S(self_sf7[1757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1758]),
        .S(self_sf7[1758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1759]),
        .S(self_sf7[1759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[175].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[175]),
        .S(self_sf7[175]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1760]),
        .S(self_sf7[1760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1761]),
        .S(self_sf7[1761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1762]),
        .S(self_sf7[1762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1763]),
        .S(self_sf7[1763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1764]),
        .S(self_sf7[1764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1765]),
        .S(self_sf7[1765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1766]),
        .S(self_sf7[1766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1767]),
        .S(self_sf7[1767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1768]),
        .S(self_sf7[1768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1769]),
        .S(self_sf7[1769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[176].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[176]),
        .S(self_sf7[176]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1770]),
        .S(self_sf7[1770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1771]),
        .S(self_sf7[1771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1772]),
        .S(self_sf7[1772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1773]),
        .S(self_sf7[1773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1774]),
        .S(self_sf7[1774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1775]),
        .S(self_sf7[1775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1776]),
        .S(self_sf7[1776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1777]),
        .S(self_sf7[1777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1778]),
        .S(self_sf7[1778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1779]),
        .S(self_sf7[1779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[177].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[177]),
        .S(self_sf7[177]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1780]),
        .S(self_sf7[1780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1781]),
        .S(self_sf7[1781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1782]),
        .S(self_sf7[1782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1783]),
        .S(self_sf7[1783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1784]),
        .S(self_sf7[1784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1785]),
        .S(self_sf7[1785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1786]),
        .S(self_sf7[1786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1787]),
        .S(self_sf7[1787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1788]),
        .S(self_sf7[1788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1789]),
        .S(self_sf7[1789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[178].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[178]),
        .S(self_sf7[178]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1790]),
        .S(self_sf7[1790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1791]),
        .S(self_sf7[1791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1792]),
        .S(self_sf7[1792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1793]),
        .S(self_sf7[1793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1794]),
        .S(self_sf7[1794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1795]),
        .S(self_sf7[1795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1796]),
        .S(self_sf7[1796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1797]),
        .S(self_sf7[1797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1798]),
        .S(self_sf7[1798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1799]),
        .S(self_sf7[1799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[179].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[179]),
        .S(self_sf7[179]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[17].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[17]),
        .S(self_sf7[17]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[180].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[180]),
        .S(self_sf7[180]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[181].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[181]),
        .S(self_sf7[181]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[182].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[182]),
        .S(self_sf7[182]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[183].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[183]),
        .S(self_sf7[183]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[184].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[184]),
        .S(self_sf7[184]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[185].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[185]),
        .S(self_sf7[185]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[186].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[186]),
        .S(self_sf7[186]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[187].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[187]),
        .S(self_sf7[187]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[188].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[188]),
        .S(self_sf7[188]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[189].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[189]),
        .S(self_sf7[189]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[18].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[18]),
        .S(self_sf7[18]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[190].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[190]),
        .S(self_sf7[190]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[191].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[191]),
        .S(self_sf7[191]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[192].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[192]),
        .S(self_sf7[192]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[193].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[193]),
        .S(self_sf7[193]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[194].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[194]),
        .S(self_sf7[194]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[195].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[195]),
        .S(self_sf7[195]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[196].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[196]),
        .S(self_sf7[196]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[197].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[197]),
        .S(self_sf7[197]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[198].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[198]),
        .S(self_sf7[198]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[199].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[199]),
        .S(self_sf7[199]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[19].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[19]),
        .S(self_sf7[19]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[1].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[1]),
        .S(info_sf7[1]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[200].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[200]),
        .S(self_sf7[200]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[201].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[201]),
        .S(self_sf7[201]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[202].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[202]),
        .S(self_sf7[202]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[203].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[203]),
        .S(self_sf7[203]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[204].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[204]),
        .S(self_sf7[204]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[205].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[205]),
        .S(self_sf7[205]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[206].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[206]),
        .S(self_sf7[206]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[207].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[207]),
        .S(self_sf7[207]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[208].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[208]),
        .S(self_sf7[208]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[209].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[209]),
        .S(self_sf7[209]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[20].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[20]),
        .S(self_sf7[20]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[210].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[210]),
        .S(self_sf7[210]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[211].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[211]),
        .S(self_sf7[211]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[212].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[212]),
        .S(self_sf7[212]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[213].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[213]),
        .S(self_sf7[213]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[214].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[214]),
        .S(self_sf7[214]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[215].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[215]),
        .S(self_sf7[215]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[216].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[216]),
        .S(self_sf7[216]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[217].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[217]),
        .S(self_sf7[217]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[218].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[218]),
        .S(self_sf7[218]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[219].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[219]),
        .S(self_sf7[219]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[21].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[21]),
        .S(self_sf7[21]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[220].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[220]),
        .S(self_sf7[220]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[221].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[221]),
        .S(self_sf7[221]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[222].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[222]),
        .S(self_sf7[222]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[223].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[223]),
        .S(self_sf7[223]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[224].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[224]),
        .S(self_sf7[224]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[225].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[225]),
        .S(self_sf7[225]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[226].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[226]),
        .S(self_sf7[226]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[227].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[227]),
        .S(self_sf7[227]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[228].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[228]),
        .S(self_sf7[228]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[229].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[229]),
        .S(self_sf7[229]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[22].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[22]),
        .S(self_sf7[22]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[230].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[230]),
        .S(self_sf7[230]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[231].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[231]),
        .S(self_sf7[231]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[232].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[232]),
        .S(self_sf7[232]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[233].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[233]),
        .S(self_sf7[233]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[234].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[234]),
        .S(self_sf7[234]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[235].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[235]),
        .S(self_sf7[235]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[236].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[236]),
        .S(self_sf7[236]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[237].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[237]),
        .S(self_sf7[237]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[238].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[238]),
        .S(self_sf7[238]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[239].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[239]),
        .S(self_sf7[239]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[23].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[23]),
        .S(self_sf7[23]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[240].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[240]),
        .S(self_sf7[240]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[241].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[241]),
        .S(self_sf7[241]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[242].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[242]),
        .S(self_sf7[242]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[243].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[243]),
        .S(self_sf7[243]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[244].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[244]),
        .S(self_sf7[244]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[245].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[245]),
        .S(self_sf7[245]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[246].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[246]),
        .S(self_sf7[246]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[247].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[247]),
        .S(self_sf7[247]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[248].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[248]),
        .S(self_sf7[248]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[249].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[249]),
        .S(self_sf7[249]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[24].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[24]),
        .S(self_sf7[24]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[250].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[250]),
        .S(self_sf7[250]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[251].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[251]),
        .S(self_sf7[251]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[252].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[252]),
        .S(self_sf7[252]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[253].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[253]),
        .S(self_sf7[253]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[254].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[254]),
        .S(self_sf7[254]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[255].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[255]),
        .S(self_sf7[255]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[256].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[256]),
        .S(self_sf7[256]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[257].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[257]),
        .S(self_sf7[257]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[258].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[258]),
        .S(self_sf7[258]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[259].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[259]),
        .S(self_sf7[259]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[25].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[25]),
        .S(self_sf7[25]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[260].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[260]),
        .S(self_sf7[260]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[261].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[261]),
        .S(self_sf7[261]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[262].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[262]),
        .S(self_sf7[262]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[263].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[263]),
        .S(self_sf7[263]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[264].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[264]),
        .S(self_sf7[264]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[265].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[265]),
        .S(self_sf7[265]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[266].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[266]),
        .S(self_sf7[266]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[267].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[267]),
        .S(self_sf7[267]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[268].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[268]),
        .S(self_sf7[268]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[269].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[269]),
        .S(self_sf7[269]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[26].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[26]),
        .S(self_sf7[26]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[270].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[270]),
        .S(self_sf7[270]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[271].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[271]),
        .S(self_sf7[271]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[272].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[272]),
        .S(self_sf7[272]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[273].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[273]),
        .S(self_sf7[273]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[274].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[274]),
        .S(self_sf7[274]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[275].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[275]),
        .S(self_sf7[275]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[276].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[276]),
        .S(self_sf7[276]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[277].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[277]),
        .S(self_sf7[277]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[278].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[278]),
        .S(self_sf7[278]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[279].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[279]),
        .S(self_sf7[279]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[27].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[27]),
        .S(self_sf7[27]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[280].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[280]),
        .S(self_sf7[280]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[281].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[281]),
        .S(self_sf7[281]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[282].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[282]),
        .S(self_sf7[282]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[283].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[283]),
        .S(self_sf7[283]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[284].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[284]),
        .S(self_sf7[284]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[285].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[285]),
        .S(self_sf7[285]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[286].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[286]),
        .S(self_sf7[286]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[287].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[287]),
        .S(self_sf7[287]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[288].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[288]),
        .S(self_sf7[288]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[289].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[289]),
        .S(self_sf7[289]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[28].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[28]),
        .S(self_sf7[28]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[290].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[290]),
        .S(self_sf7[290]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[291].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[291]),
        .S(self_sf7[291]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[292].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[292]),
        .S(self_sf7[292]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[293].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[293]),
        .S(self_sf7[293]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[294].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[294]),
        .S(self_sf7[294]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[295].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[295]),
        .S(self_sf7[295]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[296].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[296]),
        .S(self_sf7[296]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[297].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[297]),
        .S(self_sf7[297]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[298].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[298]),
        .S(self_sf7[298]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[299].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[299]),
        .S(self_sf7[299]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[29].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[29]),
        .S(self_sf7[29]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[2].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[2]),
        .S(info_sf7[2]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[300].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[300]),
        .S(self_sf7[300]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[301].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[301]),
        .S(self_sf7[301]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[302].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[302]),
        .S(self_sf7[302]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[303].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[303]),
        .S(self_sf7[303]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[304].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[304]),
        .S(self_sf7[304]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[305].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[305]),
        .S(self_sf7[305]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[306].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[306]),
        .S(self_sf7[306]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[307].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[307]),
        .S(self_sf7[307]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[308].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[308]),
        .S(self_sf7[308]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[309].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[309]),
        .S(self_sf7[309]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[30].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[30]),
        .S(self_sf7[30]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[310].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[310]),
        .S(self_sf7[310]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[311].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[311]),
        .S(self_sf7[311]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[312].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[312]),
        .S(self_sf7[312]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[313].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[313]),
        .S(self_sf7[313]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[314].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[314]),
        .S(self_sf7[314]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[315].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[315]),
        .S(self_sf7[315]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[316].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[316]),
        .S(self_sf7[316]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[317].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[317]),
        .S(self_sf7[317]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[318].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[318]),
        .S(self_sf7[318]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[319].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[319]),
        .S(self_sf7[319]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[31].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[31]),
        .S(self_sf7[31]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[320].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[320]),
        .S(self_sf7[320]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[321].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[321]),
        .S(self_sf7[321]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[322].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[322]),
        .S(self_sf7[322]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[323].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[323]),
        .S(self_sf7[323]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[324].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[324]),
        .S(self_sf7[324]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[325].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[325]),
        .S(self_sf7[325]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[326].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[326]),
        .S(self_sf7[326]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[327].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[327]),
        .S(self_sf7[327]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[328].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[328]),
        .S(self_sf7[328]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[329].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[329]),
        .S(self_sf7[329]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[32].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[32]),
        .S(self_sf7[32]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[330].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[330]),
        .S(self_sf7[330]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[331].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[331]),
        .S(self_sf7[331]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[332].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[332]),
        .S(self_sf7[332]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[333].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[333]),
        .S(self_sf7[333]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[334].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[334]),
        .S(self_sf7[334]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[335].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[335]),
        .S(self_sf7[335]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[336].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[336]),
        .S(self_sf7[336]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[337].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[337]),
        .S(self_sf7[337]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[338].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[338]),
        .S(self_sf7[338]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[339].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[339]),
        .S(self_sf7[339]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[33].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[33]),
        .S(self_sf7[33]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[340].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[340]),
        .S(self_sf7[340]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[341].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[341]),
        .S(self_sf7[341]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[342].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[342]),
        .S(self_sf7[342]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[343].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[343]),
        .S(self_sf7[343]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[344].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[344]),
        .S(self_sf7[344]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[345].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[345]),
        .S(self_sf7[345]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[346].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[346]),
        .S(self_sf7[346]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[347].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[347]),
        .S(self_sf7[347]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[348].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[348]),
        .S(self_sf7[348]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[349].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[349]),
        .S(self_sf7[349]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[34].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[34]),
        .S(self_sf7[34]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[350].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[350]),
        .S(self_sf7[350]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[351].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[351]),
        .S(self_sf7[351]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[352].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[352]),
        .S(self_sf7[352]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[353].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[353]),
        .S(self_sf7[353]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[354].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[354]),
        .S(self_sf7[354]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[355].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[355]),
        .S(self_sf7[355]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[356].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[356]),
        .S(self_sf7[356]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[357].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[357]),
        .S(self_sf7[357]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[358].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[358]),
        .S(self_sf7[358]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[359].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[359]),
        .S(self_sf7[359]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[35].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[35]),
        .S(self_sf7[35]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[360].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[360]),
        .S(self_sf7[360]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[361].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[361]),
        .S(self_sf7[361]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[362].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[362]),
        .S(self_sf7[362]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[363].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[363]),
        .S(self_sf7[363]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[364].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[364]),
        .S(self_sf7[364]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[365].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[365]),
        .S(self_sf7[365]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[366].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[366]),
        .S(self_sf7[366]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[367].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[367]),
        .S(self_sf7[367]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[368].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[368]),
        .S(self_sf7[368]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[369].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[369]),
        .S(self_sf7[369]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[36].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[36]),
        .S(self_sf7[36]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[370].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[370]),
        .S(self_sf7[370]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[371].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[371]),
        .S(self_sf7[371]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[372].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[372]),
        .S(self_sf7[372]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[373].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[373]),
        .S(self_sf7[373]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[374].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[374]),
        .S(self_sf7[374]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[375].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[375]),
        .S(self_sf7[375]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[376].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[376]),
        .S(self_sf7[376]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[377].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[377]),
        .S(self_sf7[377]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[378].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[378]),
        .S(self_sf7[378]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[379].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[379]),
        .S(self_sf7[379]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[37].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[37]),
        .S(self_sf7[37]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[380].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[380]),
        .S(self_sf7[380]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[381].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[381]),
        .S(self_sf7[381]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[382].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[382]),
        .S(self_sf7[382]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[383].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[383]),
        .S(self_sf7[383]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[384].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[384]),
        .S(self_sf7[384]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[385].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[385]),
        .S(self_sf7[385]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[386].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[386]),
        .S(self_sf7[386]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[387].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[387]),
        .S(self_sf7[387]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[388].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[388]),
        .S(self_sf7[388]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[389].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[389]),
        .S(self_sf7[389]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[38].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[38]),
        .S(self_sf7[38]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[390].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[390]),
        .S(self_sf7[390]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[391].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[391]),
        .S(self_sf7[391]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[392].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[392]),
        .S(self_sf7[392]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[393].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[393]),
        .S(self_sf7[393]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[394].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[394]),
        .S(self_sf7[394]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[395].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[395]),
        .S(self_sf7[395]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[396].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[396]),
        .S(self_sf7[396]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[397].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[397]),
        .S(self_sf7[397]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[398].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[398]),
        .S(self_sf7[398]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[399].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[399]),
        .S(self_sf7[399]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[39].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[39]),
        .S(self_sf7[39]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[3].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[3]),
        .S(info_sf7[3]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[400].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[400]),
        .S(self_sf7[400]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[401].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[401]),
        .S(self_sf7[401]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[402].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[402]),
        .S(self_sf7[402]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[403].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[403]),
        .S(self_sf7[403]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[404].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[404]),
        .S(self_sf7[404]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[405].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[405]),
        .S(self_sf7[405]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[406].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[406]),
        .S(self_sf7[406]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[407].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[407]),
        .S(self_sf7[407]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[408].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[408]),
        .S(self_sf7[408]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[409].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[409]),
        .S(self_sf7[409]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[40].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[40]),
        .S(self_sf7[40]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[410].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[410]),
        .S(self_sf7[410]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[411].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[411]),
        .S(self_sf7[411]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[412].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[412]),
        .S(self_sf7[412]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[413].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[413]),
        .S(self_sf7[413]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[414].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[414]),
        .S(self_sf7[414]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[415].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[415]),
        .S(self_sf7[415]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[416].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[416]),
        .S(self_sf7[416]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[417].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[417]),
        .S(self_sf7[417]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[418].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[418]),
        .S(self_sf7[418]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[419].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[419]),
        .S(self_sf7[419]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[41].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[41]),
        .S(self_sf7[41]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[420].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[420]),
        .S(self_sf7[420]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[421].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[421]),
        .S(self_sf7[421]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[422].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[422]),
        .S(self_sf7[422]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[423].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[423]),
        .S(self_sf7[423]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[424].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[424]),
        .S(self_sf7[424]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[425].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[425]),
        .S(self_sf7[425]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[426].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[426]),
        .S(self_sf7[426]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[427].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[427]),
        .S(self_sf7[427]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[428].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[428]),
        .S(self_sf7[428]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[429].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[429]),
        .S(self_sf7[429]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[42].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[42]),
        .S(self_sf7[42]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[430].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[430]),
        .S(self_sf7[430]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[431].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[431]),
        .S(self_sf7[431]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[432].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[432]),
        .S(self_sf7[432]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[433].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[433]),
        .S(self_sf7[433]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[434].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[434]),
        .S(self_sf7[434]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[435].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[435]),
        .S(self_sf7[435]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[436].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[436]),
        .S(self_sf7[436]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[437].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[437]),
        .S(self_sf7[437]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[438].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[438]),
        .S(self_sf7[438]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[439].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[439]),
        .S(self_sf7[439]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[43].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[43]),
        .S(self_sf7[43]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[440].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[440]),
        .S(self_sf7[440]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[441].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[441]),
        .S(self_sf7[441]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[442].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[442]),
        .S(self_sf7[442]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[443].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[443]),
        .S(self_sf7[443]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[444].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[444]),
        .S(self_sf7[444]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[445].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[445]),
        .S(self_sf7[445]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[446].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[446]),
        .S(self_sf7[446]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[447].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[447]),
        .S(self_sf7[447]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[448].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[448]),
        .S(self_sf7[448]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[449].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[449]),
        .S(self_sf7[449]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[44].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[44]),
        .S(self_sf7[44]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[450].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[450]),
        .S(self_sf7[450]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[451].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[451]),
        .S(self_sf7[451]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[452].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[452]),
        .S(self_sf7[452]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[453].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[453]),
        .S(self_sf7[453]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[454].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[454]),
        .S(self_sf7[454]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[455].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[455]),
        .S(self_sf7[455]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[456].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[456]),
        .S(self_sf7[456]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[457].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[457]),
        .S(self_sf7[457]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[458].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[458]),
        .S(self_sf7[458]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[459].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[459]),
        .S(self_sf7[459]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[45].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[45]),
        .S(self_sf7[45]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[460].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[460]),
        .S(self_sf7[460]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[461].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[461]),
        .S(self_sf7[461]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[462].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[462]),
        .S(self_sf7[462]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[463].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[463]),
        .S(self_sf7[463]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[464].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[464]),
        .S(self_sf7[464]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[465].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[465]),
        .S(self_sf7[465]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[466].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[466]),
        .S(self_sf7[466]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[467].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[467]),
        .S(self_sf7[467]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[468].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[468]),
        .S(self_sf7[468]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[469].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[469]),
        .S(self_sf7[469]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[46].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[46]),
        .S(self_sf7[46]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[470].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[470]),
        .S(self_sf7[470]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[471].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[471]),
        .S(self_sf7[471]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[472].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[472]),
        .S(self_sf7[472]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[473].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[473]),
        .S(self_sf7[473]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[474].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[474]),
        .S(self_sf7[474]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[475].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[475]),
        .S(self_sf7[475]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[476].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[476]),
        .S(self_sf7[476]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[477].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[477]),
        .S(self_sf7[477]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[478].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[478]),
        .S(self_sf7[478]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[479].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[479]),
        .S(self_sf7[479]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[47].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[47]),
        .S(self_sf7[47]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[480].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[480]),
        .S(self_sf7[480]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[481].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[481]),
        .S(self_sf7[481]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[482].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[482]),
        .S(self_sf7[482]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[483].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[483]),
        .S(self_sf7[483]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[484].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[484]),
        .S(self_sf7[484]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[485].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[485]),
        .S(self_sf7[485]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[486].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[486]),
        .S(self_sf7[486]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[487].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[487]),
        .S(self_sf7[487]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[488].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[488]),
        .S(self_sf7[488]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[489].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[489]),
        .S(self_sf7[489]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[48].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[48]),
        .S(self_sf7[48]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[490].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[490]),
        .S(self_sf7[490]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[491].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[491]),
        .S(self_sf7[491]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[492].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[492]),
        .S(self_sf7[492]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[493].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[493]),
        .S(self_sf7[493]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[494].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[494]),
        .S(self_sf7[494]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[495].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[495]),
        .S(self_sf7[495]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[496].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[496]),
        .S(self_sf7[496]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[497].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[497]),
        .S(self_sf7[497]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[498].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[498]),
        .S(self_sf7[498]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[499].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[499]),
        .S(self_sf7[499]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[49].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[49]),
        .S(self_sf7[49]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[4].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[4]),
        .S(info_sf7[4]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[500].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[500]),
        .S(self_sf7[500]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[501].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[501]),
        .S(self_sf7[501]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[502].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[502]),
        .S(self_sf7[502]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[503].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[503]),
        .S(self_sf7[503]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[504].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[504]),
        .S(self_sf7[504]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[505].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[505]),
        .S(self_sf7[505]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[506].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[506]),
        .S(self_sf7[506]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[507].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[507]),
        .S(self_sf7[507]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[508].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[508]),
        .S(self_sf7[508]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[509].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[509]),
        .S(self_sf7[509]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[50].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[50]),
        .S(self_sf7[50]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[510].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[510]),
        .S(self_sf7[510]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[511].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[511]),
        .S(self_sf7[511]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[512].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[512]),
        .S(self_sf7[512]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[513].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[513]),
        .S(self_sf7[513]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[514].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[514]),
        .S(self_sf7[514]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[515].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[515]),
        .S(self_sf7[515]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[516].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[516]),
        .S(self_sf7[516]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[517].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[517]),
        .S(self_sf7[517]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[518].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[518]),
        .S(self_sf7[518]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[519].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[519]),
        .S(self_sf7[519]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[51].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[51]),
        .S(self_sf7[51]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[520].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[520]),
        .S(self_sf7[520]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[521].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[521]),
        .S(self_sf7[521]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[522].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[522]),
        .S(self_sf7[522]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[523].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[523]),
        .S(self_sf7[523]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[524].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[524]),
        .S(self_sf7[524]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[525].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[525]),
        .S(self_sf7[525]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[526].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[526]),
        .S(self_sf7[526]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[527].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[527]),
        .S(self_sf7[527]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[528].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[528]),
        .S(self_sf7[528]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[529].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[529]),
        .S(self_sf7[529]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[52].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[52]),
        .S(self_sf7[52]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[530].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[530]),
        .S(self_sf7[530]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[531].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[531]),
        .S(self_sf7[531]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[532].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[532]),
        .S(self_sf7[532]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[533].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[533]),
        .S(self_sf7[533]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[534].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[534]),
        .S(self_sf7[534]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[535].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[535]),
        .S(self_sf7[535]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[536].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[536]),
        .S(self_sf7[536]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[537].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[537]),
        .S(self_sf7[537]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[538].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[538]),
        .S(self_sf7[538]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[539].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[539]),
        .S(self_sf7[539]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[53].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[53]),
        .S(self_sf7[53]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[540].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[540]),
        .S(self_sf7[540]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[541].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[541]),
        .S(self_sf7[541]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[542].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[542]),
        .S(self_sf7[542]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[543].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[543]),
        .S(self_sf7[543]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[544].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[544]),
        .S(self_sf7[544]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[545].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[545]),
        .S(self_sf7[545]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[546].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[546]),
        .S(self_sf7[546]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[547].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[547]),
        .S(self_sf7[547]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[548].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[548]),
        .S(self_sf7[548]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[549].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[549]),
        .S(self_sf7[549]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[54].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[54]),
        .S(self_sf7[54]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[550].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[550]),
        .S(self_sf7[550]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[551].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[551]),
        .S(self_sf7[551]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[552].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[552]),
        .S(self_sf7[552]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[553].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[553]),
        .S(self_sf7[553]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[554].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[554]),
        .S(self_sf7[554]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[555].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[555]),
        .S(self_sf7[555]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[556].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[556]),
        .S(self_sf7[556]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[557].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[557]),
        .S(self_sf7[557]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[558].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[558]),
        .S(self_sf7[558]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[559].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[559]),
        .S(self_sf7[559]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[55].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[55]),
        .S(self_sf7[55]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[560].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[560]),
        .S(self_sf7[560]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[561].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[561]),
        .S(self_sf7[561]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[562].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[562]),
        .S(self_sf7[562]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[563].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[563]),
        .S(self_sf7[563]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[564].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[564]),
        .S(self_sf7[564]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[565].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[565]),
        .S(self_sf7[565]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[566].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[566]),
        .S(self_sf7[566]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[567].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[567]),
        .S(self_sf7[567]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[568].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[568]),
        .S(self_sf7[568]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[569].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[569]),
        .S(self_sf7[569]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[56].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[56]),
        .S(self_sf7[56]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[570].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[570]),
        .S(self_sf7[570]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[571].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[571]),
        .S(self_sf7[571]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[572].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[572]),
        .S(self_sf7[572]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[573].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[573]),
        .S(self_sf7[573]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[574].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[574]),
        .S(self_sf7[574]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[575].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[575]),
        .S(self_sf7[575]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[576].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[576]),
        .S(self_sf7[576]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[577].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[577]),
        .S(self_sf7[577]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[578].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[578]),
        .S(self_sf7[578]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[579].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[579]),
        .S(self_sf7[579]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[57].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[57]),
        .S(self_sf7[57]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[580].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[580]),
        .S(self_sf7[580]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[581].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[581]),
        .S(self_sf7[581]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[582].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[582]),
        .S(self_sf7[582]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[583].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[583]),
        .S(self_sf7[583]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[584].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[584]),
        .S(self_sf7[584]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[585].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[585]),
        .S(self_sf7[585]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[586].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[586]),
        .S(self_sf7[586]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[587].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[587]),
        .S(self_sf7[587]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[588].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[588]),
        .S(self_sf7[588]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[589].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[589]),
        .S(self_sf7[589]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[58].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[58]),
        .S(self_sf7[58]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[590].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[590]),
        .S(self_sf7[590]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[591].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[591]),
        .S(self_sf7[591]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[592].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[592]),
        .S(self_sf7[592]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[593].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[593]),
        .S(self_sf7[593]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[594].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[594]),
        .S(self_sf7[594]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[595].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[595]),
        .S(self_sf7[595]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[596].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[596]),
        .S(self_sf7[596]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[597].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[597]),
        .S(self_sf7[597]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[598].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[598]),
        .S(self_sf7[598]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[599].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[599]),
        .S(self_sf7[599]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[59].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[59]),
        .S(self_sf7[59]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[5].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[5]),
        .S(info_sf7[5]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[600].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[600]),
        .S(self_sf7[600]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[601].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[601]),
        .S(self_sf7[601]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[602].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[602]),
        .S(self_sf7[602]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[603].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[603]),
        .S(self_sf7[603]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[604].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[604]),
        .S(self_sf7[604]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[605].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[605]),
        .S(self_sf7[605]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[606].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[606]),
        .S(self_sf7[606]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[607].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[607]),
        .S(self_sf7[607]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[608].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[608]),
        .S(self_sf7[608]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[609].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[609]),
        .S(self_sf7[609]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[60].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[60]),
        .S(self_sf7[60]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[610].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[610]),
        .S(self_sf7[610]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[611].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[611]),
        .S(self_sf7[611]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[612].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[612]),
        .S(self_sf7[612]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[613].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[613]),
        .S(self_sf7[613]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[614].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[614]),
        .S(self_sf7[614]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[615].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[615]),
        .S(self_sf7[615]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[616].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[616]),
        .S(self_sf7[616]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[617].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[617]),
        .S(self_sf7[617]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[618].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[618]),
        .S(self_sf7[618]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[619].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[619]),
        .S(self_sf7[619]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[61].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[61]),
        .S(self_sf7[61]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[620].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[620]),
        .S(self_sf7[620]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[621].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[621]),
        .S(self_sf7[621]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[622].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[622]),
        .S(self_sf7[622]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[623].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[623]),
        .S(self_sf7[623]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[624].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[624]),
        .S(self_sf7[624]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[625].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[625]),
        .S(self_sf7[625]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[626].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[626]),
        .S(self_sf7[626]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[627].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[627]),
        .S(self_sf7[627]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[628].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[628]),
        .S(self_sf7[628]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[629].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[629]),
        .S(self_sf7[629]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[62].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[62]),
        .S(self_sf7[62]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[630].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[630]),
        .S(self_sf7[630]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[631].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[631]),
        .S(self_sf7[631]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[632].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[632]),
        .S(self_sf7[632]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[633].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[633]),
        .S(self_sf7[633]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[634].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[634]),
        .S(self_sf7[634]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[635].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[635]),
        .S(self_sf7[635]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[636].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[636]),
        .S(self_sf7[636]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[637].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[637]),
        .S(self_sf7[637]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[638].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[638]),
        .S(self_sf7[638]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[639].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[639]),
        .S(self_sf7[639]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[63].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[63]),
        .S(self_sf7[63]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[640].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[640]),
        .S(self_sf7[640]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[641].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[641]),
        .S(self_sf7[641]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[642].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[642]),
        .S(self_sf7[642]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[643].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[643]),
        .S(self_sf7[643]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[644].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[644]),
        .S(self_sf7[644]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[645].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[645]),
        .S(self_sf7[645]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[646].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[646]),
        .S(self_sf7[646]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[647].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[647]),
        .S(self_sf7[647]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[648].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[648]),
        .S(self_sf7[648]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[649].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[649]),
        .S(self_sf7[649]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[64].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[64]),
        .S(self_sf7[64]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[650].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[650]),
        .S(self_sf7[650]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[651].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[651]),
        .S(self_sf7[651]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[652].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[652]),
        .S(self_sf7[652]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[653].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[653]),
        .S(self_sf7[653]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[654].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[654]),
        .S(self_sf7[654]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[655].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[655]),
        .S(self_sf7[655]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[656].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[656]),
        .S(self_sf7[656]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[657].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[657]),
        .S(self_sf7[657]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[658].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[658]),
        .S(self_sf7[658]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[659].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[659]),
        .S(self_sf7[659]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[65].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[65]),
        .S(self_sf7[65]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[660].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[660]),
        .S(self_sf7[660]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[661].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[661]),
        .S(self_sf7[661]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[662].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[662]),
        .S(self_sf7[662]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[663].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[663]),
        .S(self_sf7[663]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[664].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[664]),
        .S(self_sf7[664]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[665].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[665]),
        .S(self_sf7[665]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[666].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[666]),
        .S(self_sf7[666]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[667].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[667]),
        .S(self_sf7[667]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[668].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[668]),
        .S(self_sf7[668]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[669].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[669]),
        .S(self_sf7[669]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[66].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[66]),
        .S(self_sf7[66]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[670].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[670]),
        .S(self_sf7[670]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[671].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[671]),
        .S(self_sf7[671]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[672].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[672]),
        .S(self_sf7[672]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[673].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[673]),
        .S(self_sf7[673]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[674].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[674]),
        .S(self_sf7[674]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[675].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[675]),
        .S(self_sf7[675]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[676].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[676]),
        .S(self_sf7[676]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[677].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[677]),
        .S(self_sf7[677]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[678].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[678]),
        .S(self_sf7[678]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[679].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[679]),
        .S(self_sf7[679]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[67].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[67]),
        .S(self_sf7[67]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[680].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[680]),
        .S(self_sf7[680]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[681].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[681]),
        .S(self_sf7[681]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[682].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[682]),
        .S(self_sf7[682]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[683].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[683]),
        .S(self_sf7[683]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[684].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[684]),
        .S(self_sf7[684]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[685].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[685]),
        .S(self_sf7[685]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[686].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[686]),
        .S(self_sf7[686]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[687].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[687]),
        .S(self_sf7[687]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[688].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[688]),
        .S(self_sf7[688]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[689].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[689]),
        .S(self_sf7[689]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[68].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[68]),
        .S(self_sf7[68]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[690].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[690]),
        .S(self_sf7[690]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[691].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[691]),
        .S(self_sf7[691]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[692].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[692]),
        .S(self_sf7[692]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[693].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[693]),
        .S(self_sf7[693]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[694].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[694]),
        .S(self_sf7[694]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[695].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[695]),
        .S(self_sf7[695]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[696].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[696]),
        .S(self_sf7[696]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[697].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[697]),
        .S(self_sf7[697]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[698].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[698]),
        .S(self_sf7[698]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[699].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[699]),
        .S(self_sf7[699]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[69].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[69]),
        .S(self_sf7[69]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[6].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[6]),
        .S(info_sf7[6]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[700].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[700]),
        .S(self_sf7[700]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[701].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[701]),
        .S(self_sf7[701]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[702].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[702]),
        .S(self_sf7[702]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[703].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[703]),
        .S(self_sf7[703]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[704].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[704]),
        .S(self_sf7[704]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[705].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[705]),
        .S(self_sf7[705]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[706].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[706]),
        .S(self_sf7[706]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[707].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[707]),
        .S(self_sf7[707]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[708].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[708]),
        .S(self_sf7[708]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[709].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[709]),
        .S(self_sf7[709]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[70].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[70]),
        .S(self_sf7[70]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[710].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[710]),
        .S(self_sf7[710]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[711].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[711]),
        .S(self_sf7[711]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[712].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[712]),
        .S(self_sf7[712]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[713].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[713]),
        .S(self_sf7[713]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[714].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[714]),
        .S(self_sf7[714]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[715].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[715]),
        .S(self_sf7[715]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[716].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[716]),
        .S(self_sf7[716]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[717].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[717]),
        .S(self_sf7[717]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[718].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[718]),
        .S(self_sf7[718]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[719].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[719]),
        .S(self_sf7[719]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[71].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[71]),
        .S(self_sf7[71]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[720].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[720]),
        .S(self_sf7[720]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[721].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[721]),
        .S(self_sf7[721]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[722].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[722]),
        .S(self_sf7[722]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[723].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[723]),
        .S(self_sf7[723]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[724].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[724]),
        .S(self_sf7[724]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[725].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[725]),
        .S(self_sf7[725]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[726].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[726]),
        .S(self_sf7[726]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[727].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[727]),
        .S(self_sf7[727]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[728].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[728]),
        .S(self_sf7[728]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[729].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[729]),
        .S(self_sf7[729]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[72].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[72]),
        .S(self_sf7[72]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[730].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[730]),
        .S(self_sf7[730]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[731].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[731]),
        .S(self_sf7[731]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[732].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[732]),
        .S(self_sf7[732]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[733].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[733]),
        .S(self_sf7[733]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[734].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[734]),
        .S(self_sf7[734]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[735].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[735]),
        .S(self_sf7[735]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[736].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[736]),
        .S(self_sf7[736]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[737].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[737]),
        .S(self_sf7[737]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[738].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[738]),
        .S(self_sf7[738]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[739].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[739]),
        .S(self_sf7[739]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[73].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[73]),
        .S(self_sf7[73]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[740].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[740]),
        .S(self_sf7[740]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[741].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[741]),
        .S(self_sf7[741]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[742].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[742]),
        .S(self_sf7[742]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[743].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[743]),
        .S(self_sf7[743]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[744].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[744]),
        .S(self_sf7[744]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[745].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[745]),
        .S(self_sf7[745]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[746].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[746]),
        .S(self_sf7[746]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[747].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[747]),
        .S(self_sf7[747]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[748].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[748]),
        .S(self_sf7[748]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[749].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[749]),
        .S(self_sf7[749]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[74].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[74]),
        .S(self_sf7[74]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[750].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[750]),
        .S(self_sf7[750]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[751].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[751]),
        .S(self_sf7[751]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[752].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[752]),
        .S(self_sf7[752]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[753].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[753]),
        .S(self_sf7[753]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[754].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[754]),
        .S(self_sf7[754]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[755].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[755]),
        .S(self_sf7[755]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[756].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[756]),
        .S(self_sf7[756]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[757].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[757]),
        .S(self_sf7[757]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[758].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[758]),
        .S(self_sf7[758]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[759].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[759]),
        .S(self_sf7[759]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[75].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[75]),
        .S(self_sf7[75]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[760].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[760]),
        .S(self_sf7[760]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[761].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[761]),
        .S(self_sf7[761]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[762].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[762]),
        .S(self_sf7[762]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[763].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[763]),
        .S(self_sf7[763]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[764].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[764]),
        .S(self_sf7[764]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[765].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[765]),
        .S(self_sf7[765]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[766].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[766]),
        .S(self_sf7[766]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[767].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[767]),
        .S(self_sf7[767]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[768].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[768]),
        .S(self_sf7[768]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[769].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[769]),
        .S(self_sf7[769]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[76].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[76]),
        .S(self_sf7[76]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[770].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[770]),
        .S(self_sf7[770]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[771].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[771]),
        .S(self_sf7[771]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[772].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[772]),
        .S(self_sf7[772]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[773].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[773]),
        .S(self_sf7[773]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[774].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[774]),
        .S(self_sf7[774]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[775].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[775]),
        .S(self_sf7[775]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[776].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[776]),
        .S(self_sf7[776]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[777].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[777]),
        .S(self_sf7[777]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[778].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[778]),
        .S(self_sf7[778]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[779].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[779]),
        .S(self_sf7[779]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[77].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[77]),
        .S(self_sf7[77]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[780].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[780]),
        .S(self_sf7[780]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[781].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[781]),
        .S(self_sf7[781]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[782].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[782]),
        .S(self_sf7[782]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[783].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[783]),
        .S(self_sf7[783]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[784].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[784]),
        .S(self_sf7[784]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[785].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[785]),
        .S(self_sf7[785]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[786].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[786]),
        .S(self_sf7[786]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[787].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[787]),
        .S(self_sf7[787]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[788].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[788]),
        .S(self_sf7[788]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[789].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[789]),
        .S(self_sf7[789]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[78].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[78]),
        .S(self_sf7[78]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[790].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[790]),
        .S(self_sf7[790]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[791].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[791]),
        .S(self_sf7[791]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[792].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[792]),
        .S(self_sf7[792]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[793].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[793]),
        .S(self_sf7[793]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[794].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[794]),
        .S(self_sf7[794]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[795].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[795]),
        .S(self_sf7[795]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[796].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[796]),
        .S(self_sf7[796]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[797].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[797]),
        .S(self_sf7[797]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[798].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[798]),
        .S(self_sf7[798]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[799].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[799]),
        .S(self_sf7[799]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[79].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[79]),
        .S(self_sf7[79]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[7].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[7]),
        .S(info_sf7[7]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[800].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[800]),
        .S(self_sf7[800]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[801].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[801]),
        .S(self_sf7[801]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[802].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[802]),
        .S(self_sf7[802]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[803].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[803]),
        .S(self_sf7[803]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[804].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[804]),
        .S(self_sf7[804]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[805].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[805]),
        .S(self_sf7[805]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[806].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[806]),
        .S(self_sf7[806]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[807].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[807]),
        .S(self_sf7[807]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[808].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[808]),
        .S(self_sf7[808]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[809].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[809]),
        .S(self_sf7[809]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[80].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[80]),
        .S(self_sf7[80]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[810].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[810]),
        .S(self_sf7[810]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[811].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[811]),
        .S(self_sf7[811]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[812].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[812]),
        .S(self_sf7[812]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[813].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[813]),
        .S(self_sf7[813]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[814].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[814]),
        .S(self_sf7[814]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[815].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[815]),
        .S(self_sf7[815]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[816].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[816]),
        .S(self_sf7[816]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[817].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[817]),
        .S(self_sf7[817]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[818].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[818]),
        .S(self_sf7[818]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[819].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[819]),
        .S(self_sf7[819]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[81].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[81]),
        .S(self_sf7[81]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[820].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[820]),
        .S(self_sf7[820]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[821].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[821]),
        .S(self_sf7[821]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[822].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[822]),
        .S(self_sf7[822]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[823].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[823]),
        .S(self_sf7[823]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[824].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[824]),
        .S(self_sf7[824]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[825].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[825]),
        .S(self_sf7[825]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[826].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[826]),
        .S(self_sf7[826]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[827].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[827]),
        .S(self_sf7[827]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[828].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[828]),
        .S(self_sf7[828]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[829].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[829]),
        .S(self_sf7[829]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[82].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[82]),
        .S(self_sf7[82]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[830].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[830]),
        .S(self_sf7[830]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[831].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[831]),
        .S(self_sf7[831]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[832].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[832]),
        .S(self_sf7[832]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[833].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[833]),
        .S(self_sf7[833]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[834].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[834]),
        .S(self_sf7[834]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[835].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[835]),
        .S(self_sf7[835]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[836].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[836]),
        .S(self_sf7[836]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[837].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[837]),
        .S(self_sf7[837]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[838].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[838]),
        .S(self_sf7[838]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[839].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[839]),
        .S(self_sf7[839]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[83].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[83]),
        .S(self_sf7[83]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[840].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[840]),
        .S(self_sf7[840]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[841].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[841]),
        .S(self_sf7[841]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[842].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[842]),
        .S(self_sf7[842]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[843].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[843]),
        .S(self_sf7[843]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[844].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[844]),
        .S(self_sf7[844]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[845].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[845]),
        .S(self_sf7[845]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[846].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[846]),
        .S(self_sf7[846]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[847].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[847]),
        .S(self_sf7[847]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[848].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[848]),
        .S(self_sf7[848]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[849].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[849]),
        .S(self_sf7[849]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[84].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[84]),
        .S(self_sf7[84]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[850].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[850]),
        .S(self_sf7[850]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[851].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[851]),
        .S(self_sf7[851]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[852].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[852]),
        .S(self_sf7[852]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[853].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[853]),
        .S(self_sf7[853]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[854].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[854]),
        .S(self_sf7[854]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[855].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[855]),
        .S(self_sf7[855]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[856].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[856]),
        .S(self_sf7[856]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[857].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[857]),
        .S(self_sf7[857]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[858].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[858]),
        .S(self_sf7[858]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[859].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[859]),
        .S(self_sf7[859]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[85].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[85]),
        .S(self_sf7[85]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[860].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[860]),
        .S(self_sf7[860]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[861].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[861]),
        .S(self_sf7[861]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[862].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[862]),
        .S(self_sf7[862]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[863].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[863]),
        .S(self_sf7[863]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[864].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[864]),
        .S(self_sf7[864]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[865].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[865]),
        .S(self_sf7[865]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[866].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[866]),
        .S(self_sf7[866]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[867].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[867]),
        .S(self_sf7[867]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[868].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[868]),
        .S(self_sf7[868]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[869].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[869]),
        .S(self_sf7[869]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[86].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[86]),
        .S(self_sf7[86]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[870].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[870]),
        .S(self_sf7[870]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[871].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[871]),
        .S(self_sf7[871]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[872].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[872]),
        .S(self_sf7[872]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[873].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[873]),
        .S(self_sf7[873]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[874].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[874]),
        .S(self_sf7[874]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[875].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[875]),
        .S(self_sf7[875]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[876].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[876]),
        .S(self_sf7[876]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[877].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[877]),
        .S(self_sf7[877]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[878].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[878]),
        .S(self_sf7[878]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[879].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[879]),
        .S(self_sf7[879]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[87].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[87]),
        .S(self_sf7[87]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[880].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[880]),
        .S(self_sf7[880]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[881].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[881]),
        .S(self_sf7[881]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[882].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[882]),
        .S(self_sf7[882]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[883].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[883]),
        .S(self_sf7[883]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[884].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[884]),
        .S(self_sf7[884]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[885].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[885]),
        .S(self_sf7[885]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[886].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[886]),
        .S(self_sf7[886]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[887].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[887]),
        .S(self_sf7[887]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[888].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[888]),
        .S(self_sf7[888]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[889].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[889]),
        .S(self_sf7[889]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[88].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[88]),
        .S(self_sf7[88]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[890].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[890]),
        .S(self_sf7[890]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[891].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[891]),
        .S(self_sf7[891]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[892].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[892]),
        .S(self_sf7[892]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[893].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[893]),
        .S(self_sf7[893]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[894].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[894]),
        .S(self_sf7[894]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[895].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[895]),
        .S(self_sf7[895]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[896].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[896]),
        .S(self_sf7[896]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[897].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[897]),
        .S(self_sf7[897]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[898].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[898]),
        .S(self_sf7[898]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[899].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[899]),
        .S(self_sf7[899]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[89].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[89]),
        .S(self_sf7[89]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[8].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[8]),
        .S(self_sf7[8]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[900].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[900]),
        .S(self_sf7[900]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[901].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[901]),
        .S(self_sf7[901]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[902].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[902]),
        .S(self_sf7[902]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[903].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[903]),
        .S(self_sf7[903]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[904].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[904]),
        .S(self_sf7[904]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[905].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[905]),
        .S(self_sf7[905]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[906].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[906]),
        .S(self_sf7[906]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[907].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[907]),
        .S(self_sf7[907]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[908].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[908]),
        .S(self_sf7[908]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[909].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[909]),
        .S(self_sf7[909]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[90].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[90]),
        .S(self_sf7[90]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[910].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[910]),
        .S(self_sf7[910]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[911].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[911]),
        .S(self_sf7[911]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[912].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[912]),
        .S(self_sf7[912]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[913].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[913]),
        .S(self_sf7[913]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[914].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[914]),
        .S(self_sf7[914]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[915].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[915]),
        .S(self_sf7[915]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[916].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[916]),
        .S(self_sf7[916]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[917].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[917]),
        .S(self_sf7[917]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[918].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[918]),
        .S(self_sf7[918]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[919].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[919]),
        .S(self_sf7[919]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[91].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[91]),
        .S(self_sf7[91]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[920].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[920]),
        .S(self_sf7[920]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[921].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[921]),
        .S(self_sf7[921]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[922].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[922]),
        .S(self_sf7[922]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[923].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[923]),
        .S(self_sf7[923]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[924].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[924]),
        .S(self_sf7[924]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[925].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[925]),
        .S(self_sf7[925]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[926].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[926]),
        .S(self_sf7[926]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[927].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[927]),
        .S(self_sf7[927]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[928].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[928]),
        .S(self_sf7[928]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[929].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[929]),
        .S(self_sf7[929]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[92].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[92]),
        .S(self_sf7[92]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[930].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[930]),
        .S(self_sf7[930]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[931].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[931]),
        .S(self_sf7[931]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[932].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[932]),
        .S(self_sf7[932]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[933].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[933]),
        .S(self_sf7[933]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[934].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[934]),
        .S(self_sf7[934]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[935].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[935]),
        .S(self_sf7[935]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[936].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[936]),
        .S(self_sf7[936]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[937].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[937]),
        .S(self_sf7[937]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[938].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[938]),
        .S(self_sf7[938]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[939].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[939]),
        .S(self_sf7[939]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[93].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[93]),
        .S(self_sf7[93]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[940].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[940]),
        .S(self_sf7[940]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[941].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[941]),
        .S(self_sf7[941]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[942].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[942]),
        .S(self_sf7[942]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[943].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[943]),
        .S(self_sf7[943]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[944].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[944]),
        .S(self_sf7[944]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[945].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[945]),
        .S(self_sf7[945]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[946].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[946]),
        .S(self_sf7[946]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[947].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[947]),
        .S(self_sf7[947]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[948].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[948]),
        .S(self_sf7[948]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[949].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[949]),
        .S(self_sf7[949]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[94].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[94]),
        .S(self_sf7[94]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[950].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[950]),
        .S(self_sf7[950]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[951].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[951]),
        .S(self_sf7[951]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[952].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[952]),
        .S(self_sf7[952]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[953].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[953]),
        .S(self_sf7[953]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[954].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[954]),
        .S(self_sf7[954]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[955].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[955]),
        .S(self_sf7[955]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[956].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[956]),
        .S(self_sf7[956]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[957].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[957]),
        .S(self_sf7[957]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[958].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[958]),
        .S(self_sf7[958]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[959].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[959]),
        .S(self_sf7[959]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[95].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[95]),
        .S(self_sf7[95]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[960].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[960]),
        .S(self_sf7[960]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[961].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[961]),
        .S(self_sf7[961]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[962].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[962]),
        .S(self_sf7[962]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[963].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[963]),
        .S(self_sf7[963]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[964].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[964]),
        .S(self_sf7[964]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[965].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[965]),
        .S(self_sf7[965]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[966].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[966]),
        .S(self_sf7[966]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[967].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[967]),
        .S(self_sf7[967]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[968].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[968]),
        .S(self_sf7[968]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[969].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[969]),
        .S(self_sf7[969]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[96].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[96]),
        .S(self_sf7[96]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[970].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[970]),
        .S(self_sf7[970]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[971].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[971]),
        .S(self_sf7[971]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[972].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[972]),
        .S(self_sf7[972]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[973].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[973]),
        .S(self_sf7[973]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[974].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[974]),
        .S(self_sf7[974]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[975].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[975]),
        .S(self_sf7[975]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[976].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[976]),
        .S(self_sf7[976]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[977].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[977]),
        .S(self_sf7[977]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[978].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[978]),
        .S(self_sf7[978]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[979].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[979]),
        .S(self_sf7[979]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[97].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[97]),
        .S(self_sf7[97]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[980].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[980]),
        .S(self_sf7[980]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[981].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[981]),
        .S(self_sf7[981]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[982].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[982]),
        .S(self_sf7[982]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[983].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[983]),
        .S(self_sf7[983]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[984].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[984]),
        .S(self_sf7[984]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[985].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[985]),
        .S(self_sf7[985]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[986].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[986]),
        .S(self_sf7[986]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[987].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[987]),
        .S(self_sf7[987]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[988].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[988]),
        .S(self_sf7[988]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[989].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[989]),
        .S(self_sf7[989]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[98].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[98]),
        .S(self_sf7[98]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[990].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[990]),
        .S(self_sf7[990]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[991].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[991]),
        .S(self_sf7[991]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[992].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[992]),
        .S(self_sf7[992]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[993].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[993]),
        .S(self_sf7[993]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[994].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[994]),
        .S(self_sf7[994]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[995].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[995]),
        .S(self_sf7[995]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[996].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[996]),
        .S(self_sf7[996]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[997].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[997]),
        .S(self_sf7[997]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[998].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[998]),
        .S(self_sf7[998]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[999].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[999]),
        .S(self_sf7[999]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[99].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[99]),
        .S(self_sf7[99]));
  (* BOX_TYPE = "black_box" *) 
  MUXF7 \activity_ROsf7[9].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf7[9]),
        .S(self_sf7[9]));
  (* BOX_TYPE = "black_box" *) 
  MUXF8 \activity_ROsf8[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf8[0]),
        .S(self_sf8[0]));
  (* BOX_TYPE = "black_box" *) 
  MUXF9 \activity_ROsf9[0].ro_inv 
       (.I0(enable_i),
        .I1(1'b0),
        .O(self_sf9[0]),
        .S(self_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_0
       (.I0(1'b0),
        .O(self_sf7[1802]));
  LUT1 #(
    .INIT(2'h2)) 
    i_1
       (.I0(1'b0),
        .O(self_sf7[1801]));
  LUT1 #(
    .INIT(2'h2)) 
    i_10
       (.I0(1'b0),
        .O(info_sf8[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_11
       (.I0(1'b0),
        .O(info_sf8[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_12
       (.I0(1'b0),
        .O(info_sf8[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_13
       (.I0(1'b0),
        .O(info_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_14
       (.I0(1'b0),
        .O(info_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_15
       (.I0(1'b0),
        .O(info_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_16
       (.I0(1'b0),
        .O(info_sf8[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_17
       (.I0(1'b0),
        .O(info_sf9[7]));
  LUT1 #(
    .INIT(2'h2)) 
    i_18
       (.I0(1'b0),
        .O(info_sf9[6]));
  LUT1 #(
    .INIT(2'h2)) 
    i_19
       (.I0(1'b0),
        .O(info_sf9[5]));
  LUT1 #(
    .INIT(2'h2)) 
    i_2
       (.I0(1'b0),
        .O(self_sf7[1800]));
  LUT1 #(
    .INIT(2'h2)) 
    i_20
       (.I0(1'b0),
        .O(info_sf9[4]));
  LUT1 #(
    .INIT(2'h2)) 
    i_21
       (.I0(1'b0),
        .O(info_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_22
       (.I0(1'b0),
        .O(info_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_23
       (.I0(1'b0),
        .O(info_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_24
       (.I0(1'b0),
        .O(info_sf9[0]));
  LUT1 #(
    .INIT(2'h2)) 
    i_3
       (.I0(1'b0),
        .O(self_sf8[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_4
       (.I0(1'b0),
        .O(self_sf8[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_5
       (.I0(1'b0),
        .O(self_sf8[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_6
       (.I0(1'b0),
        .O(self_sf9[3]));
  LUT1 #(
    .INIT(2'h2)) 
    i_7
       (.I0(1'b0),
        .O(self_sf9[2]));
  LUT1 #(
    .INIT(2'h2)) 
    i_8
       (.I0(1'b0),
        .O(self_sf9[1]));
  LUT1 #(
    .INIT(2'h2)) 
    i_9
       (.I0(1'b0),
        .O(info_sf8[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst
       (.I0(self_sf7[7]),
        .O(info_sf7[7]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__0
       (.I0(self_sf7[6]),
        .O(info_sf7[6]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__1
       (.I0(self_sf7[5]),
        .O(info_sf7[5]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__2
       (.I0(self_sf7[4]),
        .O(info_sf7[4]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__3
       (.I0(self_sf7[3]),
        .O(info_sf7[3]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__4
       (.I0(self_sf7[2]),
        .O(info_sf7[2]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__5
       (.I0(self_sf7[1]),
        .O(info_sf7[1]));
  LUT1 #(
    .INIT(2'h2)) 
    self_sf7_inst__6
       (.I0(self_sf7[0]),
        .O(info_sf7[0]));
endmodule
`ifndef GLBL
`define GLBL
`timescale  1 ps / 1 ps

module glbl ();

    parameter ROC_WIDTH = 100000;
    parameter TOC_WIDTH = 0;

//--------   STARTUP Globals --------------
    wire GSR;
    wire GTS;
    wire GWE;
    wire PRLD;
    tri1 p_up_tmp;
    tri (weak1, strong0) PLL_LOCKG = p_up_tmp;

    wire PROGB_GLBL;
    wire CCLKO_GLBL;
    wire FCSBO_GLBL;
    wire [3:0] DO_GLBL;
    wire [3:0] DI_GLBL;
   
    reg GSR_int;
    reg GTS_int;
    reg PRLD_int;

//--------   JTAG Globals --------------
    wire JTAG_TDO_GLBL;
    wire JTAG_TCK_GLBL;
    wire JTAG_TDI_GLBL;
    wire JTAG_TMS_GLBL;
    wire JTAG_TRST_GLBL;

    reg JTAG_CAPTURE_GLBL;
    reg JTAG_RESET_GLBL;
    reg JTAG_SHIFT_GLBL;
    reg JTAG_UPDATE_GLBL;
    reg JTAG_RUNTEST_GLBL;

    reg JTAG_SEL1_GLBL = 0;
    reg JTAG_SEL2_GLBL = 0 ;
    reg JTAG_SEL3_GLBL = 0;
    reg JTAG_SEL4_GLBL = 0;

    reg JTAG_USER_TDO1_GLBL = 1'bz;
    reg JTAG_USER_TDO2_GLBL = 1'bz;
    reg JTAG_USER_TDO3_GLBL = 1'bz;
    reg JTAG_USER_TDO4_GLBL = 1'bz;

    assign (strong1, weak0) GSR = GSR_int;
    assign (strong1, weak0) GTS = GTS_int;
    assign (weak1, weak0) PRLD = PRLD_int;

    initial begin
	GSR_int = 1'b1;
	PRLD_int = 1'b1;
	#(ROC_WIDTH)
	GSR_int = 1'b0;
	PRLD_int = 1'b0;
    end

    initial begin
	GTS_int = 1'b1;
	#(TOC_WIDTH)
	GTS_int = 1'b0;
    end

endmodule
`endif
